* NGSPICE file created from NfiVe32_SYS.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt NfiVe32_SYS HADDR[0] HADDR[10] HADDR[11] HADDR[12] HADDR[13] HADDR[14] HADDR[15]
+ HADDR[16] HADDR[17] HADDR[18] HADDR[19] HADDR[1] HADDR[20] HADDR[21] HADDR[22] HADDR[23]
+ HADDR[24] HADDR[25] HADDR[26] HADDR[27] HADDR[28] HADDR[29] HADDR[2] HADDR[30] HADDR[31]
+ HADDR[3] HADDR[4] HADDR[5] HADDR[6] HADDR[7] HADDR[8] HADDR[9] HCLK HRDATA[0] HRDATA[10]
+ HRDATA[11] HRDATA[12] HRDATA[13] HRDATA[14] HRDATA[15] HRDATA[16] HRDATA[17] HRDATA[18]
+ HRDATA[19] HRDATA[1] HRDATA[20] HRDATA[21] HRDATA[22] HRDATA[23] HRDATA[24] HRDATA[25]
+ HRDATA[26] HRDATA[27] HRDATA[28] HRDATA[29] HRDATA[2] HRDATA[30] HRDATA[31] HRDATA[3]
+ HRDATA[4] HRDATA[5] HRDATA[6] HRDATA[7] HRDATA[8] HRDATA[9] HREADY HRESETn HSIZE[0]
+ HSIZE[1] HSIZE[2] HTRANS[0] HTRANS[1] HWDATA[0] HWDATA[10] HWDATA[11] HWDATA[12]
+ HWDATA[13] HWDATA[14] HWDATA[15] HWDATA[16] HWDATA[17] HWDATA[18] HWDATA[19] HWDATA[1]
+ HWDATA[20] HWDATA[21] HWDATA[22] HWDATA[23] HWDATA[24] HWDATA[25] HWDATA[26] HWDATA[27]
+ HWDATA[28] HWDATA[29] HWDATA[2] HWDATA[30] HWDATA[31] HWDATA[3] HWDATA[4] HWDATA[5]
+ HWDATA[6] HWDATA[7] HWDATA[8] HWDATA[9] HWRITE IRQ[0] IRQ[10] IRQ[11] IRQ[12] IRQ[13]
+ IRQ[14] IRQ[15] IRQ[16] IRQ[17] IRQ[18] IRQ[19] IRQ[1] IRQ[20] IRQ[21] IRQ[22] IRQ[23]
+ IRQ[24] IRQ[25] IRQ[26] IRQ[27] IRQ[28] IRQ[29] IRQ[2] IRQ[30] IRQ[31] IRQ[3] IRQ[4]
+ IRQ[5] IRQ[6] IRQ[7] IRQ[8] IRQ[9] NMI SYSTICKCLKDIV[0] SYSTICKCLKDIV[1] SYSTICKCLKDIV[2]
+ SYSTICKCLKDIV[3] SYSTICKCLKDIV[4] SYSTICKCLKDIV[5] SYSTICKCLKDIV[6] SYSTICKCLKDIV[7]
+ VPWR VGND
XANTENNA__21917__A2 _21916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15814__B _15869_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18869_ _15651_/X _18863_/X _20727_/A _18864_/X VGND VGND VPWR VPWR _24417_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18794__A1 _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20900_ HRDATA[5] VGND VGND VPWR VPWR _20900_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21880_ _21879_/X _21875_/X _15351_/B _21870_/X VGND VGND VPWR VPWR _21880_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22928__A _22927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20831_ _20782_/X _20830_/X _11523_/A _20789_/X VGND VGND VPWR VPWR _20831_/X sky130_fd_sc_hd__o22a_4
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22878__B1 _17397_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15830__A _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23550_ _23997_/CLK _21976_/X VGND VGND VPWR VPWR _23550_/Q sky130_fd_sc_hd__dfxtp_4
X_20762_ _20754_/X _20760_/X _19141_/A _20761_/X VGND VGND VPWR VPWR _20762_/X sky130_fd_sc_hd__o22a_4
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21550__B1 _23787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22501_ _22508_/A VGND VGND VPWR VPWR _22501_/X sky130_fd_sc_hd__buf_2
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23481_ _23294_/CLK _22083_/X VGND VGND VPWR VPWR _14834_/B sky130_fd_sc_hd__dfxtp_4
X_20693_ _21283_/A VGND VGND VPWR VPWR _20693_/X sky130_fd_sc_hd__buf_2
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22432_ _22117_/A VGND VGND VPWR VPWR _22432_/X sky130_fd_sc_hd__buf_2
XFILLER_149_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16309__B1 _11608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14165__B _23103_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22363_ _22097_/X _22362_/X _12128_/B _22359_/X VGND VGND VPWR VPWR _23315_/D sky130_fd_sc_hd__o22a_4
XFILLER_11_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24102_ _24102_/CLK _20615_/X VGND VGND VPWR VPWR _24102_/Q sky130_fd_sc_hd__dfxtp_4
X_21314_ _21313_/X _21305_/X _14871_/B _21239_/X VGND VGND VPWR VPWR _23926_/D sky130_fd_sc_hd__o22a_4
X_22294_ _22294_/A VGND VGND VPWR VPWR _22294_/X sky130_fd_sc_hd__buf_2
X_24033_ _23303_/CLK _24033_/D VGND VGND VPWR VPWR _24033_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_105_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21245_ _21269_/A VGND VGND VPWR VPWR _21245_/X sky130_fd_sc_hd__buf_2
XANTENNA__15277__A _14169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14181__A _14225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20813__C1 _20812_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21176_ _21136_/A VGND VGND VPWR VPWR _21176_/X sky130_fd_sc_hd__buf_2
XFILLER_104_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12413__B _23660_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20127_ _20118_/Y _20126_/X _18960_/X VGND VGND VPWR VPWR _20127_/X sky130_fd_sc_hd__and3_4
XANTENNA__21908__A2 _21902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20058_ _20040_/X _18402_/A _20046_/X _20057_/X VGND VGND VPWR VPWR _20058_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22030__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11900_ _11900_/A VGND VGND VPWR VPWR _12854_/A sky130_fd_sc_hd__buf_2
X_12880_ _12472_/A _12880_/B _12880_/C VGND VGND VPWR VPWR _12881_/C sky130_fd_sc_hd__and3_4
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23817_ _24073_/CLK _23817_/D VGND VGND VPWR VPWR _12964_/B sky130_fd_sc_hd__dfxtp_4
X_11831_ _11786_/X _11823_/X _11830_/X VGND VGND VPWR VPWR _11831_/X sky130_fd_sc_hd__and3_4
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15740__A _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14482_/X _14549_/Y VGND VGND VPWR VPWR _15389_/B sky130_fd_sc_hd__or2_4
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _23750_/CLK _23748_/D VGND VGND VPWR VPWR _23748_/Q sky130_fd_sc_hd__dfxtp_4
X_11762_ _11742_/X VGND VGND VPWR VPWR _11762_/X sky130_fd_sc_hd__buf_2
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20358__A _20358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13532_/A _23781_/Q VGND VGND VPWR VPWR _13501_/X sky130_fd_sc_hd__or2_4
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _13016_/A _14458_/X _14465_/X _14472_/X _14480_/X VGND VGND VPWR VPWR _14481_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _16205_/A VGND VGND VPWR VPWR _11693_/X sky130_fd_sc_hd__buf_2
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23679_ _23679_/CLK _21742_/X VGND VGND VPWR VPWR _23679_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16220_/A _16218_/X _16220_/C VGND VGND VPWR VPWR _16221_/C sky130_fd_sc_hd__and3_4
XANTENNA__13260__A _12978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _13431_/X _23301_/Q VGND VGND VPWR VPWR _13433_/C sky130_fd_sc_hd__or2_4
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16151_ _16116_/A _16151_/B _16150_/X VGND VGND VPWR VPWR _16151_/X sky130_fd_sc_hd__and3_4
X_13363_ _13415_/A _13363_/B _13363_/C VGND VGND VPWR VPWR _13363_/X sky130_fd_sc_hd__and3_4
XANTENNA__21844__B2 _21834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17667__A _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15102_ _15078_/A _15102_/B _15101_/X VGND VGND VPWR VPWR _15102_/X sky130_fd_sc_hd__and3_4
X_12314_ _13184_/A _12314_/B VGND VGND VPWR VPWR _12315_/C sky130_fd_sc_hd__or2_4
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16082_ _11759_/X _16078_/X _16081_/X VGND VGND VPWR VPWR _16082_/X sky130_fd_sc_hd__or3_4
X_13294_ _13320_/A _13294_/B VGND VGND VPWR VPWR _13294_/X sky130_fd_sc_hd__or2_4
XFILLER_6_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19910_ _23083_/D _19909_/X VGND VGND VPWR VPWR _19910_/X sky130_fd_sc_hd__or2_4
XANTENNA__15187__A _15076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15033_ _12495_/A _15033_/B VGND VGND VPWR VPWR _15033_/X sky130_fd_sc_hd__or2_4
X_12245_ _13301_/A _12376_/B VGND VGND VPWR VPWR _12246_/C sky130_fd_sc_hd__or2_4
XANTENNA__12604__A _12604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14091__A _14138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21072__A2 _21066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12176_ _12138_/A _12172_/X _12175_/X VGND VGND VPWR VPWR _12176_/X sky130_fd_sc_hd__or3_4
X_19841_ _19662_/B _19868_/B _19691_/Y VGND VGND VPWR VPWR _19842_/A sky130_fd_sc_hd__o21a_4
XFILLER_122_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20821__A HRDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15915__A _15849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16984_ _17708_/A _18403_/B VGND VGND VPWR VPWR _17906_/B sky130_fd_sc_hd__or2_4
X_19772_ _19469_/X _19771_/X _16684_/A _19515_/X VGND VGND VPWR VPWR _19772_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_27_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15935_ _15934_/X VGND VGND VPWR VPWR _15971_/A sky130_fd_sc_hd__buf_2
X_18723_ _16971_/A _18722_/Y _17749_/X VGND VGND VPWR VPWR _18723_/X sky130_fd_sc_hd__a21o_4
XFILLER_77_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_24_0_HCLK clkbuf_6_12_0_HCLK/X VGND VGND VPWR VPWR _24302_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_114_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13435__A _12889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18654_ _17805_/X _18054_/Y _17869_/A _18653_/X VGND VGND VPWR VPWR _18654_/X sky130_fd_sc_hd__a211o_4
X_15866_ _13540_/X _15866_/B VGND VGND VPWR VPWR _15866_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_87_0_HCLK clkbuf_7_86_0_HCLK/A VGND VGND VPWR VPWR _23290_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17605_ _18290_/A _17508_/X _17517_/A _17605_/D VGND VGND VPWR VPWR _17605_/X sky130_fd_sc_hd__or4_4
X_14817_ _14685_/A _14817_/B _14817_/C VGND VGND VPWR VPWR _14818_/C sky130_fd_sc_hd__and3_4
X_18585_ _17111_/X _18157_/Y _17869_/X _18584_/Y VGND VGND VPWR VPWR _18585_/X sky130_fd_sc_hd__a211o_4
X_15797_ _12848_/A _15797_/B VGND VGND VPWR VPWR _15797_/X sky130_fd_sc_hd__or2_4
XANTENNA__16746__A _11963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17536_ _17528_/A _17535_/X VGND VGND VPWR VPWR _17536_/Y sky130_fd_sc_hd__nor2_4
XFILLER_83_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15650__A _11668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14748_ _11913_/A _14748_/B _14748_/C VGND VGND VPWR VPWR _14749_/C sky130_fd_sc_hd__and3_4
XFILLER_32_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20268__A _20267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24332__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17467_ _12842_/X _17467_/B VGND VGND VPWR VPWR _17467_/X sky130_fd_sc_hd__or2_4
XANTENNA__14014__A1 _13951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14679_ _14679_/A _23418_/Q VGND VGND VPWR VPWR _14680_/C sky130_fd_sc_hd__or2_4
X_16418_ _13475_/A _16414_/X _16417_/X VGND VGND VPWR VPWR _16419_/B sky130_fd_sc_hd__or3_4
X_19206_ _24318_/Q _19138_/X _19205_/Y VGND VGND VPWR VPWR _19206_/X sky130_fd_sc_hd__o21a_4
XFILLER_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17398_ _17398_/A VGND VGND VPWR VPWR _17398_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19137_ _19137_/A _19211_/A VGND VGND VPWR VPWR _19138_/B sky130_fd_sc_hd__and2_4
X_16349_ _16314_/X _16347_/X _16348_/X VGND VGND VPWR VPWR _16349_/X sky130_fd_sc_hd__and3_4
XANTENNA__21835__B2 _21834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16481__A _13385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19068_ _19024_/A VGND VGND VPWR VPWR _19068_/X sky130_fd_sc_hd__buf_2
XFILLER_172_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18019_ _16933_/Y VGND VGND VPWR VPWR _18019_/X sky130_fd_sc_hd__buf_2
XANTENNA__15097__A _15081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19792__A HRDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21030_ _21030_/A VGND VGND VPWR VPWR _21134_/D sky130_fd_sc_hd__buf_2
XANTENNA__21827__A _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22260__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15825__A _12866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22012__A1 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22012__B2 _22007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22981_ _22978_/X _22981_/B _22981_/C VGND VGND VPWR VPWR _22981_/X sky130_fd_sc_hd__and3_4
XFILLER_67_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22563__A2 _22558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13345__A _13384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21932_ _21877_/X _21930_/X _14728_/B _21927_/X VGND VGND VPWR VPWR _23577_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22658__A _22658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21863_ _21808_/A VGND VGND VPWR VPWR _21863_/X sky130_fd_sc_hd__buf_2
X_23602_ _23537_/CLK _23602_/D VGND VGND VPWR VPWR _23602_/Q sky130_fd_sc_hd__dfxtp_4
X_20814_ _20814_/A VGND VGND VPWR VPWR _20814_/Y sky130_fd_sc_hd__inv_2
X_21794_ _21582_/X _21791_/X _23645_/Q _21788_/X VGND VGND VPWR VPWR _21794_/X sky130_fd_sc_hd__o22a_4
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23533_ _23533_/CLK _22005_/X VGND VGND VPWR VPWR _16167_/B sky130_fd_sc_hd__dfxtp_4
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20745_ _20745_/A VGND VGND VPWR VPWR _20745_/X sky130_fd_sc_hd__buf_2
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13080__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22079__A1 _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23464_ _23496_/CLK _22126_/X VGND VGND VPWR VPWR _13013_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22079__B2 _22078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20676_ _20447_/A VGND VGND VPWR VPWR _20676_/X sky130_fd_sc_hd__buf_2
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12408__B _24108_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20629__A2 _20443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17487__A _12680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22415_ _22412_/X _22414_/X _12114_/B _22409_/X VGND VGND VPWR VPWR _22415_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16391__A _16009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23395_ _23523_/CLK _22253_/X VGND VGND VPWR VPWR _15829_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22346_ _22346_/A VGND VGND VPWR VPWR _23324_/D sky130_fd_sc_hd__buf_2
XFILLER_124_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12319__A1 _11856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23697__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22277_ _22284_/A VGND VGND VPWR VPWR _22277_/X sky130_fd_sc_hd__buf_2
XFILLER_152_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12424__A _12466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22840__B _14483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12030_ _16595_/A VGND VGND VPWR VPWR _16702_/A sky130_fd_sc_hd__buf_2
XANTENNA__21054__A2 _21052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24016_ _24080_/CLK _21146_/X VGND VGND VPWR VPWR _16406_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_3_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21228_ _20938_/X _21226_/X _14737_/B _21223_/X VGND VGND VPWR VPWR _23961_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15735__A _12783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21159_ _21152_/A VGND VGND VPWR VPWR _21159_/X sky130_fd_sc_hd__buf_2
XANTENNA__18111__A _18111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15454__B _15454_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13981_ _13981_/A _13980_/X VGND VGND VPWR VPWR _13981_/X sky130_fd_sc_hd__and2_4
XFILLER_150_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13255__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22554__A2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15720_ _12762_/A _15658_/B VGND VGND VPWR VPWR _15720_/X sky130_fd_sc_hd__or2_4
X_12932_ _12951_/A _23945_/Q VGND VGND VPWR VPWR _12932_/X sky130_fd_sc_hd__or2_4
XFILLER_100_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15651_ _15651_/A VGND VGND VPWR VPWR _15651_/X sky130_fd_sc_hd__buf_2
X_12863_ _12863_/A _24041_/Q VGND VGND VPWR VPWR _12865_/B sky130_fd_sc_hd__or2_4
XANTENNA__24322__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22306__A2 _22301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14602_ _15408_/A _14600_/X _14601_/X VGND VGND VPWR VPWR _14602_/X sky130_fd_sc_hd__and3_4
X_11814_ _12978_/A VGND VGND VPWR VPWR _13416_/A sky130_fd_sc_hd__buf_2
X_18370_ _18358_/X _18370_/B VGND VGND VPWR VPWR _18370_/X sky130_fd_sc_hd__and2_4
X_15582_ _11855_/A _11629_/A _15551_/X _11606_/A _15581_/X VGND VGND VPWR VPWR _15582_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12833_/A _12794_/B VGND VGND VPWR VPWR _12798_/B sky130_fd_sc_hd__or2_4
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17321_ _19852_/A _17039_/X _12882_/A _17297_/X VGND VGND VPWR VPWR _17321_/X sky130_fd_sc_hd__o22a_4
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14533_ _14509_/A _14531_/X _14532_/X VGND VGND VPWR VPWR _14533_/X sky130_fd_sc_hd__and3_4
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13702__B _13702_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11745_ _12151_/A _11745_/B VGND VGND VPWR VPWR _11745_/X sky130_fd_sc_hd__or2_4
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14086__A _14086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17194__B1 _14701_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18781__A _18780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18930__A1 _14261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17252_ _17047_/X _17251_/X _17051_/X VGND VGND VPWR VPWR _17252_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14464_ _13011_/A _14464_/B _14464_/C VGND VGND VPWR VPWR _14464_/X sky130_fd_sc_hd__and3_4
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _12641_/A VGND VGND VPWR VPWR _13530_/A sky130_fd_sc_hd__buf_2
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20816__A _20857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16203_ _16219_/A _16203_/B VGND VGND VPWR VPWR _16204_/C sky130_fd_sc_hd__or2_4
XFILLER_174_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13415_ _13415_/A _13415_/B _13415_/C VGND VGND VPWR VPWR _13415_/X sky130_fd_sc_hd__and3_4
XFILLER_128_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17397__A _13863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17183_ _17132_/Y _17131_/X _15252_/X _17133_/X VGND VGND VPWR VPWR _17183_/X sky130_fd_sc_hd__o22a_4
X_14395_ _11781_/A _14384_/X _14394_/X VGND VGND VPWR VPWR _14395_/X sky130_fd_sc_hd__and3_4
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16134_ _16144_/A _16132_/X _16134_/C VGND VGND VPWR VPWR _16138_/B sky130_fd_sc_hd__and3_4
XFILLER_127_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13346_ _12834_/A VGND VGND VPWR VPWR _13385_/A sky130_fd_sc_hd__buf_2
XANTENNA__18694__B1 _17793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16065_ _16046_/A _23438_/Q VGND VGND VPWR VPWR _16066_/C sky130_fd_sc_hd__or2_4
X_13277_ _13277_/A VGND VGND VPWR VPWR _13309_/A sky130_fd_sc_hd__buf_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15016_ _13952_/A _23893_/Q VGND VGND VPWR VPWR _15016_/X sky130_fd_sc_hd__or2_4
X_12228_ _12228_/A VGND VGND VPWR VPWR _12727_/A sky130_fd_sc_hd__buf_2
XANTENNA__22242__B2 _22241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19824_ _19705_/B _19823_/X _19545_/A _19883_/A VGND VGND VPWR VPWR _19824_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15645__A _13885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12159_ _11746_/X _12159_/B VGND VGND VPWR VPWR _12159_/X sky130_fd_sc_hd__or2_4
XFILLER_110_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20270__B _19948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19755_ _19665_/A _19753_/X _19895_/A _19754_/X VGND VGND VPWR VPWR _19755_/X sky130_fd_sc_hd__a211o_4
X_16967_ _16967_/A VGND VGND VPWR VPWR _17727_/A sky130_fd_sc_hd__inv_2
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18956__A _18948_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13165__A _13301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22545__A2 _22544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18706_ _24472_/Q VGND VGND VPWR VPWR _18706_/Y sky130_fd_sc_hd__inv_2
X_15918_ _15914_/X _15917_/X VGND VGND VPWR VPWR _15919_/D sky130_fd_sc_hd__nand2_4
X_19686_ _19624_/B VGND VGND VPWR VPWR _19815_/B sky130_fd_sc_hd__buf_2
X_16898_ _16828_/X _16898_/B VGND VGND VPWR VPWR _16898_/X sky130_fd_sc_hd__and2_4
XANTENNA__22478__A _20958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15849_ _11857_/A _11631_/A _15818_/X _11607_/A _15848_/X VGND VGND VPWR VPWR _15849_/X
+ sky130_fd_sc_hd__a32o_4
X_18637_ _18095_/A _18637_/B VGND VGND VPWR VPWR _18637_/X sky130_fd_sc_hd__and2_4
XFILLER_65_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15380__A _15380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18568_ _18506_/X _18560_/Y _18561_/X _18563_/X _18567_/Y VGND VGND VPWR VPWR _18568_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17519_ _16786_/A _17378_/X _17379_/X VGND VGND VPWR VPWR _17520_/B sky130_fd_sc_hd__o21a_4
X_18499_ _18019_/X VGND VGND VPWR VPWR _18499_/X sky130_fd_sc_hd__buf_2
XANTENNA__12509__A _13042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17724__A2 _17427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20530_ _20530_/A VGND VGND VPWR VPWR _20531_/A sky130_fd_sc_hd__buf_2
XANTENNA__22925__B _22930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20461_ _20334_/A _20460_/X VGND VGND VPWR VPWR _20461_/X sky130_fd_sc_hd__or2_4
XANTENNA__14724__A _15444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22200_ _22132_/X _22194_/X _13546_/B _22198_/X VGND VGND VPWR VPWR _23429_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17100__A _17100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21284__A2 _21281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23180_ _23728_/CLK _23180_/D VGND VGND VPWR VPWR _12361_/B sky130_fd_sc_hd__dfxtp_4
X_20392_ _20358_/A _20391_/X VGND VGND VPWR VPWR _20392_/Y sky130_fd_sc_hd__nand2_4
XFILLER_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22941__A _22940_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22481__B2 _22421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22131_ _22129_/X _22123_/X _23462_/Q _22130_/X VGND VGND VPWR VPWR _23462_/D sky130_fd_sc_hd__o22a_4
XFILLER_173_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22062_ _21841_/X _22060_/X _23496_/Q _22057_/X VGND VGND VPWR VPWR _23496_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22233__B2 _22227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20461__A _20334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21013_ _20470_/A _21012_/X _24373_/Q _18893_/A VGND VGND VPWR VPWR _21013_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15555__A _11886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22964_ _22946_/X _18533_/A _22959_/X _22963_/X VGND VGND VPWR VPWR _22964_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21292__A _20801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21915_ _21848_/X _21909_/X _13447_/B _21913_/X VGND VGND VPWR VPWR _23589_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_70_0_HCLK clkbuf_6_35_0_HCLK/X VGND VGND VPWR VPWR _23095_/CLK sky130_fd_sc_hd__clkbuf_1
X_22895_ _19915_/X _22837_/X _15453_/Y _20665_/X VGND VGND VPWR VPWR _22895_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13803__A _14307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24495__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21846_ _21834_/A VGND VGND VPWR VPWR _21846_/X sky130_fd_sc_hd__buf_2
XFILLER_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14618__B _14618_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19697__A HRDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21777_ _21770_/A VGND VGND VPWR VPWR _21777_/X sky130_fd_sc_hd__buf_2
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18912__A1 _12678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ _11530_/A _11530_/B VGND VGND VPWR VPWR _11530_/X sky130_fd_sc_hd__or2_4
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23516_ _23515_/CLK _23516_/D VGND VGND VPWR VPWR _14339_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_141_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20728_ _24449_/Q VGND VGND VPWR VPWR _20730_/A sky130_fd_sc_hd__inv_2
X_24496_ _24158_/CLK _24496_/D HRESETn VGND VGND VPWR VPWR _19999_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20636__A _20895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23447_ _23095_/CLK _23447_/D VGND VGND VPWR VPWR _15150_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20659_ _21280_/A VGND VGND VPWR VPWR _20659_/X sky130_fd_sc_hd__buf_2
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ _12362_/A VGND VGND VPWR VPWR _13200_/X sky130_fd_sc_hd__buf_2
X_14180_ _14229_/A VGND VGND VPWR VPWR _14225_/A sky130_fd_sc_hd__buf_2
XFILLER_104_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23378_ _23537_/CLK _23378_/D VGND VGND VPWR VPWR _16615_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22472__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13131_ _12273_/A _23751_/Q VGND VGND VPWR VPWR _13131_/X sky130_fd_sc_hd__or2_4
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22329_ _23341_/Q VGND VGND VPWR VPWR _23341_/D sky130_fd_sc_hd__buf_2
XFILLER_3_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13062_ _13091_/A _13057_/X _13061_/X VGND VGND VPWR VPWR _13062_/X sky130_fd_sc_hd__or3_4
XFILLER_97_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12013_ _11951_/A _12013_/B _12013_/C VGND VGND VPWR VPWR _12013_/X sky130_fd_sc_hd__and3_4
XFILLER_105_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17870_ _17869_/X VGND VGND VPWR VPWR _17870_/X sky130_fd_sc_hd__buf_2
XANTENNA__17651__A1 _16943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16821_ _16821_/A _16821_/B VGND VGND VPWR VPWR _16822_/A sky130_fd_sc_hd__or2_4
XANTENNA__17651__B2 _17650_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16752_ _16639_/A _23537_/Q VGND VGND VPWR VPWR _16753_/C sky130_fd_sc_hd__or2_4
X_19540_ _24169_/Q _19481_/X HRDATA[21] _19482_/X VGND VGND VPWR VPWR _19540_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13964_ _13964_/A _23296_/Q VGND VGND VPWR VPWR _13965_/C sky130_fd_sc_hd__or2_4
XFILLER_93_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22298__A _22291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15703_ _12738_/A _15701_/X _15702_/X VGND VGND VPWR VPWR _15703_/X sky130_fd_sc_hd__and3_4
XFILLER_4_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12915_ _12948_/A _12915_/B VGND VGND VPWR VPWR _12915_/X sky130_fd_sc_hd__or2_4
XFILLER_59_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16683_ _16683_/A _16683_/B _16683_/C VGND VGND VPWR VPWR _16684_/C sky130_fd_sc_hd__and3_4
X_19471_ _19439_/A VGND VGND VPWR VPWR _19471_/X sky130_fd_sc_hd__buf_2
XFILLER_46_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13895_ _11780_/A VGND VGND VPWR VPWR _13928_/A sky130_fd_sc_hd__buf_2
X_18422_ _17396_/D _18421_/X _17448_/Y VGND VGND VPWR VPWR _18422_/Y sky130_fd_sc_hd__o21ai_4
X_15634_ _15610_/A _15634_/B VGND VGND VPWR VPWR _15634_/X sky130_fd_sc_hd__or2_4
XFILLER_64_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12846_ _12846_/A _12846_/B VGND VGND VPWR VPWR _12846_/X sky130_fd_sc_hd__or2_4
X_18353_ _18301_/A _18352_/X _18301_/A _18352_/X VGND VGND VPWR VPWR _18353_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21930__A _21923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15565_ _12186_/A _15561_/X _15564_/X VGND VGND VPWR VPWR _15565_/X sky130_fd_sc_hd__or3_4
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12604_/A VGND VGND VPWR VPWR _13051_/A sky130_fd_sc_hd__buf_2
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12329__A _12329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18903__A1 _17255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22745__B _22737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17304_ _17632_/A _17621_/B VGND VGND VPWR VPWR _17304_/X sky130_fd_sc_hd__and2_4
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14516_/A _14452_/B VGND VGND VPWR VPWR _14516_/X sky130_fd_sc_hd__or2_4
X_11728_ _16454_/A VGND VGND VPWR VPWR _16033_/A sky130_fd_sc_hd__buf_2
XANTENNA__15717__A1 _11856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18284_ _18284_/A VGND VGND VPWR VPWR _18284_/Y sky130_fd_sc_hd__inv_2
X_15496_ _13744_/A _15432_/B VGND VGND VPWR VPWR _15496_/X sky130_fd_sc_hd__or2_4
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17235_ _17128_/A VGND VGND VPWR VPWR _17825_/A sky130_fd_sc_hd__buf_2
X_14447_ _13601_/A _14503_/B VGND VGND VPWR VPWR _14447_/X sky130_fd_sc_hd__or2_4
X_11659_ _11659_/A VGND VGND VPWR VPWR _11660_/A sky130_fd_sc_hd__buf_2
XANTENNA__24218__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17166_ _15653_/X _17144_/X _17165_/Y _17146_/X VGND VGND VPWR VPWR _17166_/X sky130_fd_sc_hd__o22a_4
X_14378_ _14378_/A _23964_/Q VGND VGND VPWR VPWR _14378_/X sky130_fd_sc_hd__or2_4
XANTENNA__22463__B2 _22457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16117_ _16142_/A _23341_/Q VGND VGND VPWR VPWR _16117_/X sky130_fd_sc_hd__or2_4
X_13329_ _13320_/A _23654_/Q VGND VGND VPWR VPWR _13330_/C sky130_fd_sc_hd__or2_4
X_17097_ _17097_/A VGND VGND VPWR VPWR _18485_/A sky130_fd_sc_hd__buf_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16048_ _16048_/A _16048_/B VGND VGND VPWR VPWR _16048_/X sky130_fd_sc_hd__or2_4
XANTENNA__21377__A _21391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12999__A _12906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15375__A _11697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19807_ _19807_/A VGND VGND VPWR VPWR _19807_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17999_ _18288_/A _17998_/X VGND VGND VPWR VPWR _17999_/Y sky130_fd_sc_hd__nor2_4
X_19738_ _19619_/A _19736_/X _19603_/X _19737_/Y VGND VGND VPWR VPWR _19738_/X sky130_fd_sc_hd__a211o_4
XANTENNA__23392__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19669_ _19630_/X _19879_/C _19600_/X _19668_/X VGND VGND VPWR VPWR _19670_/B sky130_fd_sc_hd__a211o_4
Xclkbuf_6_57_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14719__A _14301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21700_ _21592_/X _21698_/X _14760_/B _21695_/X VGND VGND VPWR VPWR _23705_/D sky130_fd_sc_hd__o22a_4
XFILLER_77_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22680_ _22473_/X _22679_/X _14590_/B _22676_/X VGND VGND VPWR VPWR _22680_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22936__A _22910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21631_ _21624_/A VGND VGND VPWR VPWR _21631_/X sky130_fd_sc_hd__buf_2
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24350_ _24382_/CLK _19086_/X HRESETn VGND VGND VPWR VPWR _11524_/A sky130_fd_sc_hd__dfstp_4
X_21562_ _21560_/X _21554_/X _23782_/Q _21561_/X VGND VGND VPWR VPWR _21562_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20456__A _20313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23301_ _23397_/CLK _22382_/X VGND VGND VPWR VPWR _23301_/Q sky130_fd_sc_hd__dfxtp_4
X_20513_ _20251_/A _20512_/X _20306_/X VGND VGND VPWR VPWR _20513_/Y sky130_fd_sc_hd__o21ai_4
X_21493_ _21268_/X _21492_/X _12964_/B _21489_/X VGND VGND VPWR VPWR _23817_/D sky130_fd_sc_hd__o22a_4
X_24281_ _24292_/CLK _24281_/D HRESETn VGND VGND VPWR VPWR _19230_/A sky130_fd_sc_hd__dfrtp_4
X_20444_ _18779_/X VGND VGND VPWR VPWR _20444_/X sky130_fd_sc_hd__buf_2
X_23232_ _23617_/CLK _22521_/X VGND VGND VPWR VPWR _23232_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20375_ _20358_/A _20374_/X VGND VGND VPWR VPWR _20375_/Y sky130_fd_sc_hd__nand2_4
X_23163_ _24096_/CLK _22628_/X VGND VGND VPWR VPWR _14502_/B sky130_fd_sc_hd__dfxtp_4
X_22114_ _22113_/X _22111_/X _16196_/B _22106_/X VGND VGND VPWR VPWR _23469_/D sky130_fd_sc_hd__o22a_4
X_23094_ _23095_/CLK _23094_/D VGND VGND VPWR VPWR _14902_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22206__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22045_ _22041_/A VGND VGND VPWR VPWR _22060_/A sky130_fd_sc_hd__buf_2
XANTENNA__12702__A _12702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22509__A2 _22508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23996_ _23592_/CLK _23996_/D VGND VGND VPWR VPWR _23996_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23007__A _22908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22947_ _23080_/A VGND VGND VPWR VPWR _22947_/X sky130_fd_sc_hd__buf_2
XANTENNA__21193__B2 _21188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13533__A _12402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12700_ _13152_/A VGND VGND VPWR VPWR _13277_/A sky130_fd_sc_hd__buf_2
XFILLER_16_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13680_ _12300_/A _13678_/X _13680_/C VGND VGND VPWR VPWR _13680_/X sky130_fd_sc_hd__and3_4
X_22878_ _22876_/X _22820_/X _17397_/Y _22877_/X VGND VGND VPWR VPWR _22878_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22846__A _18780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12631_ _12646_/A _12500_/B VGND VGND VPWR VPWR _12631_/X sky130_fd_sc_hd__or2_4
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21829_ _20464_/A VGND VGND VPWR VPWR _21829_/X sky130_fd_sc_hd__buf_2
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_0_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR _24287_/CLK sky130_fd_sc_hd__clkbuf_1
X_15350_ _15372_/A _15348_/X _15349_/X VGND VGND VPWR VPWR _15354_/B sky130_fd_sc_hd__and3_4
X_12562_ _12903_/A _12559_/X _12562_/C VGND VGND VPWR VPWR _12562_/X sky130_fd_sc_hd__and3_4
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14301_ _14301_/A _14297_/X _14301_/C VGND VGND VPWR VPWR _14301_/X sky130_fd_sc_hd__or3_4
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11513_ _24406_/Q VGND VGND VPWR VPWR _11513_/Y sky130_fd_sc_hd__inv_2
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ _15281_/A _15280_/X VGND VGND VPWR VPWR _15281_/X sky130_fd_sc_hd__and2_4
X_12493_ _12493_/A VGND VGND VPWR VPWR _12903_/A sky130_fd_sc_hd__buf_2
X_24479_ _24137_/CLK _18552_/X HRESETn VGND VGND VPWR VPWR _24479_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17020_ _17019_/X VGND VGND VPWR VPWR _17020_/X sky130_fd_sc_hd__buf_2
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _14635_/A _14230_/X _14231_/X VGND VGND VPWR VPWR _14232_/X sky130_fd_sc_hd__and3_4
XANTENNA__21248__A2 _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23265__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14163_ _13791_/A _14161_/X _14163_/C VGND VGND VPWR VPWR _14164_/C sky130_fd_sc_hd__and3_4
XANTENNA__17321__B1 _12882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13114_ _13090_/A _13114_/B _13114_/C VGND VGND VPWR VPWR _13114_/X sky130_fd_sc_hd__and3_4
XANTENNA__15907__B _15837_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18971_ _18948_/A _18948_/B _18964_/A VGND VGND VPWR VPWR _18971_/X sky130_fd_sc_hd__o21a_4
X_14094_ _14094_/A VGND VGND VPWR VPWR _14103_/A sky130_fd_sc_hd__buf_2
XFILLER_4_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20208__B1 _20200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22748__A2 _22736_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13045_ _13045_/A _13045_/B _13045_/C VGND VGND VPWR VPWR _13045_/X sky130_fd_sc_hd__or3_4
XFILLER_26_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17922_ _17922_/A VGND VGND VPWR VPWR _17922_/X sky130_fd_sc_hd__buf_2
XFILLER_105_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17853_ _17922_/A _17851_/X _17836_/X _17852_/X VGND VGND VPWR VPWR _17854_/A sky130_fd_sc_hd__o22a_4
X_16804_ _16811_/A _23825_/Q VGND VGND VPWR VPWR _16804_/X sky130_fd_sc_hd__or2_4
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17784_ _17655_/X _17782_/Y _17783_/X VGND VGND VPWR VPWR _17784_/X sky130_fd_sc_hd__o21a_4
X_14996_ _13952_/A _24021_/Q VGND VGND VPWR VPWR _14998_/B sky130_fd_sc_hd__or2_4
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19523_ _19499_/A VGND VGND VPWR VPWR _19524_/A sky130_fd_sc_hd__inv_2
XFILLER_47_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13947_ _13946_/Y VGND VGND VPWR VPWR _13947_/X sky130_fd_sc_hd__buf_2
X_16735_ _12059_/X _24113_/Q VGND VGND VPWR VPWR _16736_/C sky130_fd_sc_hd__or2_4
XANTENNA__17388__B1 _17358_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13443__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19454_ _19454_/A VGND VGND VPWR VPWR _19454_/X sky130_fd_sc_hd__buf_2
X_16666_ _16678_/A _16664_/X _16666_/C VGND VGND VPWR VPWR _16666_/X sky130_fd_sc_hd__and3_4
XANTENNA__20931__A1 _18681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13878_ _14377_/A _23741_/Q VGND VGND VPWR VPWR _13879_/C sky130_fd_sc_hd__or2_4
XANTENNA__21660__A _21667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18405_ _18405_/A _17387_/A VGND VGND VPWR VPWR _18405_/X sky130_fd_sc_hd__or2_4
X_15617_ _13928_/A _15609_/X _15617_/C VGND VGND VPWR VPWR _15618_/C sky130_fd_sc_hd__and3_4
XANTENNA__13162__B _23975_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12829_ _12829_/A VGND VGND VPWR VPWR _13370_/A sky130_fd_sc_hd__buf_2
X_16597_ _16594_/A _23890_/Q VGND VGND VPWR VPWR _16597_/X sky130_fd_sc_hd__or2_4
X_19385_ _19383_/X VGND VGND VPWR VPWR _19385_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16754__A _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12059__A _11990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21487__A2 _21485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18336_ _18282_/A _18336_/B VGND VGND VPWR VPWR _18337_/D sky130_fd_sc_hd__and2_4
X_15548_ _12427_/A _15548_/B _15547_/X VGND VGND VPWR VPWR _15548_/X sky130_fd_sc_hd__and3_4
XFILLER_148_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22906__D _19910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20144__C1 _20192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22684__B2 _22648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23608__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11898__A _11898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18267_ _18168_/A _18266_/X VGND VGND VPWR VPWR _18267_/Y sky130_fd_sc_hd__nor2_4
XFILLER_72_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15479_ _12650_/A _15479_/B _15478_/X VGND VGND VPWR VPWR _15479_/X sky130_fd_sc_hd__and3_4
XANTENNA__14274__A _12454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17218_ _17137_/X _17210_/X _17112_/X _17217_/X VGND VGND VPWR VPWR _17218_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22436__B2 _22433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19784__B HRDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18198_ _18198_/A VGND VGND VPWR VPWR _18198_/X sky130_fd_sc_hd__buf_2
XANTENNA__15089__B _24053_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22491__A _22498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17585__A _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17149_ _17128_/X _17142_/X _17113_/X _17148_/X VGND VGND VPWR VPWR _17149_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20160_ IRQ[15] VGND VGND VPWR VPWR _20160_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14721__B _14721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13618__A _15395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20091_ _20091_/A VGND VGND VPWR VPWR _20091_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12522__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21411__A2 _21405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16929__A _16927_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23850_ _23531_/CLK _23850_/D VGND VGND VPWR VPWR _12817_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_38_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22801_ _18738_/X _22800_/Y _16918_/X VGND VGND VPWR VPWR _22801_/X sky130_fd_sc_hd__o21a_4
X_23781_ _23493_/CLK _23781_/D VGND VGND VPWR VPWR _23781_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14449__A _14310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20993_ _20490_/A _20992_/Y _24278_/Q _20347_/X VGND VGND VPWR VPWR _20993_/X sky130_fd_sc_hd__o22a_4
XFILLER_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21175__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22732_ _20959_/A _22729_/X _15304_/B _22726_/X VGND VGND VPWR VPWR _23096_/D sky130_fd_sc_hd__o22a_4
XFILLER_164_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22663_ _22444_/X _22658_/X _13316_/B _22662_/X VGND VGND VPWR VPWR _22663_/X sky130_fd_sc_hd__o22a_4
XFILLER_129_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24402_ _23281_/CLK _18903_/X HRESETn VGND VGND VPWR VPWR _24402_/Q sky130_fd_sc_hd__dfstp_4
X_21614_ _21528_/X _21613_/X _23763_/Q _21610_/X VGND VGND VPWR VPWR _23763_/D sky130_fd_sc_hd__o22a_4
X_22594_ _22608_/A VGND VGND VPWR VPWR _22594_/X sky130_fd_sc_hd__buf_2
XANTENNA__22675__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20686__B1 _20538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24333_ _24294_/CLK _19176_/X HRESETn VGND VGND VPWR VPWR _19154_/A sky130_fd_sc_hd__dfrtp_4
X_21545_ _21544_/X _21542_/X _16178_/B _21537_/X VGND VGND VPWR VPWR _21545_/X sky130_fd_sc_hd__o22a_4
XFILLER_21_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11601__A _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22427__B2 _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24264_ _24271_/CLK _19352_/X HRESETn VGND VGND VPWR VPWR _20570_/A sky130_fd_sc_hd__dfrtp_4
X_21476_ _21469_/Y _21475_/X _21241_/X _21475_/X VGND VGND VPWR VPWR _23828_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_14_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20914__A _22158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23215_ _23760_/CLK _23215_/D VGND VGND VPWR VPWR _16256_/B sky130_fd_sc_hd__dfxtp_4
X_20427_ _20427_/A VGND VGND VPWR VPWR _20427_/X sky130_fd_sc_hd__buf_2
X_24195_ _23511_/CLK _19814_/X HRESETn VGND VGND VPWR VPWR _11706_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14912__A _11659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23146_ _23531_/CLK _23146_/D VGND VGND VPWR VPWR _12816_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15727__B _23780_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20358_ _20358_/A _20357_/X VGND VGND VPWR VPWR _20358_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21650__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23077_ _23076_/X VGND VGND VPWR VPWR HADDR[30] sky130_fd_sc_hd__inv_2
X_20289_ _20315_/A VGND VGND VPWR VPWR _20344_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_2_0_HCLK_A clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13340__A1 _13453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21745__A _21724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22028_ _22007_/A VGND VGND VPWR VPWR _22028_/X sky130_fd_sc_hd__buf_2
XFILLER_48_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15743__A _13205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14850_ _12218_/A _14850_/B VGND VGND VPWR VPWR _14850_/X sky130_fd_sc_hd__or2_4
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13801_ _15394_/A _13801_/B _13801_/C VGND VGND VPWR VPWR _13801_/X sky130_fd_sc_hd__and3_4
XFILLER_21_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24384__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15462__B _15399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14781_ _14667_/A _14781_/B _14781_/C VGND VGND VPWR VPWR _14782_/C sky130_fd_sc_hd__and3_4
X_23979_ _23558_/CLK _21203_/X VGND VGND VPWR VPWR _23979_/Q sky130_fd_sc_hd__dfxtp_4
X_11993_ _16744_/A _11824_/B VGND VGND VPWR VPWR _11993_/X sky130_fd_sc_hd__or2_4
X_16520_ _11815_/X _16504_/X _16519_/X VGND VGND VPWR VPWR _16520_/X sky130_fd_sc_hd__or3_4
XANTENNA__13263__A _13262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13732_ _15486_/A _13732_/B VGND VGND VPWR VPWR _13732_/X sky130_fd_sc_hd__or2_4
XFILLER_43_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_40_0_HCLK clkbuf_5_20_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_40_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14078__B _23232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16451_ _11858_/A _11631_/X _16420_/X _11608_/A _16450_/X VGND VGND VPWR VPWR _16451_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13663_ _13663_/A VGND VGND VPWR VPWR _14331_/A sky130_fd_sc_hd__buf_2
X_15402_ _15402_/A _15465_/B VGND VGND VPWR VPWR _15404_/B sky130_fd_sc_hd__or2_4
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12614_ _12977_/A _12595_/X _12614_/C VGND VGND VPWR VPWR _12614_/X sky130_fd_sc_hd__and3_4
X_19170_ _24336_/Q _19157_/B _19169_/Y VGND VGND VPWR VPWR _19170_/X sky130_fd_sc_hd__o21a_4
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16382_ _16381_/X VGND VGND VPWR VPWR _16383_/A sky130_fd_sc_hd__inv_2
XANTENNA__22666__B2 _22662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20096__A _11635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13594_ _13974_/A VGND VGND VPWR VPWR _13983_/A sky130_fd_sc_hd__buf_2
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18121_ _17878_/X _17928_/X _17823_/X _17937_/X VGND VGND VPWR VPWR _18122_/A sky130_fd_sc_hd__o22a_4
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15333_ _15328_/A _15333_/B VGND VGND VPWR VPWR _15333_/X sky130_fd_sc_hd__or2_4
X_12545_ _15449_/A VGND VGND VPWR VPWR _12546_/A sky130_fd_sc_hd__buf_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12607__A _12623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18052_ _17810_/X _17855_/X _17880_/A VGND VGND VPWR VPWR _18052_/X sky130_fd_sc_hd__o21a_4
X_15264_ _14148_/A _15264_/B VGND VGND VPWR VPWR _15264_/X sky130_fd_sc_hd__or2_4
X_12476_ _14325_/A VGND VGND VPWR VPWR _12477_/A sky130_fd_sc_hd__buf_2
X_17003_ _17727_/A VGND VGND VPWR VPWR _17006_/A sky130_fd_sc_hd__buf_2
X_14215_ _13868_/A VGND VGND VPWR VPWR _14240_/A sky130_fd_sc_hd__buf_2
X_15195_ _14786_/A _15195_/B _15195_/C VGND VGND VPWR VPWR _15201_/B sky130_fd_sc_hd__and3_4
XFILLER_126_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14146_ _14003_/A _14144_/X _14146_/C VGND VGND VPWR VPWR _14150_/B sky130_fd_sc_hd__and3_4
XFILLER_99_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14541__B _14469_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13438__A _13474_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18954_ _18949_/A _18949_/B _18950_/Y _18953_/X VGND VGND VPWR VPWR _18955_/A sky130_fd_sc_hd__o22a_4
X_14077_ _11736_/A _14075_/X _14077_/C VGND VGND VPWR VPWR _14081_/B sky130_fd_sc_hd__and3_4
X_13028_ _12510_/A _13028_/B VGND VGND VPWR VPWR _13028_/X sky130_fd_sc_hd__or2_4
XFILLER_117_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17905_ _17905_/A VGND VGND VPWR VPWR _17906_/A sky130_fd_sc_hd__buf_2
X_18885_ _16866_/X _18840_/A _24405_/Q _18843_/A VGND VGND VPWR VPWR _18885_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20601__B1 _20157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17836_ _17836_/A VGND VGND VPWR VPWR _17836_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_122_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR _23241_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17767_ _17767_/A _17714_/X _17767_/C VGND VGND VPWR VPWR _17768_/C sky130_fd_sc_hd__or3_4
XANTENNA__21157__B2 _21152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14979_ _14783_/X _14975_/X _14979_/C VGND VGND VPWR VPWR _14979_/X sky130_fd_sc_hd__or3_4
XANTENNA__14269__A _14269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13173__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19506_ _19506_/A VGND VGND VPWR VPWR _19507_/B sky130_fd_sc_hd__inv_2
X_16718_ _11973_/X _16718_/B VGND VGND VPWR VPWR _16718_/X sky130_fd_sc_hd__and2_4
X_17698_ _17698_/A _17689_/X _17698_/C VGND VGND VPWR VPWR _17698_/X sky130_fd_sc_hd__and3_4
XANTENNA__19770__A1 _19519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19437_ _24128_/Q VGND VGND VPWR VPWR _19438_/B sky130_fd_sc_hd__buf_2
X_16649_ _16677_/A _23570_/Q VGND VGND VPWR VPWR _16649_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_4_13_0_HCLK_A clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13901__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16915__C _16915_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22657__B2 _22655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19368_ _19365_/X _18592_/X _19365_/X _24253_/Q VGND VGND VPWR VPWR _19368_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14716__B _14716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18319_ _18131_/X _17865_/X _18053_/X VGND VGND VPWR VPWR _18319_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__12517__A _12878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19299_ _19237_/B VGND VGND VPWR VPWR _19299_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21330_ _21249_/X _21327_/X _23921_/Q _21324_/X VGND VGND VPWR VPWR _23921_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21880__A2 _21875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21261_ _20486_/A VGND VGND VPWR VPWR _21261_/X sky130_fd_sc_hd__buf_2
XANTENNA__18204__A _18320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23000_ _19438_/A VGND VGND VPWR VPWR _23043_/A sky130_fd_sc_hd__buf_2
XFILLER_150_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20212_ _24129_/Q VGND VGND VPWR VPWR _20218_/A sky130_fd_sc_hd__inv_2
XANTENNA__21632__A2 _21627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21192_ _20337_/X _21191_/X _23987_/Q _21188_/X VGND VGND VPWR VPWR _23987_/D sky130_fd_sc_hd__o22a_4
XFILLER_132_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20143_ _11576_/X _20141_/X _20142_/Y VGND VGND VPWR VPWR _20143_/Y sky130_fd_sc_hd__o21ai_4
X_20074_ _20074_/A VGND VGND VPWR VPWR _20074_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21396__B2 _21395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16659__A _16659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23902_ _23518_/CLK _21357_/X VGND VGND VPWR VPWR _13750_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24086__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23833_ _23641_/CLK _21464_/X VGND VGND VPWR VPWR _14744_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13083__A _13100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23764_ _23764_/CLK _21611_/X VGND VGND VPWR VPWR _23764_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22896__A1 _16687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _20305_/X _20967_/Y _20974_/X _20975_/Y _20255_/A VGND VGND VPWR VPWR _20976_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_27_0_HCLK clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22715_ _22708_/A VGND VGND VPWR VPWR _22715_/X sky130_fd_sc_hd__buf_2
XPHY_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16394__A _16007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23695_ _23662_/CLK _21719_/X VGND VGND VPWR VPWR _16338_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_80_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14907__A _13955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13811__A _13656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22646_ _22416_/X _22644_/X _16661_/B _22641_/X VGND VGND VPWR VPWR _23154_/D sky130_fd_sc_hd__o22a_4
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22577_ _22468_/X _22572_/X _14349_/B _22576_/X VGND VGND VPWR VPWR _23196_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12427__A _12427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22843__B _17273_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12330_ _12625_/A VGND VGND VPWR VPWR _13205_/A sky130_fd_sc_hd__buf_2
X_24316_ _24292_/CLK _24316_/D HRESETn VGND VGND VPWR VPWR _19137_/A sky130_fd_sc_hd__dfrtp_4
X_21528_ _21528_/A VGND VGND VPWR VPWR _21528_/X sky130_fd_sc_hd__buf_2
XFILLER_139_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21871__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23020__A _22949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12261_ _12266_/A _12261_/B _12260_/X VGND VGND VPWR VPWR _12261_/X sky130_fd_sc_hd__or3_4
XANTENNA__15738__A _15778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24247_ _23126_/CLK _19379_/X HRESETn VGND VGND VPWR VPWR _24247_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21459_ _21438_/A VGND VGND VPWR VPWR _21459_/X sky130_fd_sc_hd__buf_2
XANTENNA__14642__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14000_ _11618_/A VGND VGND VPWR VPWR _14003_/A sky130_fd_sc_hd__buf_2
XFILLER_108_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21623__A2 _21620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12192_ _13042_/A VGND VGND VPWR VPWR _12568_/A sky130_fd_sc_hd__buf_2
X_24178_ _23383_/CLK _19927_/X HRESETn VGND VGND VPWR VPWR _24178_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17953__A _18413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23129_ _23641_/CLK _22681_/X VGND VGND VPWR VPWR _14743_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_150_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21475__A _21482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15951_ _15982_/A _23790_/Q VGND VGND VPWR VPWR _15952_/C sky130_fd_sc_hd__or2_4
XFILLER_114_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21387__B2 _21381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16569__A _11973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14902_ _14905_/A _14902_/B VGND VGND VPWR VPWR _14902_/X sky130_fd_sc_hd__or2_4
X_15882_ _13532_/A _15820_/B VGND VGND VPWR VPWR _15883_/C sky130_fd_sc_hd__or2_4
X_18670_ _18670_/A VGND VGND VPWR VPWR _18670_/X sky130_fd_sc_hd__buf_2
XFILLER_48_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17621_ _17308_/X _17621_/B _17620_/X VGND VGND VPWR VPWR _17621_/X sky130_fd_sc_hd__and3_4
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14833_ _14660_/A _14833_/B _14832_/X VGND VGND VPWR VPWR _14833_/X sky130_fd_sc_hd__or3_4
XANTENNA__21139__B2 _21138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14089__A _11623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18784__A _18837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22887__A1 _17556_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17552_ _17642_/A VGND VGND VPWR VPWR _17971_/B sky130_fd_sc_hd__inv_2
X_14764_ _13853_/A _14763_/X VGND VGND VPWR VPWR _14764_/X sky130_fd_sc_hd__and2_4
X_11976_ _12012_/A _23604_/Q VGND VGND VPWR VPWR _11977_/C sky130_fd_sc_hd__or2_4
XANTENNA__16015__B1 _11608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20819__A _20819_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16503_ _16362_/X _16499_/X _16502_/X VGND VGND VPWR VPWR _16504_/C sky130_fd_sc_hd__or3_4
X_13715_ _14372_/A _13708_/X _13714_/X VGND VGND VPWR VPWR _13715_/X sky130_fd_sc_hd__or3_4
XANTENNA__20898__B1 HRDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22737__C _20598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17483_ _17482_/X VGND VGND VPWR VPWR _17483_/Y sky130_fd_sc_hd__inv_2
X_14695_ _15620_/A _14601_/B VGND VGND VPWR VPWR _14696_/C sky130_fd_sc_hd__or2_4
X_19222_ _24310_/Q _19131_/B _19221_/Y VGND VGND VPWR VPWR _19222_/X sky130_fd_sc_hd__o21a_4
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16434_ _15934_/X _16434_/B _16433_/X VGND VGND VPWR VPWR _16434_/X sky130_fd_sc_hd__or3_4
X_13646_ _13628_/A _13736_/B VGND VGND VPWR VPWR _13646_/X sky130_fd_sc_hd__or2_4
XFILLER_20_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16365_ _16313_/A _16363_/X _16364_/X VGND VGND VPWR VPWR _16365_/X sky130_fd_sc_hd__and3_4
XFILLER_13_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19153_ _19153_/A _19153_/B VGND VGND VPWR VPWR _19154_/B sky130_fd_sc_hd__and2_4
XFILLER_82_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20114__A2 _20113_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13577_ _12846_/A _12984_/Y _12845_/A VGND VGND VPWR VPWR _13578_/B sky130_fd_sc_hd__o21ai_4
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18104_ _17673_/X _18103_/X _17673_/X _18103_/X VGND VGND VPWR VPWR _18104_/X sky130_fd_sc_hd__a2bb2o_4
X_15316_ _15319_/A _23512_/Q VGND VGND VPWR VPWR _15317_/C sky130_fd_sc_hd__or2_4
XFILLER_160_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12528_ _15000_/A VGND VGND VPWR VPWR _14295_/A sky130_fd_sc_hd__buf_2
X_16296_ _15944_/A _16296_/B VGND VGND VPWR VPWR _16296_/X sky130_fd_sc_hd__or2_4
X_19084_ _24382_/Q VGND VGND VPWR VPWR _19084_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_47_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR _24077_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18035_ _18310_/A _18035_/B VGND VGND VPWR VPWR _18035_/X sky130_fd_sc_hd__or2_4
X_15247_ _13882_/A _15247_/B _15247_/C VGND VGND VPWR VPWR _15248_/C sky130_fd_sc_hd__or3_4
XANTENNA__15648__A _13894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12459_ _12857_/A _12440_/X _12459_/C VGND VGND VPWR VPWR _12459_/X sky130_fd_sc_hd__or3_4
XFILLER_172_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23064__B2 _22930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21075__B1 _24057_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17818__A1 _17816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21614__A2 _21613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15178_ _13954_/A _15176_/X _15178_/C VGND VGND VPWR VPWR _15178_/X sky130_fd_sc_hd__and3_4
XANTENNA__13168__A _13164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14129_ _14094_/A _14129_/B _14129_/C VGND VGND VPWR VPWR _14129_/X sky130_fd_sc_hd__and3_4
XANTENNA__24120__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19986_ _18670_/X _16945_/X _19956_/X _19985_/X VGND VGND VPWR VPWR _19987_/A sky130_fd_sc_hd__o22a_4
XANTENNA__12072__A _11990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18937_ _17290_/X _18934_/X _24378_/Q _18935_/X VGND VGND VPWR VPWR _18937_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16479__A _13384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21378__B2 _21374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22575__B1 _13807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12800__A _12800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18868_ _17169_/X _18863_/X _24418_/Q _18864_/X VGND VGND VPWR VPWR _24418_/D sky130_fd_sc_hd__o22a_4
X_17819_ _17825_/A VGND VGND VPWR VPWR _17819_/X sky130_fd_sc_hd__buf_2
XFILLER_82_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18799_ _17139_/X _18796_/X _24462_/Q _18797_/X VGND VGND VPWR VPWR _24462_/D sky130_fd_sc_hd__o22a_4
X_20830_ _20726_/X _20829_/Y _19234_/A _20347_/X VGND VGND VPWR VPWR _20830_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20761_ _20761_/A VGND VGND VPWR VPWR _20761_/X sky130_fd_sc_hd__buf_2
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21550__B2 _21549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14727__A _13990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22500_ _22423_/X _22494_/X _16296_/B _22498_/X VGND VGND VPWR VPWR _23247_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13631__A _14329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23480_ _23098_/CLK _22084_/X VGND VGND VPWR VPWR _23480_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20692_ _20692_/A VGND VGND VPWR VPWR _21283_/A sky130_fd_sc_hd__buf_2
XFILLER_11_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14446__B _14502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22431_ _22430_/X _22426_/X _12193_/B _22421_/X VGND VGND VPWR VPWR _22431_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16309__A1 _11858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16309__B2 _16308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16942__A _16941_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22362_ _22376_/A VGND VGND VPWR VPWR _22362_/X sky130_fd_sc_hd__buf_2
XANTENNA__24279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24101_ _23493_/CLK _20634_/X VGND VGND VPWR VPWR _13470_/B sky130_fd_sc_hd__dfxtp_4
X_21313_ _21313_/A VGND VGND VPWR VPWR _21313_/X sky130_fd_sc_hd__buf_2
XANTENNA__15558__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14462__A _12537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22293_ _22120_/X _22287_/X _12768_/B _22291_/X VGND VGND VPWR VPWR _22293_/X sky130_fd_sc_hd__o22a_4
XFILLER_163_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24032_ _23523_/CLK _24032_/D VGND VGND VPWR VPWR _24032_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15277__B _23160_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21244_ _21238_/A VGND VGND VPWR VPWR _21269_/A sky130_fd_sc_hd__buf_2
XFILLER_172_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14181__B _23263_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_4_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13078__A _13067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21175_ _20892_/X _21169_/X _23995_/Q _21173_/X VGND VGND VPWR VPWR _21175_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21295__A _20819_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20126_ _20119_/Y _20123_/Y _11583_/X _20125_/X VGND VGND VPWR VPWR _20126_/X sky130_fd_sc_hd__a211o_4
XANTENNA__23476__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15293__A _14267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20057_ _18430_/X _20055_/X _20056_/Y _20042_/X VGND VGND VPWR VPWR _20057_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13806__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19431__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22030__A2 _22024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20592__A2 _20443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23816_ _23592_/CLK _21494_/X VGND VGND VPWR VPWR _13110_/B sky130_fd_sc_hd__dfxtp_4
X_11830_ _12169_/A _11826_/X _11829_/X VGND VGND VPWR VPWR _11830_/X sky130_fd_sc_hd__or3_4
XANTENNA__22869__A1 _14483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23015__A _18299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23747_ _23111_/CLK _23747_/D VGND VGND VPWR VPWR _15854_/B sky130_fd_sc_hd__dfxtp_4
X_11761_ _11760_/X VGND VGND VPWR VPWR _12138_/A sky130_fd_sc_hd__buf_2
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ _20959_/A VGND VGND VPWR VPWR _20959_/X sky130_fd_sc_hd__buf_2
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14637__A _14677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13531_/A _13500_/B VGND VGND VPWR VPWR _13500_/X sky130_fd_sc_hd__or2_4
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14480_/A _14479_/X VGND VGND VPWR VPWR _14480_/X sky130_fd_sc_hd__and2_4
XFILLER_14_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11692_ _13407_/A VGND VGND VPWR VPWR _16205_/A sky130_fd_sc_hd__buf_2
XPHY_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23678_ _23678_/CLK _21743_/X VGND VGND VPWR VPWR _13741_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _12864_/A VGND VGND VPWR VPWR _13431_/X sky130_fd_sc_hd__buf_2
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22629_ _22622_/A VGND VGND VPWR VPWR _22629_/X sky130_fd_sc_hd__buf_2
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19498__B1 HRDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12157__A _11705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16150_ _16147_/A _16150_/B VGND VGND VPWR VPWR _16150_/X sky130_fd_sc_hd__or2_4
X_13362_ _13392_/A _13358_/X _13362_/C VGND VGND VPWR VPWR _13363_/C sky130_fd_sc_hd__or3_4
XFILLER_155_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21844__A2 _21839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15101_ _15096_/A _15038_/B VGND VGND VPWR VPWR _15101_/X sky130_fd_sc_hd__or2_4
X_12313_ _13183_/A _23724_/Q VGND VGND VPWR VPWR _12315_/B sky130_fd_sc_hd__or2_4
X_16081_ _16035_/A _16081_/B _16081_/C VGND VGND VPWR VPWR _16081_/X sky130_fd_sc_hd__and3_4
X_13293_ _13304_/A VGND VGND VPWR VPWR _13320_/A sky130_fd_sc_hd__buf_2
XFILLER_155_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24251__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15032_ _11912_/A _15030_/X _15031_/X VGND VGND VPWR VPWR _15036_/B sky130_fd_sc_hd__and3_4
X_12244_ _12311_/A VGND VGND VPWR VPWR _13301_/A sky130_fd_sc_hd__buf_2
XFILLER_108_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14091__B _23519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19840_ _19752_/B VGND VGND VPWR VPWR _19868_/B sky130_fd_sc_hd__buf_2
X_12175_ _11834_/A _12173_/X _12175_/C VGND VGND VPWR VPWR _12175_/X sky130_fd_sc_hd__and3_4
XANTENNA__18473__B2 _18472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19771_ _19576_/X _19762_/X _19768_/Y _19603_/X _19770_/Y VGND VGND VPWR VPWR _19771_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_110_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16983_ _16983_/A _18433_/A VGND VGND VPWR VPWR _18403_/B sky130_fd_sc_hd__or2_4
XFILLER_27_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13716__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18722_ _17329_/X VGND VGND VPWR VPWR _18722_/Y sky130_fd_sc_hd__inv_2
X_15934_ _12516_/A VGND VGND VPWR VPWR _15934_/X sky130_fd_sc_hd__buf_2
XFILLER_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18653_ _17249_/X _18653_/B VGND VGND VPWR VPWR _18653_/X sky130_fd_sc_hd__and2_4
XFILLER_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15865_ _13539_/A _15865_/B VGND VGND VPWR VPWR _15865_/X sky130_fd_sc_hd__or2_4
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17984__B1 _17813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21780__B2 _21774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17604_ _17639_/A _17603_/X VGND VGND VPWR VPWR _17640_/C sky130_fd_sc_hd__or2_4
X_14816_ _14823_/A _24057_/Q VGND VGND VPWR VPWR _14817_/C sky130_fd_sc_hd__or2_4
XFILLER_91_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18584_ _18168_/A _18161_/X VGND VGND VPWR VPWR _18584_/Y sky130_fd_sc_hd__nor2_4
X_15796_ _11888_/A _15796_/B VGND VGND VPWR VPWR _15796_/X sky130_fd_sc_hd__or2_4
XANTENNA__20549__A _20264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17535_ _17165_/Y _18280_/B _17517_/Y _17534_/X VGND VGND VPWR VPWR _17535_/X sky130_fd_sc_hd__o22a_4
X_11959_ _11891_/X VGND VGND VPWR VPWR _11960_/A sky130_fd_sc_hd__buf_2
X_14747_ _14329_/A _23417_/Q VGND VGND VPWR VPWR _14748_/C sky130_fd_sc_hd__or2_4
XANTENNA__14547__A _15517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20335__A2 _20304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13451__A _12869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_10_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17466_ _17156_/A _17467_/B VGND VGND VPWR VPWR _17469_/A sky130_fd_sc_hd__and2_4
X_14678_ _14691_/A _23386_/Q VGND VGND VPWR VPWR _14680_/B sky130_fd_sc_hd__or2_4
X_19205_ _19205_/A VGND VGND VPWR VPWR _19205_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16417_ _11882_/X _16415_/X _16416_/X VGND VGND VPWR VPWR _16417_/X sky130_fd_sc_hd__and3_4
X_13629_ _13658_/A _13741_/B VGND VGND VPWR VPWR _13629_/X sky130_fd_sc_hd__or2_4
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17397_ _13863_/X VGND VGND VPWR VPWR _17397_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19136_ _19136_/A _19213_/A VGND VGND VPWR VPWR _19211_/A sky130_fd_sc_hd__and2_4
XFILLER_34_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21835__A2 _21827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16348_ _16195_/A _16280_/B VGND VGND VPWR VPWR _16348_/X sky130_fd_sc_hd__or2_4
XFILLER_121_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16279_ _16282_/A _16279_/B VGND VGND VPWR VPWR _16279_/X sky130_fd_sc_hd__or2_4
XANTENNA__24301__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19067_ _19046_/X _19065_/X _19066_/Y _19049_/X VGND VGND VPWR VPWR _19067_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14282__A _13601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21048__B1 _24076_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18018_ _17900_/X _18017_/X _19999_/A _17900_/X VGND VGND VPWR VPWR _24496_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12514__B _12514_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21599__B2 _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22260__A2 _22258_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19969_ _17807_/X _18753_/Y _17870_/X _19968_/Y VGND VGND VPWR VPWR _19969_/X sky130_fd_sc_hd__a211o_4
XFILLER_80_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22012__A2 _22010_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13626__A _15405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12530__A _12530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22980_ _18472_/X _22973_/B VGND VGND VPWR VPWR _22981_/C sky130_fd_sc_hd__or2_4
XANTENNA__16002__A _16110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22939__A _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21220__B1 _23967_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21931_ _21874_/X _21930_/X _14645_/B _21927_/X VGND VGND VPWR VPWR _23578_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21771__B2 _21767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15841__A _12487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21862_ _20801_/A VGND VGND VPWR VPWR _21862_/X sky130_fd_sc_hd__buf_2
X_23601_ _23761_/CLK _23601_/D VGND VGND VPWR VPWR _23601_/Q sky130_fd_sc_hd__dfxtp_4
X_20813_ _18568_/X _20702_/X _20753_/X _20812_/Y VGND VGND VPWR VPWR _20813_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24124__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14457__A _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21793_ _21580_/X _21791_/X _13776_/B _21788_/X VGND VGND VPWR VPWR _23646_/D sky130_fd_sc_hd__o22a_4
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23532_ _23500_/CLK _23532_/D VGND VGND VPWR VPWR _23532_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20744_ _20744_/A VGND VGND VPWR VPWR _20745_/A sky130_fd_sc_hd__buf_2
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22079__A2 _22074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23463_ _23303_/CLK _23463_/D VGND VGND VPWR VPWR _13217_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20675_ _20259_/A VGND VGND VPWR VPWR _20675_/X sky130_fd_sc_hd__buf_2
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16672__A _16672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22414_ _22438_/A VGND VGND VPWR VPWR _22414_/X sky130_fd_sc_hd__buf_2
X_23394_ _23523_/CLK _23394_/D VGND VGND VPWR VPWR _15432_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_52_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22345_ _13818_/B VGND VGND VPWR VPWR _23325_/D sky130_fd_sc_hd__buf_2
XANTENNA__19983__A _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14192__A _14615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12705__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_30_0_HCLK clkbuf_7_31_0_HCLK/A VGND VGND VPWR VPWR _23281_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_151_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22276_ _22291_/A VGND VGND VPWR VPWR _22284_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_93_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR _24057_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_151_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24015_ _23983_/CLK _24015_/D VGND VGND VPWR VPWR _16339_/B sky130_fd_sc_hd__dfxtp_4
X_21227_ _20915_/X _21226_/X _14584_/B _21223_/X VGND VGND VPWR VPWR _21227_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21158_ _20596_/X _21155_/X _24007_/Q _21152_/X VGND VGND VPWR VPWR _21158_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18111__B _18148_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20109_ _11574_/X VGND VGND VPWR VPWR _20109_/Y sky130_fd_sc_hd__inv_2
X_13980_ _11930_/A _13976_/X _13980_/C VGND VGND VPWR VPWR _13980_/X sky130_fd_sc_hd__or3_4
X_21089_ _21118_/A VGND VGND VPWR VPWR _21104_/A sky130_fd_sc_hd__buf_2
XANTENNA__20014__A1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12931_ _12977_/A _12921_/X _12930_/X VGND VGND VPWR VPWR _12947_/B sky130_fd_sc_hd__and3_4
XFILLER_150_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15751__A _12641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12862_ _12862_/A VGND VGND VPWR VPWR _12889_/A sky130_fd_sc_hd__buf_2
X_15650_ _11668_/A _15618_/X _15649_/X VGND VGND VPWR VPWR _15651_/A sky130_fd_sc_hd__and3_4
XFILLER_74_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11813_ _11813_/A VGND VGND VPWR VPWR _12978_/A sky130_fd_sc_hd__buf_2
X_14601_ _13632_/A _14601_/B VGND VGND VPWR VPWR _14601_/X sky130_fd_sc_hd__or2_4
XANTENNA__15470__B _15470_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15581_ _11969_/A _15558_/X _15565_/X _15572_/X _15580_/X VGND VGND VPWR VPWR _15581_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12793_ _15770_/A VGND VGND VPWR VPWR _12833_/A sky130_fd_sc_hd__buf_2
XANTENNA__21514__A1 _21304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21514__B2 _21510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14520_/A _14474_/B VGND VGND VPWR VPWR _14532_/X sky130_fd_sc_hd__or2_4
X_17320_ _21028_/A VGND VGND VPWR VPWR _19852_/A sky130_fd_sc_hd__inv_2
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11744_ _16079_/A VGND VGND VPWR VPWR _12151_/A sky130_fd_sc_hd__buf_2
XANTENNA__17194__A1 _16383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18391__B1 _18320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14086__B _14084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14463_ _13010_/A _14463_/B VGND VGND VPWR VPWR _14464_/C sky130_fd_sc_hd__or2_4
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _17251_/A _17251_/B VGND VGND VPWR VPWR _17251_/X sky130_fd_sc_hd__and2_4
X_11675_ _11675_/A VGND VGND VPWR VPWR _12641_/A sky130_fd_sc_hd__buf_2
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16202_ _16202_/A _23341_/Q VGND VGND VPWR VPWR _16202_/X sky130_fd_sc_hd__or2_4
X_13414_ _13414_/A _13414_/B _13414_/C VGND VGND VPWR VPWR _13415_/C sky130_fd_sc_hd__or3_4
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17182_ _12027_/X VGND VGND VPWR VPWR _17847_/A sky130_fd_sc_hd__buf_2
X_14394_ _14513_/A _14389_/X _14393_/X VGND VGND VPWR VPWR _14394_/X sky130_fd_sc_hd__or3_4
XFILLER_155_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16133_ _16109_/A _23981_/Q VGND VGND VPWR VPWR _16134_/C sky130_fd_sc_hd__or2_4
X_13345_ _13384_/A _13273_/B VGND VGND VPWR VPWR _13345_/X sky130_fd_sc_hd__or2_4
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12615__A _11781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16064_ _16057_/A _23406_/Q VGND VGND VPWR VPWR _16064_/X sky130_fd_sc_hd__or2_4
X_13276_ _13276_/A VGND VGND VPWR VPWR _13321_/A sky130_fd_sc_hd__buf_2
XFILLER_170_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15015_ _14012_/A _14991_/X _14999_/X _15006_/X _15014_/X VGND VGND VPWR VPWR _15015_/X
+ sky130_fd_sc_hd__a32o_4
X_12227_ _11880_/A VGND VGND VPWR VPWR _12704_/A sky130_fd_sc_hd__buf_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22242__A2 _22237_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19823_ _19823_/A _19823_/B VGND VGND VPWR VPWR _19823_/X sky130_fd_sc_hd__or2_4
XFILLER_110_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12158_ _12151_/A _12158_/B VGND VGND VPWR VPWR _12158_/X sky130_fd_sc_hd__or2_4
XFILLER_64_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13446__A _12863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19754_ _19705_/A _19665_/B _19659_/Y _19879_/C VGND VGND VPWR VPWR _19754_/X sky130_fd_sc_hd__and4_4
XFILLER_110_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16966_ _24140_/Q VGND VGND VPWR VPWR _17726_/A sky130_fd_sc_hd__inv_2
X_12089_ _12058_/A _12158_/B VGND VGND VPWR VPWR _12089_/X sky130_fd_sc_hd__or2_4
XANTENNA__20005__A1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21663__A _21677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18705_ _16933_/Y _18700_/X _16933_/Y _18704_/X VGND VGND VPWR VPWR _18705_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24147__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15917_ _15915_/Y _15916_/X VGND VGND VPWR VPWR _15917_/X sky130_fd_sc_hd__or2_4
X_19685_ _19684_/X VGND VGND VPWR VPWR _19685_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13691__B1 _11606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16897_ _16829_/X _16897_/B _16838_/X _16897_/D VGND VGND VPWR VPWR _16898_/B sky130_fd_sc_hd__and4_4
XANTENNA__16757__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21753__B2 _21717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15661__A _12690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18636_ _17351_/B _18634_/X VGND VGND VPWR VPWR _18636_/Y sky130_fd_sc_hd__nand2_4
X_15848_ _13307_/A _15825_/X _15832_/X _15839_/X _15847_/X VGND VGND VPWR VPWR _15848_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_91_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18567_ _18567_/A VGND VGND VPWR VPWR _18567_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15779_ _11701_/A _15779_/B _15779_/C VGND VGND VPWR VPWR _15779_/X sky130_fd_sc_hd__and3_4
XANTENNA__14277__A _14277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23171__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21505__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13181__A _12741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24297__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17518_ _13192_/X VGND VGND VPWR VPWR _17518_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22494__A _22508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18498_ _18453_/X _18497_/X _20071_/A _18453_/X VGND VGND VPWR VPWR _18498_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17588__A _16381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17449_ _17396_/D _17447_/X _17448_/Y VGND VGND VPWR VPWR _17449_/X sky130_fd_sc_hd__o21a_4
XFILLER_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20460_ _24269_/Q _20443_/X _20459_/X VGND VGND VPWR VPWR _20460_/X sky130_fd_sc_hd__o21a_4
XFILLER_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19119_ _11516_/A _11515_/Y _11518_/B VGND VGND VPWR VPWR _19119_/X sky130_fd_sc_hd__o21a_4
XFILLER_174_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20391_ _20231_/X _20381_/Y _20389_/X _20390_/Y _20255_/X VGND VGND VPWR VPWR _20391_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19882__B1 _22039_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_17_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_34_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22130_ _22118_/A VGND VGND VPWR VPWR _22130_/X sky130_fd_sc_hd__buf_2
XFILLER_106_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20742__A _20535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22061_ _21838_/X _22060_/X _23497_/Q _22057_/X VGND VGND VPWR VPWR _23497_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15836__A _12871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22233__A2 _22230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14740__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21012_ _24405_/Q _20427_/A _24437_/Q _20282_/A VGND VGND VPWR VPWR _21012_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13356__A _13384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12260__A _11880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21573__A _21549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19937__B2 _20866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22963_ _22947_/X _22963_/B _22963_/C VGND VGND VPWR VPWR _22963_/X sky130_fd_sc_hd__and3_4
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16667__A _16675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21744__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21914_ _21845_/X _21909_/X _13365_/B _21913_/X VGND VGND VPWR VPWR _23590_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15571__A _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22894_ _22897_/A _22894_/B VGND VGND VPWR VPWR HWDATA[28] sky130_fd_sc_hd__nor2_4
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15290__B _23128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21845_ _21560_/A VGND VGND VPWR VPWR _21845_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13091__A _13091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21776_ _21551_/X _21770_/X _23658_/Q _21774_/X VGND VGND VPWR VPWR _21776_/X sky130_fd_sc_hd__o22a_4
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23515_ _23515_/CLK _22030_/X VGND VGND VPWR VPWR _14485_/B sky130_fd_sc_hd__dfxtp_4
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20727_ _20727_/A _20617_/B VGND VGND VPWR VPWR _20727_/Y sky130_fd_sc_hd__nand2_4
X_24495_ _24495_/CLK _24495_/D HRESETn VGND VGND VPWR VPWR _20003_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14915__A _11697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23446_ _23095_/CLK _23446_/D VGND VGND VPWR VPWR _14875_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20658_ _20658_/A VGND VGND VPWR VPWR _21280_/A sky130_fd_sc_hd__buf_2
XFILLER_109_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23377_ _23537_/CLK _22283_/X VGND VGND VPWR VPWR _16756_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12435__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20589_ _18325_/X _20446_/X _20538_/X _20588_/Y VGND VGND VPWR VPWR _20589_/X sky130_fd_sc_hd__a211o_4
XFILLER_152_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13130_ _12696_/A _13199_/B VGND VGND VPWR VPWR _13130_/X sky130_fd_sc_hd__or2_4
XFILLER_109_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22328_ _16048_/B VGND VGND VPWR VPWR _23342_/D sky130_fd_sc_hd__buf_2
XANTENNA__21748__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13061_ _13096_/A _13059_/X _13061_/C VGND VGND VPWR VPWR _13061_/X sky130_fd_sc_hd__and3_4
XFILLER_140_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22259_ _22146_/X _22258_/X _23391_/Q _22255_/X VGND VGND VPWR VPWR _23391_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14650__A _14658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20371__B _20371_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12012_ _12012_/A _23828_/Q VGND VGND VPWR VPWR _12013_/C sky130_fd_sc_hd__or2_4
XANTENNA__15465__B _15465_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21983__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16820_ _16819_/X VGND VGND VPWR VPWR _16821_/B sky130_fd_sc_hd__inv_2
XANTENNA__13266__A _13125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22579__A _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19928__B2 _20339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16751_ _16788_/A _16751_/B VGND VGND VPWR VPWR _16753_/B sky130_fd_sc_hd__or2_4
XFILLER_4_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13963_ _13990_/A _24032_/Q VGND VGND VPWR VPWR _13965_/B sky130_fd_sc_hd__or2_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16577__A _16592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21735__B2 _21731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15702_ _13304_/A _15702_/B VGND VGND VPWR VPWR _15702_/X sky130_fd_sc_hd__or2_4
XANTENNA__15481__A _12626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12914_ _11857_/A _11631_/A _12883_/X _11607_/A _12913_/X VGND VGND VPWR VPWR _12914_/X
+ sky130_fd_sc_hd__a32o_4
X_19470_ _19441_/X _19467_/X _18027_/X _19469_/X VGND VGND VPWR VPWR _24212_/D sky130_fd_sc_hd__o22a_4
X_16682_ _16682_/A _16682_/B _16681_/X VGND VGND VPWR VPWR _16683_/C sky130_fd_sc_hd__or3_4
XFILLER_74_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13894_ _13894_/A _13894_/B _13894_/C VGND VGND VPWR VPWR _13912_/B sky130_fd_sc_hd__and3_4
XANTENNA__20099__A _20124_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18421_ _17396_/B _18420_/X _17446_/X VGND VGND VPWR VPWR _18421_/X sky130_fd_sc_hd__o21a_4
X_12845_ _12845_/A VGND VGND VPWR VPWR _12846_/B sky130_fd_sc_hd__inv_2
X_15633_ _13928_/A _15633_/B _15632_/X VGND VGND VPWR VPWR _15633_/X sky130_fd_sc_hd__and3_4
XFILLER_34_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18352_ _18180_/X _17773_/X _17694_/X VGND VGND VPWR VPWR _18352_/X sky130_fd_sc_hd__o21a_4
X_12776_ _12773_/X _12774_/X _12775_/X VGND VGND VPWR VPWR _12776_/X sky130_fd_sc_hd__and3_4
X_15564_ _14431_/A _15562_/X _15563_/X VGND VGND VPWR VPWR _15564_/X sky130_fd_sc_hd__and3_4
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _14548_/X _17303_/B VGND VGND VPWR VPWR _17621_/B sky130_fd_sc_hd__or2_4
XANTENNA__22160__B2 _22154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11727_/A VGND VGND VPWR VPWR _16454_/A sky130_fd_sc_hd__buf_2
X_14515_ _13229_/A _14498_/X _14514_/X VGND VGND VPWR VPWR _14547_/B sky130_fd_sc_hd__or3_4
XFILLER_148_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15495_ _13743_/A _15493_/X _15495_/C VGND VGND VPWR VPWR _15495_/X sky130_fd_sc_hd__and3_4
XFILLER_30_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18283_ _18283_/A _18283_/B _18281_/Y _18283_/D VGND VGND VPWR VPWR _18284_/A sky130_fd_sc_hd__or4_4
XANTENNA__14825__A _15106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17234_ _17231_/X _17187_/X _17233_/X _17184_/X VGND VGND VPWR VPWR _17234_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11658_ _14772_/A VGND VGND VPWR VPWR _11659_/A sky130_fd_sc_hd__buf_2
X_14446_ _14311_/A _14502_/B VGND VGND VPWR VPWR _14446_/X sky130_fd_sc_hd__or2_4
XFILLER_122_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _14377_/A VGND VGND VPWR VPWR _14378_/A sky130_fd_sc_hd__buf_2
X_17165_ _13266_/X VGND VGND VPWR VPWR _17165_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11589_ _16901_/A VGND VGND VPWR VPWR _16921_/A sky130_fd_sc_hd__buf_2
XFILLER_155_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13328_ _13319_/A _23238_/Q VGND VGND VPWR VPWR _13328_/X sky130_fd_sc_hd__or2_4
X_16116_ _16116_/A _16116_/B _16116_/C VGND VGND VPWR VPWR _16116_/X sky130_fd_sc_hd__and3_4
XFILLER_170_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21658__A _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17096_ _17096_/A _17082_/B VGND VGND VPWR VPWR _17097_/A sky130_fd_sc_hd__or2_4
X_16047_ _16047_/A _16047_/B _16047_/C VGND VGND VPWR VPWR _16051_/B sky130_fd_sc_hd__and3_4
X_13259_ _11682_/A _13259_/B _13259_/C VGND VGND VPWR VPWR _13260_/C sky130_fd_sc_hd__and3_4
XANTENNA__14560__A _14278_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19806_ _19806_/A _19705_/A VGND VGND VPWR VPWR _19806_/X sky130_fd_sc_hd__or2_4
XFILLER_69_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23537__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17998_ _17809_/X _17992_/X _17848_/X _17997_/X VGND VGND VPWR VPWR _17998_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22489__A _22489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19737_ _19898_/B _19684_/X _19714_/X VGND VGND VPWR VPWR _19737_/Y sky130_fd_sc_hd__a21oi_4
X_16949_ _16949_/A VGND VGND VPWR VPWR _17660_/A sky130_fd_sc_hd__inv_2
XANTENNA__16487__A _16362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21726__B2 _21724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13904__A _13916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19668_ _19589_/X _19642_/A _19596_/X VGND VGND VPWR VPWR _19668_/X sky130_fd_sc_hd__o21a_4
XFILLER_37_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_8_0_HCLK clkbuf_5_8_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16602__B1 _11608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23687__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18619_ _16927_/Y _18597_/Y _18614_/Y _17013_/X _18618_/X VGND VGND VPWR VPWR _18619_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19798__A _19823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19599_ _19661_/A VGND VGND VPWR VPWR _19744_/A sky130_fd_sc_hd__buf_2
XFILLER_52_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21630_ _21558_/X _21627_/X _23751_/Q _21624_/X VGND VGND VPWR VPWR _23751_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19698__A3 _21007_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21561_ _21549_/A VGND VGND VPWR VPWR _21561_/X sky130_fd_sc_hd__buf_2
XFILLER_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23300_ _23588_/CLK _23300_/D VGND VGND VPWR VPWR _15668_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20512_ _20380_/A _20512_/B VGND VGND VPWR VPWR _20512_/X sky130_fd_sc_hd__and2_4
X_24280_ _24287_/CLK _19314_/X HRESETn VGND VGND VPWR VPWR _24280_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21492_ _21492_/A VGND VGND VPWR VPWR _21492_/X sky130_fd_sc_hd__buf_2
XFILLER_159_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23231_ _24096_/CLK _23231_/D VGND VGND VPWR VPWR _23231_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_140_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20443_ _20229_/X VGND VGND VPWR VPWR _20443_/X sky130_fd_sc_hd__buf_2
XANTENNA__12255__A _12279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20465__A1 _20418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20465__B2 _20396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_opt_0_HCLK _24472_/CLK VGND VGND VPWR VPWR _23509_/CLK sky130_fd_sc_hd__clkbuf_16
X_23162_ _23641_/CLK _23162_/D VGND VGND VPWR VPWR _14649_/B sky130_fd_sc_hd__dfxtp_4
X_20374_ _20231_/X _20365_/Y _20372_/X _20373_/Y _20255_/X VGND VGND VPWR VPWR _20374_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17330__A1 _17327_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24312__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22113_ _22113_/A VGND VGND VPWR VPWR _22113_/X sky130_fd_sc_hd__buf_2
XANTENNA__22206__A2 _22201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14470__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23093_ _23392_/CLK _22735_/X VGND VGND VPWR VPWR _23093_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22044_ _22038_/Y _22043_/X _21811_/X _22043_/X VGND VGND VPWR VPWR _23508_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21965__B2 _21964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13086__A _13103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18830__A1 _15251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23995_ _23592_/CLK _21175_/X VGND VGND VPWR VPWR _23995_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16397__A _16007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22946_ _19319_/X VGND VGND VPWR VPWR _22946_/X sky130_fd_sc_hd__buf_2
XFILLER_21_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21193__A2 _21191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22877_ _20665_/X VGND VGND VPWR VPWR _22877_/X sky130_fd_sc_hd__buf_2
XFILLER_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12630_ _12630_/A VGND VGND VPWR VPWR _12945_/A sky130_fd_sc_hd__buf_2
XANTENNA__22846__B _22846_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21828_ _21826_/X _21827_/X _16057_/B _21822_/X VGND VGND VPWR VPWR _21828_/X sky130_fd_sc_hd__o22a_4
XFILLER_19_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _12561_/A _12672_/B VGND VGND VPWR VPWR _12562_/C sky130_fd_sc_hd__or2_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21759_ _21774_/A VGND VGND VPWR VPWR _21767_/A sky130_fd_sc_hd__buf_2
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11512_ _24163_/Q VGND VGND VPWR VPWR _11638_/A sky130_fd_sc_hd__inv_2
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17021__A _17020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14300_ _12469_/A _14298_/X _14300_/C VGND VGND VPWR VPWR _14301_/C sky130_fd_sc_hd__and3_4
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15280_ _15022_/A _15276_/X _15279_/X VGND VGND VPWR VPWR _15280_/X sky130_fd_sc_hd__or3_4
X_12492_ _12492_/A VGND VGND VPWR VPWR _12493_/A sky130_fd_sc_hd__buf_2
X_24478_ _24137_/CLK _18573_/X HRESETn VGND VGND VPWR VPWR _24478_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ _14240_/A _24063_/Q VGND VGND VPWR VPWR _14231_/X sky130_fd_sc_hd__or2_4
X_23429_ _23397_/CLK _23429_/D VGND VGND VPWR VPWR _13546_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24344__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21478__A _21492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14162_ _12453_/A _23647_/Q VGND VGND VPWR VPWR _14163_/C sky130_fd_sc_hd__or2_4
XANTENNA__17675__B _17473_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20382__A _20847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13113_ _13089_/A _23880_/Q VGND VGND VPWR VPWR _13114_/C sky130_fd_sc_hd__or2_4
XANTENNA__14135__A1 _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18970_ _18959_/X _18969_/X _18959_/X _24370_/Q VGND VGND VPWR VPWR _18970_/X sky130_fd_sc_hd__a2bb2o_4
X_14093_ _11910_/A VGND VGND VPWR VPWR _14094_/A sky130_fd_sc_hd__buf_2
XANTENNA__20208__A1 _19402_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_63_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13044_ _11915_/A _13044_/B _13044_/C VGND VGND VPWR VPWR _13045_/C sky130_fd_sc_hd__and3_4
X_17921_ _17815_/X _17123_/B _17820_/X _17142_/X VGND VGND VPWR VPWR _17921_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18787__A _18796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21956__B2 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18821__A1 _17153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17852_ _17233_/X _17199_/X _17231_/X _17183_/X VGND VGND VPWR VPWR _17852_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16803_ _16791_/A _23121_/Q VGND VGND VPWR VPWR _16803_/X sky130_fd_sc_hd__or2_4
XFILLER_94_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17783_ _17655_/A _17252_/Y VGND VGND VPWR VPWR _17783_/X sky130_fd_sc_hd__or2_4
X_14995_ _14171_/A _14992_/X _14995_/C VGND VGND VPWR VPWR _14995_/X sky130_fd_sc_hd__and3_4
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13724__A _13697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19522_ _19680_/A VGND VGND VPWR VPWR _19687_/D sky130_fd_sc_hd__buf_2
X_16734_ _12051_/A _23505_/Q VGND VGND VPWR VPWR _16736_/B sky130_fd_sc_hd__or2_4
X_13946_ _13945_/X VGND VGND VPWR VPWR _13946_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16100__A _16099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22381__B2 _22380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21941__A _21941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19453_ _19452_/X VGND VGND VPWR VPWR _19454_/A sky130_fd_sc_hd__buf_2
XANTENNA__24145__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16665_ _16658_/A _16665_/B VGND VGND VPWR VPWR _16666_/C sky130_fd_sc_hd__or2_4
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13877_ _13877_/A VGND VGND VPWR VPWR _14377_/A sky130_fd_sc_hd__buf_2
XANTENNA__20931__A2 _20313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18404_ _18370_/B _18402_/X _18358_/X _22990_/C VGND VGND VPWR VPWR _18404_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19411__A _19406_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15616_ _15616_/A _15612_/X _15616_/C VGND VGND VPWR VPWR _15617_/C sky130_fd_sc_hd__or3_4
X_12828_ _13387_/A _23722_/Q VGND VGND VPWR VPWR _12831_/B sky130_fd_sc_hd__or2_4
X_19384_ _19328_/Y _17000_/Y _19328_/A _16999_/X VGND VGND VPWR VPWR _23078_/B sky130_fd_sc_hd__o22a_4
X_16596_ _16593_/A _23730_/Q VGND VGND VPWR VPWR _16598_/B sky130_fd_sc_hd__or2_4
XANTENNA__22133__B2 _22130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18335_ _18335_/A _18335_/B VGND VGND VPWR VPWR _18337_/C sky130_fd_sc_hd__and2_4
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15547_ _14421_/A _15607_/B VGND VGND VPWR VPWR _15547_/X sky130_fd_sc_hd__or2_4
X_12759_ _12759_/A _12759_/B VGND VGND VPWR VPWR _12759_/X sky130_fd_sc_hd__or2_4
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22684__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14555__A _12427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18266_ _17809_/X _17997_/X _17882_/X VGND VGND VPWR VPWR _18266_/X sky130_fd_sc_hd__o21a_4
X_15478_ _12592_/A _15478_/B VGND VGND VPWR VPWR _15478_/X sky130_fd_sc_hd__or2_4
XANTENNA__17560__A1 _17556_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17217_ _17128_/A _17213_/X _17113_/X _17216_/X VGND VGND VPWR VPWR _17217_/X sky130_fd_sc_hd__o22a_4
X_14429_ _12435_/A _14491_/B VGND VGND VPWR VPWR _14431_/B sky130_fd_sc_hd__or2_4
XFILLER_156_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22436__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18197_ _18197_/A VGND VGND VPWR VPWR _18197_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12075__A _11984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21388__A _21388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17148_ _17130_/X _17143_/X _17124_/X _17147_/X VGND VGND VPWR VPWR _17148_/X sky130_fd_sc_hd__o22a_4
XFILLER_157_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14290__A _12504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17079_ _17078_/X VGND VGND VPWR VPWR _17079_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12803__A _12833_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24485__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13618__B _13721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20090_ _19402_/A _17006_/A _20070_/X _20089_/X VGND VGND VPWR VPWR _20091_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21947__B2 _21943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17076__B1 _16918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18812__A1 _13567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16929__B _17087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15833__B _15833_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22800_ _16922_/C _18774_/X VGND VGND VPWR VPWR _22800_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13634__A _11623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23780_ _23111_/CLK _23780_/D VGND VGND VPWR VPWR _23780_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16010__A _16009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20992_ _20992_/A VGND VGND VPWR VPWR _20992_/Y sky130_fd_sc_hd__inv_2
XFILLER_168_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21175__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22372__B2 _22366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22731_ _20938_/A _22729_/X _14827_/B _22726_/X VGND VGND VPWR VPWR _22731_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21851__A _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20383__B1 _24464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22662_ _22655_/A VGND VGND VPWR VPWR _22662_/X sky130_fd_sc_hd__buf_2
XFILLER_164_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22124__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24401_ _23281_/CLK _24401_/D HRESETn VGND VGND VPWR VPWR _24401_/Q sky130_fd_sc_hd__dfstp_4
X_21613_ _21620_/A VGND VGND VPWR VPWR _21613_/X sky130_fd_sc_hd__buf_2
XANTENNA__18879__A1 _14548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22593_ _22622_/A VGND VGND VPWR VPWR _22608_/A sky130_fd_sc_hd__buf_2
XANTENNA__14465__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20686__A1 _18448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24332_ _24277_/CLK _19178_/X HRESETn VGND VGND VPWR VPWR _19153_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_166_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21544_ _20464_/A VGND VGND VPWR VPWR _21544_/X sky130_fd_sc_hd__buf_2
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14184__B _23519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24263_ _24271_/CLK _19353_/X HRESETn VGND VGND VPWR VPWR _24263_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11601__B _17398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22427__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21475_ _21482_/A VGND VGND VPWR VPWR _21475_/X sky130_fd_sc_hd__buf_2
XFILLER_135_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23214_ _23662_/CLK _23214_/D VGND VGND VPWR VPWR _23214_/Q sky130_fd_sc_hd__dfxtp_4
X_20426_ _18835_/X VGND VGND VPWR VPWR _20427_/A sky130_fd_sc_hd__buf_2
X_24194_ _23383_/CLK _19821_/Y HRESETn VGND VGND VPWR VPWR _11643_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_174_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23145_ _23561_/CLK _22659_/X VGND VGND VPWR VPWR _23145_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15296__A _13788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13809__A _12445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20357_ _20231_/X _20340_/Y _20355_/X _20356_/Y _20255_/X VGND VGND VPWR VPWR _20357_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12713__A _12702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23076_ _19953_/A _16945_/X _23048_/X _23075_/X VGND VGND VPWR VPWR _23076_/X sky130_fd_sc_hd__a211o_4
X_20288_ _20267_/X VGND VGND VPWR VPWR _20315_/A sky130_fd_sc_hd__inv_2
XFILLER_121_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22027_ _21867_/X _22024_/X _13800_/B _22021_/X VGND VGND VPWR VPWR _23517_/D sky130_fd_sc_hd__o22a_4
XFILLER_76_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18400__A _18399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13544__A _13543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13800_ _15393_/A _13800_/B VGND VGND VPWR VPWR _13801_/C sky130_fd_sc_hd__or2_4
XANTENNA__24208__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14780_ _14675_/A _14780_/B VGND VGND VPWR VPWR _14781_/C sky130_fd_sc_hd__or2_4
X_11992_ _11939_/X _11987_/X _11992_/C VGND VGND VPWR VPWR _11992_/X sky130_fd_sc_hd__or3_4
X_23978_ _24074_/CLK _21204_/X VGND VGND VPWR VPWR _23978_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22363__B2 _22359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13731_ _12576_/A _13715_/X _13730_/X VGND VGND VPWR VPWR _13749_/B sky130_fd_sc_hd__and3_4
X_22929_ _22929_/A _24136_/Q VGND VGND VPWR VPWR _22933_/B sky130_fd_sc_hd__or2_4
XFILLER_21_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16450_ _16130_/A _16427_/X _16434_/X _16441_/X _16449_/X VGND VGND VPWR VPWR _16450_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_32_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13662_ _13662_/A VGND VGND VPWR VPWR _13663_/A sky130_fd_sc_hd__buf_2
XANTENNA__20377__A _20377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15401_ _15401_/A _15399_/X _15401_/C VGND VGND VPWR VPWR _15401_/X sky130_fd_sc_hd__and3_4
X_12613_ _12954_/A _12603_/X _12613_/C VGND VGND VPWR VPWR _12614_/C sky130_fd_sc_hd__or3_4
XANTENNA__11999__A _12108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13593_ _13593_/A VGND VGND VPWR VPWR _14448_/A sky130_fd_sc_hd__buf_2
X_16381_ _16380_/X VGND VGND VPWR VPWR _16381_/X sky130_fd_sc_hd__buf_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18120_ _18120_/A VGND VGND VPWR VPWR _18120_/Y sky130_fd_sc_hd__inv_2
X_12544_ _12890_/A _12536_/X _12544_/C VGND VGND VPWR VPWR _12544_/X sky130_fd_sc_hd__or3_4
XFILLER_129_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15332_ _15318_/A _23928_/Q VGND VGND VPWR VPWR _15334_/B sky130_fd_sc_hd__or2_4
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18051_ _18051_/A VGND VGND VPWR VPWR _18653_/B sky130_fd_sc_hd__inv_2
X_15263_ _14154_/A _24024_/Q VGND VGND VPWR VPWR _15263_/X sky130_fd_sc_hd__or2_4
X_12475_ _13642_/A VGND VGND VPWR VPWR _14325_/A sky130_fd_sc_hd__buf_2
X_17002_ _24212_/Q VGND VGND VPWR VPWR _17009_/A sky130_fd_sc_hd__inv_2
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14214_ _14199_/A _23679_/Q VGND VGND VPWR VPWR _14217_/B sky130_fd_sc_hd__or2_4
X_15194_ _14196_/A _15130_/B VGND VGND VPWR VPWR _15195_/C sky130_fd_sc_hd__or2_4
XANTENNA__14822__B _23385_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14145_ _11898_/A _23839_/Q VGND VGND VPWR VPWR _14146_/C sky130_fd_sc_hd__or2_4
XANTENNA__13719__A _13719_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12623__A _12623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18953_ _18952_/Y _18953_/B VGND VGND VPWR VPWR _18953_/X sky130_fd_sc_hd__and2_4
X_14076_ _12581_/A _24096_/Q VGND VGND VPWR VPWR _14077_/C sky130_fd_sc_hd__or2_4
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20840__A _20840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21929__B2 _21927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13027_ _12472_/A _13027_/B _13027_/C VGND VGND VPWR VPWR _13031_/B sky130_fd_sc_hd__and3_4
X_17904_ _17659_/A VGND VGND VPWR VPWR _17904_/X sky130_fd_sc_hd__buf_2
XANTENNA__15934__A _12516_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19406__A _19324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18884_ _15118_/X _18840_/A _24406_/Q _18843_/A VGND VGND VPWR VPWR _24406_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18310__A _18310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17835_ _17233_/A _17157_/X _17817_/A _17163_/X VGND VGND VPWR VPWR _17835_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24326__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17766_ _16982_/A _17368_/X _17715_/X _17765_/X VGND VGND VPWR VPWR _17767_/C sky130_fd_sc_hd__o22a_4
X_14978_ _14771_/A _14976_/X _14978_/C VGND VGND VPWR VPWR _14979_/C sky130_fd_sc_hd__and3_4
XANTENNA__21157__A2 _21155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19505_ _19560_/A _19528_/B VGND VGND VPWR VPWR _19680_/A sky130_fd_sc_hd__or2_4
X_16717_ _16568_/A _16717_/B _16716_/X VGND VGND VPWR VPWR _16718_/B sky130_fd_sc_hd__or3_4
XANTENNA__20365__B1 _20235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13929_ _13916_/A _13929_/B VGND VGND VPWR VPWR _13929_/X sky130_fd_sc_hd__or2_4
X_17697_ _17697_/A _17697_/B _17696_/X VGND VGND VPWR VPWR _17698_/C sky130_fd_sc_hd__or3_4
X_19436_ _22910_/B VGND VGND VPWR VPWR _19438_/A sky130_fd_sc_hd__buf_2
XANTENNA__19770__A2 HRDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16648_ _16672_/A _23346_/Q VGND VGND VPWR VPWR _16648_/X sky130_fd_sc_hd__or2_4
XFILLER_35_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20117__B1 _19399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19367_ _19365_/X _18571_/X _19365_/X _20814_/A VGND VGND VPWR VPWR _19367_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22657__A2 _22651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14285__A _14307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16579_ _16539_/X _23858_/Q VGND VGND VPWR VPWR _16580_/C sky130_fd_sc_hd__or2_4
XFILLER_163_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11702__A _13367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18318_ _18318_/A VGND VGND VPWR VPWR _18464_/B sky130_fd_sc_hd__inv_2
XFILLER_124_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19298_ _19237_/A _19237_/B _19297_/Y VGND VGND VPWR VPWR _24288_/D sky130_fd_sc_hd__o21a_4
XANTENNA__12517__B _12618_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18249_ _16958_/A _18248_/X VGND VGND VPWR VPWR _18249_/X sky130_fd_sc_hd__and2_4
XFILLER_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21260_ _21259_/X _21257_/X _23949_/Q _21252_/X VGND VGND VPWR VPWR _21260_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22007__A _22007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20211_ _22687_/A _19852_/A _19863_/A VGND VGND VPWR VPWR _22487_/A sky130_fd_sc_hd__or3_4
XANTENNA__13629__A _13658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21093__B2 _21087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21191_ _21198_/A VGND VGND VPWR VPWR _21191_/X sky130_fd_sc_hd__buf_2
XANTENNA__24390__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12533__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20142_ _20142_/A VGND VGND VPWR VPWR _20142_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15844__A _12906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20073_ _20064_/X _18478_/A _20070_/X _20072_/X VGND VGND VPWR VPWR _20074_/A sky130_fd_sc_hd__o22a_4
XFILLER_112_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21396__A2 _21391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23901_ _23518_/CLK _23901_/D VGND VGND VPWR VPWR _13831_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23832_ _23098_/CLK _23832_/D VGND VGND VPWR VPWR _23832_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23763_ _23760_/CLK _23763_/D VGND VGND VPWR VPWR _23763_/Q sky130_fd_sc_hd__dfxtp_4
X_20975_ _24247_/Q VGND VGND VPWR VPWR _20975_/Y sky130_fd_sc_hd__inv_2
XPHY_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16675__A _16675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24500__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22714_ _21848_/A _22708_/X _13476_/B _22712_/X VGND VGND VPWR VPWR _23109_/D sky130_fd_sc_hd__o22a_4
XFILLER_0_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23694_ _23501_/CLK _21721_/X VGND VGND VPWR VPWR _23694_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22645_ _22412_/X _22644_/X _12155_/B _22641_/X VGND VGND VPWR VPWR _23155_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14195__A _14225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22576_ _22555_/A VGND VGND VPWR VPWR _22576_/X sky130_fd_sc_hd__buf_2
XFILLER_167_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21527_ _21520_/Y _21525_/X _21526_/X _21525_/X VGND VGND VPWR VPWR _23796_/D sky130_fd_sc_hd__a2bb2o_4
X_24315_ _24287_/CLK _19212_/X HRESETn VGND VGND VPWR VPWR _19136_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_127_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12260_ _11880_/A _12260_/B _12259_/X VGND VGND VPWR VPWR _12260_/X sky130_fd_sc_hd__and3_4
X_24246_ _24248_/CLK _19380_/X HRESETn VGND VGND VPWR VPWR _24246_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21458_ _21297_/X _21455_/X _13839_/B _21452_/X VGND VGND VPWR VPWR _23837_/D sky130_fd_sc_hd__o22a_4
X_20409_ _18062_/X _20847_/A _20638_/A _20408_/Y VGND VGND VPWR VPWR _20409_/X sky130_fd_sc_hd__a211o_4
X_12191_ _12191_/A VGND VGND VPWR VPWR _13042_/A sky130_fd_sc_hd__buf_2
XFILLER_107_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24177_ _24184_/CLK _24177_/D HRESETn VGND VGND VPWR VPWR _24177_/Q sky130_fd_sc_hd__dfrtp_4
X_21389_ _21263_/X _21384_/X _12665_/B _21388_/X VGND VGND VPWR VPWR _23883_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12443__A _15018_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11572__A1 _20157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23128_ _23192_/CLK _23128_/D VGND VGND VPWR VPWR _23128_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15754__A _13090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15950_ _15944_/A _23214_/Q VGND VGND VPWR VPWR _15952_/B sky130_fd_sc_hd__or2_4
XFILLER_110_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23059_ _22922_/A _17902_/Y _17965_/X VGND VGND VPWR VPWR _23061_/B sky130_fd_sc_hd__or3_4
XANTENNA__19226__A _24129_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24490__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21387__A2 _21384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14901_ _14133_/A _14896_/X _14901_/C VGND VGND VPWR VPWR _14901_/X sky130_fd_sc_hd__or3_4
XANTENNA__22584__B2 _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15473__B _15473_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15881_ _13531_/A _15819_/B VGND VGND VPWR VPWR _15883_/B sky130_fd_sc_hd__or2_4
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13274__A _12561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17620_ _17618_/Y _17620_/B VGND VGND VPWR VPWR _17620_/X sky130_fd_sc_hd__or2_4
X_14832_ _14680_/A _14832_/B _14831_/X VGND VGND VPWR VPWR _14832_/X sky130_fd_sc_hd__and3_4
XFILLER_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14089__B _23263_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24180__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17551_ _17120_/Y _17551_/B VGND VGND VPWR VPWR _17642_/A sky130_fd_sc_hd__or2_4
X_14763_ _13663_/A _14759_/X _14762_/X VGND VGND VPWR VPWR _14763_/X sky130_fd_sc_hd__or3_4
X_11975_ _11975_/A _23956_/Q VGND VGND VPWR VPWR _11977_/B sky130_fd_sc_hd__or2_4
XANTENNA__16015__A1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16015__B2 _16014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16502_ _16474_/A _16500_/X _16502_/C VGND VGND VPWR VPWR _16502_/X sky130_fd_sc_hd__and3_4
XANTENNA__17212__B1 _17153_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23748__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13714_ _13774_/A _13711_/X _13713_/X VGND VGND VPWR VPWR _13714_/X sky130_fd_sc_hd__and3_4
X_17482_ _17047_/A _17481_/X _17050_/X VGND VGND VPWR VPWR _17482_/X sky130_fd_sc_hd__o21a_4
X_14694_ _14657_/A _14600_/B VGND VGND VPWR VPWR _14696_/B sky130_fd_sc_hd__or2_4
X_19221_ _19131_/X VGND VGND VPWR VPWR _19221_/Y sky130_fd_sc_hd__inv_2
X_16433_ _16094_/A _16431_/X _16432_/X VGND VGND VPWR VPWR _16433_/X sky130_fd_sc_hd__and3_4
XANTENNA__13721__B _13721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13645_ _11913_/A _13643_/X _13644_/X VGND VGND VPWR VPWR _13649_/B sky130_fd_sc_hd__and3_4
XFILLER_72_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19152_ _24331_/Q _19151_/X VGND VGND VPWR VPWR _19153_/B sky130_fd_sc_hd__and2_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16364_ _16318_/A _16301_/B VGND VGND VPWR VPWR _16364_/X sky130_fd_sc_hd__or2_4
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _12987_/X _16832_/A VGND VGND VPWR VPWR _15932_/A sky130_fd_sc_hd__or2_4
XANTENNA__20835__A _20834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ _18013_/C _18013_/B _17667_/X VGND VGND VPWR VPWR _18103_/X sky130_fd_sc_hd__o21a_4
XFILLER_40_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15315_ _11720_/A VGND VGND VPWR VPWR _15319_/A sky130_fd_sc_hd__buf_2
X_19083_ _11524_/A _11524_/B _19076_/Y VGND VGND VPWR VPWR _19083_/Y sky130_fd_sc_hd__a21oi_4
X_12527_ _13974_/A VGND VGND VPWR VPWR _15000_/A sky130_fd_sc_hd__buf_2
XFILLER_157_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16295_ _15952_/A _16293_/X _16294_/X VGND VGND VPWR VPWR _16295_/X sky130_fd_sc_hd__and3_4
XFILLER_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18034_ _18517_/A VGND VGND VPWR VPWR _18310_/A sky130_fd_sc_hd__buf_2
X_15246_ _14635_/A _15246_/B _15246_/C VGND VGND VPWR VPWR _15247_/C sky130_fd_sc_hd__and3_4
XFILLER_68_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12458_ _12536_/A _12458_/B _12458_/C VGND VGND VPWR VPWR _12459_/C sky130_fd_sc_hd__and3_4
XFILLER_172_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13449__A _12867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24400__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21075__B2 _21070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12389_ _12827_/A _12389_/B VGND VGND VPWR VPWR _12389_/X sky130_fd_sc_hd__or2_4
XANTENNA__12353__A _13123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15177_ _15017_/A _15177_/B VGND VGND VPWR VPWR _15178_/C sky130_fd_sc_hd__or2_4
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14128_ _14110_/A _23583_/Q VGND VGND VPWR VPWR _14129_/C sky130_fd_sc_hd__or2_4
XFILLER_141_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19985_ _17786_/X _19983_/X _19984_/Y _19979_/X VGND VGND VPWR VPWR _19985_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18936_ _14548_/X _18934_/X _19101_/A _18935_/X VGND VGND VPWR VPWR _24379_/D sky130_fd_sc_hd__o22a_4
X_14059_ _13700_/A _23136_/Q VGND VGND VPWR VPWR _14059_/X sky130_fd_sc_hd__or2_4
XFILLER_140_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21378__A2 _21377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22575__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18867_ _15916_/X _18863_/X _20677_/A _18864_/X VGND VGND VPWR VPWR _24419_/D sky130_fd_sc_hd__o22a_4
XFILLER_94_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13184__A _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17818_ _17816_/X _17134_/X _17817_/X _17117_/X VGND VGND VPWR VPWR _17818_/X sky130_fd_sc_hd__o22a_4
X_18798_ _16381_/X _18796_/X _24463_/Q _18797_/X VGND VGND VPWR VPWR _24463_/D sky130_fd_sc_hd__o22a_4
XFILLER_130_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17749_ _17749_/A _17329_/X VGND VGND VPWR VPWR _17749_/X sky130_fd_sc_hd__and2_4
XFILLER_78_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13912__A _11675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20760_ _20755_/X _20759_/X _24352_/Q _20708_/X VGND VGND VPWR VPWR _20760_/X sky130_fd_sc_hd__o22a_4
XFILLER_35_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21550__A2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19419_ _19418_/X _18482_/Y _19418_/X _24225_/Q VGND VGND VPWR VPWR _24225_/D sky130_fd_sc_hd__a2bb2o_4
X_20691_ _24227_/Q _20636_/X _20690_/X VGND VGND VPWR VPWR _20692_/A sky130_fd_sc_hd__o21a_4
XANTENNA__12528__A _15000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22430_ _20485_/A VGND VGND VPWR VPWR _22430_/X sky130_fd_sc_hd__buf_2
XANTENNA__16309__A2 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15839__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22361_ _22357_/A VGND VGND VPWR VPWR _22376_/A sky130_fd_sc_hd__buf_2
XFILLER_164_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14743__A _13652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24100_ _23908_/CLK _20660_/X VGND VGND VPWR VPWR _15702_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18215__A _18019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21312_ _21311_/X _21305_/X _15146_/B _21239_/X VGND VGND VPWR VPWR _23927_/D sky130_fd_sc_hd__o22a_4
X_22292_ _22117_/X _22287_/X _23371_/Q _22291_/X VGND VGND VPWR VPWR _22292_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22960__A _19438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14462__B _14462_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24031_ _23880_/CLK _24031_/D VGND VGND VPWR VPWR _24031_/Q sky130_fd_sc_hd__dfxtp_4
X_21243_ _21528_/A VGND VGND VPWR VPWR _21243_/X sky130_fd_sc_hd__buf_2
XANTENNA__22263__B1 _14391_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24053__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20813__A1 _18568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21174_ _20860_/X _21169_/X _23996_/Q _21173_/X VGND VGND VPWR VPWR _23996_/D sky130_fd_sc_hd__o22a_4
XFILLER_132_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24248__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20125_ _20125_/A _20125_/B VGND VGND VPWR VPWR _20125_/X sky130_fd_sc_hd__or2_4
XANTENNA__15574__A _14421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22566__B2 _22562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20056_ _24484_/Q VGND VGND VPWR VPWR _20056_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19431__A1 _19399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16245__A1 _16162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13094__A _13094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22318__B2 _22312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23815_ _23111_/CLK _23815_/D VGND VGND VPWR VPWR _23815_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13822__A _14325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11760_ _11759_/X VGND VGND VPWR VPWR _11760_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_53_0_HCLK clkbuf_7_53_0_HCLK/A VGND VGND VPWR VPWR _23203_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23746_ _23656_/CLK _21637_/X VGND VGND VPWR VPWR _23746_/Q sky130_fd_sc_hd__dfxtp_4
X_20958_ _20958_/A VGND VGND VPWR VPWR _20959_/A sky130_fd_sc_hd__buf_2
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _13399_/A VGND VGND VPWR VPWR _13407_/A sky130_fd_sc_hd__buf_2
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12438__A _12854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23677_ _23678_/CLK _23677_/D VGND VGND VPWR VPWR _23677_/Q sky130_fd_sc_hd__dfxtp_4
X_20889_ _20935_/A _20888_/X VGND VGND VPWR VPWR _20889_/X sky130_fd_sc_hd__or2_4
XPHY_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _13462_/A _24037_/Q VGND VGND VPWR VPWR _13433_/B sky130_fd_sc_hd__or2_4
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22628_ _22471_/X _22622_/X _14502_/B _22626_/X VGND VGND VPWR VPWR _22628_/X sky130_fd_sc_hd__o22a_4
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _13376_/A _13361_/B _13361_/C VGND VGND VPWR VPWR _13362_/C sky130_fd_sc_hd__and3_4
XANTENNA__23031__A _22910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22559_ _22437_/X _22558_/X _12922_/B _22555_/X VGND VGND VPWR VPWR _23209_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15749__A _11689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15100_ _15095_/A _23093_/Q VGND VGND VPWR VPWR _15102_/B sky130_fd_sc_hd__or2_4
XFILLER_154_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12312_ _12745_/A _12312_/B _12312_/C VGND VGND VPWR VPWR _12312_/X sky130_fd_sc_hd__and3_4
XFILLER_10_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13292_ _13319_/A _23686_/Q VGND VGND VPWR VPWR _13292_/X sky130_fd_sc_hd__or2_4
X_16080_ _16080_/A _23662_/Q VGND VGND VPWR VPWR _16081_/C sky130_fd_sc_hd__or2_4
XANTENNA__23046__A2 _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21057__B2 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12243_ _12258_/A VGND VGND VPWR VPWR _12311_/A sky130_fd_sc_hd__buf_2
X_15031_ _13607_/A _24085_/Q VGND VGND VPWR VPWR _15031_/X sky130_fd_sc_hd__or2_4
X_24229_ _24134_/CLK _19413_/X HRESETn VGND VGND VPWR VPWR _24229_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12174_ _12167_/A _23667_/Q VGND VGND VPWR VPWR _12175_/C sky130_fd_sc_hd__or2_4
XFILLER_174_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15484__A _12354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19770_ _19519_/X HRDATA[3] _20561_/B _19518_/X VGND VGND VPWR VPWR _19770_/Y sky130_fd_sc_hd__a22oi_4
X_16982_ _16982_/A _16981_/X VGND VGND VPWR VPWR _18433_/A sky130_fd_sc_hd__or2_4
XFILLER_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22557__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18721_ _18721_/A VGND VGND VPWR VPWR _18721_/Y sky130_fd_sc_hd__inv_2
X_15933_ _15933_/A VGND VGND VPWR VPWR _15933_/X sky130_fd_sc_hd__buf_2
XFILLER_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18652_ _18519_/X _18651_/Y _17292_/X VGND VGND VPWR VPWR _18652_/X sky130_fd_sc_hd__o21a_4
X_15864_ _13564_/A _15856_/X _15863_/X VGND VGND VPWR VPWR _15864_/X sky130_fd_sc_hd__and3_4
XANTENNA__23570__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22309__B2 _22305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21780__A2 _21777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17603_ _17513_/X _17603_/B VGND VGND VPWR VPWR _17603_/X sky130_fd_sc_hd__and2_4
X_14815_ _14834_/A _14739_/B VGND VGND VPWR VPWR _14817_/B sky130_fd_sc_hd__or2_4
X_18583_ _17436_/A _18581_/X VGND VGND VPWR VPWR _18583_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22110__A _22110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15795_ _12857_/A _15791_/X _15795_/C VGND VGND VPWR VPWR _15795_/X sky130_fd_sc_hd__or3_4
XFILLER_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17534_ _17527_/D _17532_/X _17533_/Y VGND VGND VPWR VPWR _17534_/X sky130_fd_sc_hd__o21a_4
XFILLER_83_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14746_ _13628_/A _23385_/Q VGND VGND VPWR VPWR _14748_/B sky130_fd_sc_hd__or2_4
X_11958_ _16148_/A VGND VGND VPWR VPWR _11963_/A sky130_fd_sc_hd__buf_2
XFILLER_33_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17465_ _12753_/Y _17021_/X _17021_/X _17464_/X VGND VGND VPWR VPWR _17467_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20740__B1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14677_ _14677_/A VGND VGND VPWR VPWR _14691_/A sky130_fd_sc_hd__buf_2
X_11889_ _13455_/A VGND VGND VPWR VPWR _11889_/X sky130_fd_sc_hd__buf_2
XANTENNA__12348__A _13235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19204_ _24319_/Q _19205_/A _19203_/Y VGND VGND VPWR VPWR _24319_/D sky130_fd_sc_hd__o21a_4
XFILLER_33_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16416_ _16413_/A _16476_/B VGND VGND VPWR VPWR _16416_/X sky130_fd_sc_hd__or2_4
X_13628_ _13628_/A VGND VGND VPWR VPWR _13658_/A sky130_fd_sc_hd__buf_2
XFILLER_34_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17396_ _17396_/A _17396_/B _17387_/Y _17396_/D VGND VGND VPWR VPWR _17437_/A sky130_fd_sc_hd__or4_4
XFILLER_9_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19135_ _19135_/A _19215_/A VGND VGND VPWR VPWR _19213_/A sky130_fd_sc_hd__and2_4
X_16347_ _16192_/A _16279_/B VGND VGND VPWR VPWR _16347_/X sky130_fd_sc_hd__or2_4
XANTENNA__15659__A _11881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21296__B2 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13559_ _13547_/A _13559_/B _13558_/X VGND VGND VPWR VPWR _13563_/B sky130_fd_sc_hd__and3_4
XFILLER_34_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18035__A _18310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14563__A _14304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19066_ _19066_/A VGND VGND VPWR VPWR _19066_/Y sky130_fd_sc_hd__inv_2
X_16278_ _16160_/A _16255_/X _16262_/X _16269_/X _16277_/X VGND VGND VPWR VPWR _16278_/X
+ sky130_fd_sc_hd__a32o_4
X_18017_ _16935_/X _18012_/X _17653_/X _18016_/X VGND VGND VPWR VPWR _18017_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21048__B2 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15229_ _15196_/X _15165_/B VGND VGND VPWR VPWR _15229_/X sky130_fd_sc_hd__or2_4
XFILLER_160_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15394__A _15394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12811__A _12773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19968_ _17807_/A _18755_/X VGND VGND VPWR VPWR _19968_/Y sky130_fd_sc_hd__nor2_4
XFILLER_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18919_ _17172_/X _18913_/X _24390_/Q _18914_/X VGND VGND VPWR VPWR _24390_/D sky130_fd_sc_hd__o22a_4
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19899_ _19899_/A _19899_/B VGND VGND VPWR VPWR _19899_/X sky130_fd_sc_hd__or2_4
XANTENNA__21220__B2 _21216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21930_ _21923_/A VGND VGND VPWR VPWR _21930_/X sky130_fd_sc_hd__buf_2
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21771__A2 _21770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16937__B _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21861_ _21860_/X _21851_/X _23616_/Q _21858_/X VGND VGND VPWR VPWR _23616_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14738__A _15415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23600_ _23500_/CLK _21900_/X VGND VGND VPWR VPWR _16413_/B sky130_fd_sc_hd__dfxtp_4
X_20812_ _20652_/A _20812_/B VGND VGND VPWR VPWR _20812_/Y sky130_fd_sc_hd__nor2_4
XFILLER_36_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17114__A _12097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21792_ _21577_/X _21791_/X _23647_/Q _21788_/X VGND VGND VPWR VPWR _21792_/X sky130_fd_sc_hd__o22a_4
XFILLER_169_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22955__A _18568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22720__B2 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23531_ _23531_/CLK _23531_/D VGND VGND VPWR VPWR _12584_/B sky130_fd_sc_hd__dfxtp_4
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20743_ _24225_/Q _20636_/X _20742_/X VGND VGND VPWR VPWR _20744_/A sky130_fd_sc_hd__o21a_4
XFILLER_51_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12258__A _12258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23462_ _24102_/CLK _23462_/D VGND VGND VPWR VPWR _23462_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20674_ _20641_/X _20673_/X VGND VGND VPWR VPWR _20674_/X sky130_fd_sc_hd__or2_4
XFILLER_17_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22413_ _22462_/A VGND VGND VPWR VPWR _22438_/A sky130_fd_sc_hd__buf_2
XANTENNA__15569__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23393_ _23617_/CLK _23393_/D VGND VGND VPWR VPWR _15562_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14473__A _15395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22344_ _23326_/Q VGND VGND VPWR VPWR _22344_/X sky130_fd_sc_hd__buf_2
XFILLER_163_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22690__A _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21039__B2 _21035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22275_ _22275_/A VGND VGND VPWR VPWR _22291_/A sky130_fd_sc_hd__inv_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24014_ _23438_/CLK _24014_/D VGND VGND VPWR VPWR _24014_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21226_ _21219_/A VGND VGND VPWR VPWR _21226_/X sky130_fd_sc_hd__buf_2
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21157_ _20575_/X _21155_/X _24008_/Q _21152_/X VGND VGND VPWR VPWR _24008_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12721__A _12721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20108_ _11572_/X VGND VGND VPWR VPWR _20108_/Y sky130_fd_sc_hd__inv_2
X_21088_ _21080_/Y _21087_/X _20299_/X _21087_/X VGND VGND VPWR VPWR _21088_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20014__A2 _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21211__B2 _21209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12930_ _12954_/A _12924_/X _12930_/C VGND VGND VPWR VPWR _12930_/X sky130_fd_sc_hd__or3_4
XANTENNA__19504__A _19624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20039_ _20038_/X VGND VGND VPWR VPWR _24150_/D sky130_fd_sc_hd__inv_2
XFILLER_150_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23026__A _18238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ _12886_/A _12861_/B _12861_/C VGND VGND VPWR VPWR _12861_/X sky130_fd_sc_hd__and3_4
XANTENNA__14648__A _13866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14600_ _13658_/A _14600_/B VGND VGND VPWR VPWR _14600_/X sky130_fd_sc_hd__or2_4
XFILLER_15_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11812_ _11812_/A VGND VGND VPWR VPWR _11813_/A sky130_fd_sc_hd__buf_2
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15580_ _13689_/A _15579_/X VGND VGND VPWR VPWR _15580_/X sky130_fd_sc_hd__and2_4
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _13230_/A VGND VGND VPWR VPWR _15770_/A sky130_fd_sc_hd__buf_2
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21514__A2 _21513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22711__B2 _22705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14519_/A _14531_/B VGND VGND VPWR VPWR _14531_/X sky130_fd_sc_hd__or2_4
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _23760_/CLK _21666_/X VGND VGND VPWR VPWR _23729_/Q sky130_fd_sc_hd__dfxtp_4
X_11743_ _11742_/X VGND VGND VPWR VPWR _12168_/A sky130_fd_sc_hd__buf_2
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18391__A1 _17594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18391__B2 _17452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17249_/X VGND VGND VPWR VPWR _17250_/X sky130_fd_sc_hd__buf_2
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _12537_/A _14462_/B VGND VGND VPWR VPWR _14464_/B sky130_fd_sc_hd__or2_4
XFILLER_30_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17678__B _17464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11674_ _11674_/A VGND VGND VPWR VPWR _11675_/A sky130_fd_sc_hd__buf_2
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ _16163_/X _16199_/X _16201_/C VGND VGND VPWR VPWR _16205_/B sky130_fd_sc_hd__and3_4
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _13413_/A _13411_/X _13412_/X VGND VGND VPWR VPWR _13414_/C sky130_fd_sc_hd__and3_4
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15479__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22475__B1 _14618_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17181_ _12077_/X _17150_/X _17151_/X _17180_/X VGND VGND VPWR VPWR _17181_/Y sky130_fd_sc_hd__a22oi_4
X_14393_ _14512_/A _14393_/B _14392_/X VGND VGND VPWR VPWR _14393_/X sky130_fd_sc_hd__and3_4
XFILLER_155_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16132_ _16108_/A _16132_/B VGND VGND VPWR VPWR _16132_/X sky130_fd_sc_hd__or2_4
XFILLER_6_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13344_ _12833_/A VGND VGND VPWR VPWR _13384_/A sky130_fd_sc_hd__buf_2
XFILLER_154_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16063_ _16047_/A _16061_/X _16063_/C VGND VGND VPWR VPWR _16063_/X sky130_fd_sc_hd__and3_4
X_13275_ _13318_/A _13273_/X _13274_/X VGND VGND VPWR VPWR _13275_/X sky130_fd_sc_hd__and3_4
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15014_ _13981_/A _15014_/B VGND VGND VPWR VPWR _15014_/X sky130_fd_sc_hd__and2_4
XFILLER_68_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12226_ _13045_/A VGND VGND VPWR VPWR _12708_/A sky130_fd_sc_hd__buf_2
XFILLER_64_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22105__A _22420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19822_ _19806_/A _19687_/A VGND VGND VPWR VPWR _19822_/X sky130_fd_sc_hd__or2_4
X_12157_ _11705_/X _12155_/X _12156_/X VGND VGND VPWR VPWR _12157_/X sky130_fd_sc_hd__and3_4
XANTENNA__21450__B2 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19753_ _19879_/C _19748_/X _19752_/X VGND VGND VPWR VPWR _19753_/X sky130_fd_sc_hd__a21bo_4
X_16965_ _24141_/Q VGND VGND VPWR VPWR _17721_/A sky130_fd_sc_hd__inv_2
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12088_ _16725_/A _12086_/X _12087_/X VGND VGND VPWR VPWR _12092_/B sky130_fd_sc_hd__and3_4
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15942__A _13327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18704_ _18701_/Y _18703_/X _18701_/Y _18703_/X VGND VGND VPWR VPWR _18704_/X sky130_fd_sc_hd__a2bb2o_4
X_15916_ _15912_/X VGND VGND VPWR VPWR _15916_/X sky130_fd_sc_hd__buf_2
X_19684_ _19683_/X VGND VGND VPWR VPWR _19684_/X sky130_fd_sc_hd__buf_2
XANTENNA__19414__A _19406_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13691__A1 _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16896_ _16896_/A _16852_/X _16887_/X _16896_/D VGND VGND VPWR VPWR _16897_/D sky130_fd_sc_hd__and4_4
XANTENNA__21753__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18635_ _17351_/B _18634_/X VGND VGND VPWR VPWR _18635_/X sky130_fd_sc_hd__or2_4
X_15847_ _12912_/A _15846_/X VGND VGND VPWR VPWR _15847_/X sky130_fd_sc_hd__and2_4
XFILLER_65_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14558__A _14280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13462__A _13462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23316__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18566_ _17412_/B _18564_/X _17890_/X _18565_/X VGND VGND VPWR VPWR _18567_/A sky130_fd_sc_hd__a211o_4
X_15778_ _15778_/A _15705_/B VGND VGND VPWR VPWR _15779_/C sky130_fd_sc_hd__or2_4
XFILLER_80_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21505__A2 _21499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22702__B2 _22698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17517_ _17517_/A VGND VGND VPWR VPWR _17517_/Y sky130_fd_sc_hd__inv_2
X_14729_ _11912_/A _14727_/X _14729_/C VGND VGND VPWR VPWR _14729_/X sky130_fd_sc_hd__and3_4
X_18497_ _18356_/X _18495_/X _18396_/X _18496_/X VGND VGND VPWR VPWR _18497_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12078__A _16568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17448_ _15916_/X _17448_/B VGND VGND VPWR VPWR _17448_/Y sky130_fd_sc_hd__nand2_4
XFILLER_123_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17379_ _17358_/Y VGND VGND VPWR VPWR _17379_/X sky130_fd_sc_hd__buf_2
XANTENNA__12806__A _13556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14293__A _11930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19118_ _19109_/X _19117_/X _19109_/X _11518_/A VGND VGND VPWR VPWR _24344_/D sky130_fd_sc_hd__a2bb2o_4
X_20390_ _24272_/Q VGND VGND VPWR VPWR _20390_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17893__B1 _17014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19049_ _18960_/X VGND VGND VPWR VPWR _19049_/X sky130_fd_sc_hd__buf_2
XFILLER_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22060_ _22060_/A VGND VGND VPWR VPWR _22060_/X sky130_fd_sc_hd__buf_2
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15836__B _15836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14740__B _24057_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21011_ _21009_/X _21010_/X _20262_/X VGND VGND VPWR VPWR _21011_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_82_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12541__A _12906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16013__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15120__A1 _15048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19398__B1 _19396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15852__A _13542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19324__A _19324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22962_ _18548_/X _22938_/B VGND VGND VPWR VPWR _22963_/C sky130_fd_sc_hd__or2_4
XFILLER_114_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17948__A1 _17813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21744__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21913_ _21906_/A VGND VGND VPWR VPWR _21913_/X sky130_fd_sc_hd__buf_2
XFILLER_167_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14468__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22893_ _17261_/Y _22885_/X _22875_/X _22892_/X VGND VGND VPWR VPWR _22894_/B sky130_fd_sc_hd__o22a_4
XANTENNA__13372__A _13413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21844_ _21843_/X _21839_/X _23623_/Q _21834_/X VGND VGND VPWR VPWR _21844_/X sky130_fd_sc_hd__o22a_4
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21775_ _21548_/X _21770_/X _12672_/B _21774_/X VGND VGND VPWR VPWR _21775_/X sky130_fd_sc_hd__o22a_4
XFILLER_130_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16683__A _16683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20917__B _20917_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20726_ _20490_/A VGND VGND VPWR VPWR _20726_/X sky130_fd_sc_hd__buf_2
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23514_ _24090_/CLK _23514_/D VGND VGND VPWR VPWR _23514_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24494_ _24306_/CLK _24494_/D HRESETn VGND VGND VPWR VPWR _20008_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15299__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20657_ _24228_/Q _20636_/X _20656_/Y VGND VGND VPWR VPWR _20658_/A sky130_fd_sc_hd__o21a_4
XANTENNA__19994__A _19950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23445_ _23392_/CLK _23445_/D VGND VGND VPWR VPWR _23445_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12716__A _11970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11620__A _13792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23959__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23376_ _23760_/CLK _22285_/X VGND VGND VPWR VPWR _16390_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_137_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20588_ _20501_/A _20587_/X VGND VGND VPWR VPWR _20588_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22327_ _16266_/B VGND VGND VPWR VPWR _23343_/D sky130_fd_sc_hd__buf_2
XANTENNA__21680__B2 _21674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14931__A _11752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13060_ _13095_/A _23752_/Q VGND VGND VPWR VPWR _13061_/C sky130_fd_sc_hd__or2_4
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22258_ _22258_/A VGND VGND VPWR VPWR _22258_/X sky130_fd_sc_hd__buf_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12011_ _11960_/A _23124_/Q VGND VGND VPWR VPWR _12013_/B sky130_fd_sc_hd__or2_4
XANTENNA__13547__A _13547_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21209_ _21202_/A VGND VGND VPWR VPWR _21209_/X sky130_fd_sc_hd__buf_2
XANTENNA__21432__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22189_ _22113_/X _22187_/X _16219_/B _22184_/X VGND VGND VPWR VPWR _22189_/X sky130_fd_sc_hd__o22a_4
XFILLER_160_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21983__A2 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23339__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16750_ _12027_/X _11632_/X _16719_/X _11609_/X _16749_/X VGND VGND VPWR VPWR _16821_/A
+ sky130_fd_sc_hd__a32o_4
X_13962_ _13985_/A _13960_/X _13962_/C VGND VGND VPWR VPWR _13966_/B sky130_fd_sc_hd__and3_4
XFILLER_24_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21735__A2 _21734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15701_ _13303_/A _15701_/B VGND VGND VPWR VPWR _15701_/X sky130_fd_sc_hd__or2_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12913_ _13453_/A _12890_/X _12897_/X _12904_/X _12912_/X VGND VGND VPWR VPWR _12913_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_24_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18061__B1 _18060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16681_ _16659_/A _16679_/X _16681_/C VGND VGND VPWR VPWR _16681_/X sky130_fd_sc_hd__and3_4
X_13893_ _14348_/A _13893_/B _13893_/C VGND VGND VPWR VPWR _13894_/C sky130_fd_sc_hd__or3_4
XANTENNA__24367__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13282__A _12516_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18420_ _17396_/A _18419_/X _17445_/Y VGND VGND VPWR VPWR _18420_/X sky130_fd_sc_hd__o21a_4
X_15632_ _15616_/A _15628_/X _15632_/C VGND VGND VPWR VPWR _15632_/X sky130_fd_sc_hd__or3_4
XFILLER_34_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12844_ _12753_/Y _12842_/X VGND VGND VPWR VPWR _12845_/A sky130_fd_sc_hd__or2_4
XANTENNA__19888__B _19888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18351_ _18330_/X _18332_/X _18219_/X _18350_/X VGND VGND VPWR VPWR _18351_/X sky130_fd_sc_hd__o22a_4
X_15563_ _11900_/A _15563_/B VGND VGND VPWR VPWR _15563_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_23_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12775_ _12775_/A _23786_/Q VGND VGND VPWR VPWR _12775_/X sky130_fd_sc_hd__or2_4
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _14549_/Y _17302_/B VGND VGND VPWR VPWR _17632_/A sky130_fd_sc_hd__or2_4
XANTENNA__22160__A2 _22159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _11781_/A _14505_/X _14514_/C VGND VGND VPWR VPWR _14514_/X sky130_fd_sc_hd__and3_4
XFILLER_15_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _12370_/A VGND VGND VPWR VPWR _11727_/A sky130_fd_sc_hd__buf_2
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18282_ _18282_/A _18282_/B VGND VGND VPWR VPWR _18283_/D sky130_fd_sc_hd__and2_4
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _13742_/A _15494_/B VGND VGND VPWR VPWR _15495_/C sky130_fd_sc_hd__or2_4
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21004__A _21313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17233_ _17233_/A VGND VGND VPWR VPWR _17233_/X sky130_fd_sc_hd__buf_2
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14445_ _12445_/A _14445_/B _14445_/C VGND VGND VPWR VPWR _14445_/X sky130_fd_sc_hd__and3_4
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _11706_/A VGND VGND VPWR VPWR _14772_/A sky130_fd_sc_hd__buf_2
XANTENNA__12626__A _12626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15002__A _13965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17164_ _17164_/A VGND VGND VPWR VPWR _17838_/A sky130_fd_sc_hd__buf_2
X_14376_ _14516_/A _14376_/B VGND VGND VPWR VPWR _14376_/X sky130_fd_sc_hd__or2_4
XANTENNA__20843__A HRDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11588_ _11643_/A VGND VGND VPWR VPWR _17091_/A sky130_fd_sc_hd__buf_2
XANTENNA__12345__B _23788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16115_ _16147_/A _24013_/Q VGND VGND VPWR VPWR _16116_/C sky130_fd_sc_hd__or2_4
XFILLER_128_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13327_ _13327_/A _13325_/X _13326_/X VGND VGND VPWR VPWR _13331_/B sky130_fd_sc_hd__and3_4
XANTENNA__21671__B2 _21667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17095_ _17094_/Y VGND VGND VPWR VPWR _17095_/X sky130_fd_sc_hd__buf_2
XANTENNA__14841__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19427__A2_N _18633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16046_ _16046_/A _24014_/Q VGND VGND VPWR VPWR _16047_/C sky130_fd_sc_hd__or2_4
X_13258_ _13258_/A _13258_/B _13258_/C VGND VGND VPWR VPWR _13259_/C sky130_fd_sc_hd__or3_4
XANTENNA__14560__B _14560_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13457__A _13327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12209_ _12693_/A _12344_/B VGND VGND VPWR VPWR _12211_/B sky130_fd_sc_hd__or2_4
XFILLER_124_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13189_ _11872_/A _13189_/B _13189_/C VGND VGND VPWR VPWR _13189_/X sky130_fd_sc_hd__or3_4
XANTENNA__21674__A _21674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19805_ _19441_/X _19804_/X _16659_/A _19700_/X VGND VGND VPWR VPWR _19805_/X sky130_fd_sc_hd__o22a_4
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17997_ _17985_/X _17948_/X _17877_/X _17996_/Y VGND VGND VPWR VPWR _17997_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16768__A _16768_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19736_ _19528_/A _19665_/A _19622_/B _19705_/A _19787_/A VGND VGND VPWR VPWR _19736_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24264__CLK _24271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16948_ _16948_/A VGND VGND VPWR VPWR _17659_/A sky130_fd_sc_hd__inv_2
XFILLER_56_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21726__A2 _21720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_105_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR _23750_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19667_ _19642_/A VGND VGND VPWR VPWR _19879_/C sky130_fd_sc_hd__buf_2
X_16879_ _16830_/X _16831_/B _16830_/X _16831_/B VGND VGND VPWR VPWR _16880_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14288__A _12470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16602__A1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18618_ _18615_/Y _22943_/B _18615_/Y _22943_/B VGND VGND VPWR VPWR _18618_/X sky130_fd_sc_hd__a2bb2o_4
X_19598_ _19560_/A VGND VGND VPWR VPWR _19661_/A sky130_fd_sc_hd__inv_2
XFILLER_64_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18549_ _18477_/X _18537_/Y _18504_/X _18548_/X VGND VGND VPWR VPWR _18549_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13920__A _14348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21560_ _21560_/A VGND VGND VPWR VPWR _21560_/X sky130_fd_sc_hd__buf_2
XFILLER_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20511_ _20418_/X _20509_/X _12669_/B _20510_/X VGND VGND VPWR VPWR _20511_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21491_ _21266_/X _21485_/X _12825_/B _21489_/X VGND VGND VPWR VPWR _23818_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16008__A _16007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23230_ _23646_/CLK _22524_/X VGND VGND VPWR VPWR _13775_/B sky130_fd_sc_hd__dfxtp_4
X_20442_ _20418_/X _20441_/X _24110_/Q _20396_/X VGND VGND VPWR VPWR _24110_/D sky130_fd_sc_hd__o22a_4
XFILLER_118_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23161_ _23641_/CLK _23161_/D VGND VGND VPWR VPWR _14798_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_173_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15847__A _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19319__A _24129_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20373_ _20373_/A VGND VGND VPWR VPWR _20373_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14751__A _15447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18223__A _18335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22112_ _22110_/X _22111_/X _23470_/Q _22106_/X VGND VGND VPWR VPWR _22112_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23092_ _17060_/A VGND VGND VPWR VPWR HSIZE[1] sky130_fd_sc_hd__buf_2
XFILLER_133_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13367__A _13367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22043_ _22042_/X VGND VGND VPWR VPWR _22043_/X sky130_fd_sc_hd__buf_2
XANTENNA__21414__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21965__A2 _21960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21584__A _20860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16678__A _16678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21178__B1 _14721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23994_ _24057_/CLK _23994_/D VGND VGND VPWR VPWR _14568_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_21_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22945_ _22945_/A _22942_/X _22945_/C VGND VGND VPWR VPWR HADDR[7] sky130_fd_sc_hd__and3_4
XANTENNA__14198__A _11654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11615__A _11928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22876_ _19915_/X VGND VGND VPWR VPWR _22876_/X sky130_fd_sc_hd__buf_2
XFILLER_71_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21827_ _21839_/A VGND VGND VPWR VPWR _21827_/X sky130_fd_sc_hd__buf_2
XANTENNA__22678__B1 _14523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14926__A _14772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19543__B1 HRDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17302__A _14549_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12560_ _12569_/A VGND VGND VPWR VPWR _12561_/A sky130_fd_sc_hd__buf_2
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20153__A1 _19906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21758_ _21791_/A VGND VGND VPWR VPWR _21774_/A sky130_fd_sc_hd__inv_2
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11511_ _11511_/A VGND VGND VPWR VPWR _19957_/A sky130_fd_sc_hd__inv_2
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20709_ _20516_/X _20707_/X _11528_/A _20708_/X VGND VGND VPWR VPWR _20709_/X sky130_fd_sc_hd__o22a_4
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12571_/A VGND VGND VPWR VPWR _12516_/A sky130_fd_sc_hd__buf_2
X_24477_ _24137_/CLK _24477_/D HRESETn VGND VGND VPWR VPWR _20088_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21689_ _21572_/X _21684_/X _23713_/Q _21688_/X VGND VGND VPWR VPWR _21689_/X sky130_fd_sc_hd__o22a_4
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _14623_/A _23615_/Q VGND VGND VPWR VPWR _14230_/X sky130_fd_sc_hd__or2_4
XFILLER_138_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23428_ _23588_/CLK _23428_/D VGND VGND VPWR VPWR _15698_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21102__B1 _12608_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24137__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20663__A _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15757__A _12778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14161_ _14267_/A _23231_/Q VGND VGND VPWR VPWR _14161_/X sky130_fd_sc_hd__or2_4
XFILLER_153_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21653__B2 _21617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23359_ _23582_/CLK _23359_/D VGND VGND VPWR VPWR _23359_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14661__A _13928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13112_ _13088_/A _23720_/Q VGND VGND VPWR VPWR _13114_/B sky130_fd_sc_hd__or2_4
X_14092_ _14003_/A _14092_/B _14092_/C VGND VGND VPWR VPWR _14100_/B sky130_fd_sc_hd__and3_4
XANTENNA__13277__A _13277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13043_ _12512_/A _23880_/Q VGND VGND VPWR VPWR _13044_/C sky130_fd_sc_hd__or2_4
XANTENNA__17972__A _17793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17920_ _17919_/X VGND VGND VPWR VPWR _17920_/X sky130_fd_sc_hd__buf_2
XANTENNA__12181__A _12180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24287__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21956__A2 _21953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17851_ _17837_/X _17194_/X _17838_/X _17196_/X VGND VGND VPWR VPWR _17851_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16802_ _16786_/A _16794_/X _16801_/X VGND VGND VPWR VPWR _16818_/B sky130_fd_sc_hd__and3_4
X_17782_ _17781_/X VGND VGND VPWR VPWR _17782_/Y sky130_fd_sc_hd__inv_2
X_14994_ _14994_/A _23765_/Q VGND VGND VPWR VPWR _14995_/C sky130_fd_sc_hd__or2_4
XFILLER_94_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19521_ _19509_/X VGND VGND VPWR VPWR _19521_/Y sky130_fd_sc_hd__inv_2
X_16733_ _16561_/A _16733_/B _16733_/C VGND VGND VPWR VPWR _16733_/X sky130_fd_sc_hd__or3_4
X_13945_ _11668_/A _13945_/B _13945_/C VGND VGND VPWR VPWR _13945_/X sky130_fd_sc_hd__and3_4
XANTENNA__17388__A2 _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22381__A2 _22376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19782__B1 _16683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19452_ _17005_/X _24128_/Q VGND VGND VPWR VPWR _19452_/X sky130_fd_sc_hd__or2_4
XFILLER_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16664_ _16676_/A _16664_/B VGND VGND VPWR VPWR _16664_/X sky130_fd_sc_hd__or2_4
XFILLER_90_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13876_ _14386_/A _13876_/B VGND VGND VPWR VPWR _13876_/X sky130_fd_sc_hd__or2_4
XFILLER_46_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18403_ _18402_/A _18403_/B VGND VGND VPWR VPWR _22990_/C sky130_fd_sc_hd__and2_4
XFILLER_62_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15615_ _13886_/A _15615_/B _15615_/C VGND VGND VPWR VPWR _15616_/C sky130_fd_sc_hd__and3_4
X_12827_ _12827_/A VGND VGND VPWR VPWR _13387_/A sky130_fd_sc_hd__buf_2
X_19383_ _17008_/A _17009_/B _18148_/A VGND VGND VPWR VPWR _19383_/X sky130_fd_sc_hd__o21a_4
X_16595_ _16595_/A _16593_/X _16594_/X VGND VGND VPWR VPWR _16599_/B sky130_fd_sc_hd__and3_4
XFILLER_90_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22133__A2 _22123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18334_ _18406_/A _18334_/B VGND VGND VPWR VPWR _18337_/B sky130_fd_sc_hd__and2_4
XFILLER_91_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15546_ _12434_/A _15546_/B VGND VGND VPWR VPWR _15548_/B sky130_fd_sc_hd__or2_4
X_12758_ _12758_/A VGND VGND VPWR VPWR _12759_/A sky130_fd_sc_hd__buf_2
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18265_ _18265_/A VGND VGND VPWR VPWR _18265_/X sky130_fd_sc_hd__buf_2
X_11709_ _13866_/A VGND VGND VPWR VPWR _11710_/A sky130_fd_sc_hd__buf_2
X_15477_ _15477_/A _15477_/B VGND VGND VPWR VPWR _15479_/B sky130_fd_sc_hd__or2_4
XFILLER_129_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12689_ _12689_/A _12768_/B VGND VGND VPWR VPWR _12691_/B sky130_fd_sc_hd__or2_4
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17216_ _17114_/X _17214_/X _17119_/X _17215_/X VGND VGND VPWR VPWR _17216_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14428_ _12546_/A _14423_/X _14427_/X VGND VGND VPWR VPWR _14428_/X sky130_fd_sc_hd__or3_4
XFILLER_163_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18196_ _17095_/X _18196_/B _18196_/C _18196_/D VGND VGND VPWR VPWR _18197_/A sky130_fd_sc_hd__or4_4
XANTENNA__15667__A _12727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17147_ _13947_/X _17144_/X _17145_/Y _17146_/X VGND VGND VPWR VPWR _17147_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21644__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14359_ _14366_/A _14359_/B VGND VGND VPWR VPWR _14359_/X sky130_fd_sc_hd__or2_4
XANTENNA__14571__A _15423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17078_ _11643_/A _17077_/A _17078_/C _18888_/B VGND VGND VPWR VPWR _17078_/X sky130_fd_sc_hd__or4_4
XFILLER_118_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16029_ _16056_/A _16027_/X _16029_/C VGND VGND VPWR VPWR _16029_/X sky130_fd_sc_hd__and3_4
XANTENNA__13187__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21947__A2 _21946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19719_ _19719_/A VGND VGND VPWR VPWR _19719_/X sky130_fd_sc_hd__buf_2
X_20991_ _20447_/A _20987_/X _20989_/X _20990_/Y _20495_/A VGND VGND VPWR VPWR _20992_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_77_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22372__A2 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22730_ _21304_/A _22729_/X _14604_/B _22726_/X VGND VGND VPWR VPWR _23098_/D sky130_fd_sc_hd__o22a_4
XFILLER_93_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24350__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22661_ _22442_/X _22658_/X _13237_/B _22655_/X VGND VGND VPWR VPWR _23143_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22124__A2 _22123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13650__A _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20467__B _20844_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24400_ _23281_/CLK _18905_/X HRESETn VGND VGND VPWR VPWR _24400_/Q sky130_fd_sc_hd__dfstp_4
X_21612_ _21608_/A VGND VGND VPWR VPWR _21620_/A sky130_fd_sc_hd__buf_2
X_22592_ _22586_/Y _22591_/X _22410_/X _22591_/X VGND VGND VPWR VPWR _22592_/X sky130_fd_sc_hd__a2bb2o_4
X_24331_ _24277_/CLK _24331_/D HRESETn VGND VGND VPWR VPWR _24331_/Q sky130_fd_sc_hd__dfrtp_4
X_21543_ _21541_/X _21542_/X _23790_/Q _21537_/X VGND VGND VPWR VPWR _23790_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12266__A _12266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21474_ _21489_/A VGND VGND VPWR VPWR _21482_/A sky130_fd_sc_hd__buf_2
X_24262_ _24127_/CLK _24262_/D HRESETn VGND VGND VPWR VPWR _20608_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20483__A _20438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11601__C _17048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19694__D _19687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23213_ _24045_/CLK _22553_/X VGND VGND VPWR VPWR _16177_/B sky130_fd_sc_hd__dfxtp_4
X_20425_ _20425_/A VGND VGND VPWR VPWR _20425_/X sky130_fd_sc_hd__buf_2
XANTENNA__15577__A _14270_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21635__B2 _21631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24193_ _23383_/CLK _24193_/D HRESETn VGND VGND VPWR VPWR _17060_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_49_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23144_ _23496_/CLK _22660_/X VGND VGND VPWR VPWR _13025_/B sky130_fd_sc_hd__dfxtp_4
X_20356_ _24274_/Q VGND VGND VPWR VPWR _20356_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18888__A _11609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23075_ _23080_/A _23075_/B _23074_/X VGND VGND VPWR VPWR _23075_/X sky130_fd_sc_hd__and3_4
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20287_ _20287_/A VGND VGND VPWR VPWR _20343_/A sky130_fd_sc_hd__buf_2
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17067__A1 _18782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22026_ _21865_/X _22024_/X _13707_/B _22021_/X VGND VGND VPWR VPWR _23518_/D sky130_fd_sc_hd__o22a_4
XFILLER_49_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13825__A _13666_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16201__A _16163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23977_ _24073_/CLK _23977_/D VGND VGND VPWR VPWR _23977_/Q sky130_fd_sc_hd__dfxtp_4
X_11991_ _11943_/X _11991_/B _11990_/X VGND VGND VPWR VPWR _11992_/C sky130_fd_sc_hd__and3_4
XFILLER_5_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22363__A2 _22362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13730_ _13756_/A _13723_/X _13730_/C VGND VGND VPWR VPWR _13730_/X sky130_fd_sc_hd__or3_4
XFILLER_21_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22928_ _22927_/X VGND VGND VPWR VPWR HADDR[4] sky130_fd_sc_hd__inv_2
XANTENNA__21571__B1 _23778_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20658__A _20658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13661_ _11933_/A _13661_/B _13661_/C VGND VGND VPWR VPWR _13661_/X sky130_fd_sc_hd__or3_4
X_22859_ _22859_/A VGND VGND VPWR VPWR HWDATA[18] sky130_fd_sc_hd__inv_2
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14656__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15400_ _15400_/A _23778_/Q VGND VGND VPWR VPWR _15401_/C sky130_fd_sc_hd__or2_4
X_12612_ _12953_/A _12612_/B _12611_/X VGND VGND VPWR VPWR _12613_/C sky130_fd_sc_hd__and3_4
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16380_ _13417_/A _16346_/X _16379_/X VGND VGND VPWR VPWR _16380_/X sky130_fd_sc_hd__and3_4
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13592_ _13965_/A VGND VGND VPWR VPWR _13593_/A sky130_fd_sc_hd__buf_2
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15331_ _15377_/A _15331_/B _15331_/C VGND VGND VPWR VPWR _15347_/B sky130_fd_sc_hd__and3_4
X_12543_ _12903_/A _12543_/B _12543_/C VGND VGND VPWR VPWR _12544_/C sky130_fd_sc_hd__and3_4
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17967__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18050_ _17873_/X _18047_/X _17847_/A _18049_/X VGND VGND VPWR VPWR _18051_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21489__A _21489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15262_ _14103_/A _15262_/B _15262_/C VGND VGND VPWR VPWR _15262_/X sky130_fd_sc_hd__and3_4
XANTENNA__17686__B _17511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12474_ _12474_/A VGND VGND VPWR VPWR _13642_/A sky130_fd_sc_hd__buf_2
XANTENNA__16750__B1 _11609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17001_ _16945_/X _16999_/B _17000_/Y VGND VGND VPWR VPWR _23073_/B sky130_fd_sc_hd__a21o_4
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14213_ _13882_/A _14213_/B _14212_/X VGND VGND VPWR VPWR _14213_/X sky130_fd_sc_hd__or3_4
XANTENNA__21626__B2 _21624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15193_ _14773_/A _15129_/B VGND VGND VPWR VPWR _15195_/B sky130_fd_sc_hd__or2_4
XANTENNA__14391__A _14510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12904__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20834__C1 _20833_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14144_ _14137_/A _23135_/Q VGND VGND VPWR VPWR _14144_/X sky130_fd_sc_hd__or2_4
XFILLER_152_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18952_ _24403_/Q VGND VGND VPWR VPWR _18952_/Y sky130_fd_sc_hd__inv_2
X_14075_ _14075_/A _23488_/Q VGND VGND VPWR VPWR _14075_/X sky130_fd_sc_hd__or2_4
XFILLER_106_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21929__A2 _21923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13026_ _12506_/A _23848_/Q VGND VGND VPWR VPWR _13027_/C sky130_fd_sc_hd__or2_4
X_17903_ _17903_/A _17902_/Y VGND VGND VPWR VPWR _17908_/A sky130_fd_sc_hd__or2_4
XANTENNA__22051__B2 _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18948__D _18948_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18883_ _15251_/A _18877_/X _24407_/Q _18878_/X VGND VGND VPWR VPWR _24407_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22113__A _22113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13735__A _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17834_ _17825_/A VGND VGND VPWR VPWR _17922_/A sky130_fd_sc_hd__buf_2
XANTENNA__16111__A _16138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17765_ _18478_/A _17360_/X _17717_/X _17764_/X VGND VGND VPWR VPWR _17765_/X sky130_fd_sc_hd__o22a_4
X_14977_ _15076_/A _23638_/Q VGND VGND VPWR VPWR _14978_/C sky130_fd_sc_hd__or2_4
XFILLER_82_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19504_ _19624_/A _19504_/B VGND VGND VPWR VPWR _19560_/A sky130_fd_sc_hd__or2_4
XFILLER_75_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16716_ _16595_/A _16714_/X _16715_/X VGND VGND VPWR VPWR _16716_/X sky130_fd_sc_hd__and3_4
X_13928_ _13928_/A _13928_/B _13927_/X VGND VGND VPWR VPWR _13944_/B sky130_fd_sc_hd__and3_4
X_17696_ _17693_/X _17694_/X _17772_/A VGND VGND VPWR VPWR _17696_/X sky130_fd_sc_hd__a21o_4
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16647_ _16647_/A VGND VGND VPWR VPWR _16678_/A sky130_fd_sc_hd__buf_2
X_19435_ _18670_/X _24213_/Q _19399_/X _24131_/Q VGND VGND VPWR VPWR _24213_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24302__CLK _24302_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13859_ _12251_/A _13859_/B _13859_/C VGND VGND VPWR VPWR _13859_/X sky130_fd_sc_hd__and3_4
XANTENNA__14566__A _14310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13470__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19366_ _19362_/X _18550_/X _19365_/X _24255_/Q VGND VGND VPWR VPWR _24255_/D sky130_fd_sc_hd__a2bb2o_4
X_16578_ _16558_/A _16661_/B VGND VGND VPWR VPWR _16578_/X sky130_fd_sc_hd__or2_4
XFILLER_128_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15529_ _12239_/A _23201_/Q VGND VGND VPWR VPWR _15529_/X sky130_fd_sc_hd__or2_4
X_18317_ _17874_/X _18316_/X _18200_/X _17881_/X VGND VGND VPWR VPWR _18318_/A sky130_fd_sc_hd__o22a_4
X_19297_ _19237_/X VGND VGND VPWR VPWR _19297_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18248_ _17009_/A _17906_/C _18248_/C VGND VGND VPWR VPWR _18248_/X sky130_fd_sc_hd__and3_4
XFILLER_124_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15397__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18179_ _17963_/X _18149_/X _18033_/X _18178_/X VGND VGND VPWR VPWR _18179_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12814__A _13343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20210_ _24116_/Q VGND VGND VPWR VPWR _20210_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21093__A2 _21090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21190_ _21219_/A VGND VGND VPWR VPWR _21198_/A sky130_fd_sc_hd__buf_2
XFILLER_171_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22290__B2 _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12533__B _12533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20141_ _11557_/X _20139_/X _20140_/Y VGND VGND VPWR VPWR _20141_/X sky130_fd_sc_hd__o21a_4
XFILLER_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20072_ _18497_/X _20055_/X _20071_/Y _20066_/X VGND VGND VPWR VPWR _20072_/X sky130_fd_sc_hd__o22a_4
XFILLER_83_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23900_ _23515_/CLK _21360_/X VGND VGND VPWR VPWR _14376_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_100_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13645__A _11913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22958__A _22957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23831_ _23862_/CLK _23831_/D VGND VGND VPWR VPWR _15227_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21862__A _20801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18549__B2 _18548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23762_ _23728_/CLK _21615_/X VGND VGND VPWR VPWR _23762_/Q sky130_fd_sc_hd__dfxtp_4
X_20974_ _18717_/X _20342_/X _20662_/X _20973_/Y VGND VGND VPWR VPWR _20974_/X sky130_fd_sc_hd__a211o_4
XPHY_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22713_ _21560_/A _22708_/X _23110_/Q _22712_/X VGND VGND VPWR VPWR _23110_/D sky130_fd_sc_hd__o22a_4
XFILLER_26_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23693_ _23501_/CLK _21722_/X VGND VGND VPWR VPWR _16199_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13380__A _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22644_ _22658_/A VGND VGND VPWR VPWR _22644_/X sky130_fd_sc_hd__buf_2
XFILLER_94_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14195__B _23199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22693__A _22722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21856__B2 _21846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22575_ _22466_/X _22572_/X _13807_/B _22569_/X VGND VGND VPWR VPWR _23197_/D sky130_fd_sc_hd__o22a_4
XFILLER_142_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24314_ _24287_/CLK _19214_/X HRESETn VGND VGND VPWR VPWR _19135_/A sky130_fd_sc_hd__dfrtp_4
X_21526_ _21526_/A VGND VGND VPWR VPWR _21526_/X sky130_fd_sc_hd__buf_2
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24245_ _23126_/CLK _19382_/X HRESETn VGND VGND VPWR VPWR _24245_/Q sky130_fd_sc_hd__dfrtp_4
X_21457_ _21295_/X _21455_/X _13758_/B _21452_/X VGND VGND VPWR VPWR _21457_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12724__A _13279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12190_ _12190_/A VGND VGND VPWR VPWR _12191_/A sky130_fd_sc_hd__buf_2
X_20408_ _20313_/X _20407_/X VGND VGND VPWR VPWR _20408_/Y sky130_fd_sc_hd__nor2_4
X_21388_ _21388_/A VGND VGND VPWR VPWR _21388_/X sky130_fd_sc_hd__buf_2
X_24176_ _24184_/CLK _24176_/D HRESETn VGND VGND VPWR VPWR _24176_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22281__B2 _22277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_13_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR _24428_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11572__A2 IRQ[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23127_ _23862_/CLK _23127_/D VGND VGND VPWR VPWR _15162_/B sky130_fd_sc_hd__dfxtp_4
X_20339_ _18780_/X _20339_/B VGND VGND VPWR VPWR _20339_/X sky130_fd_sc_hd__and2_4
Xclkbuf_7_76_0_HCLK clkbuf_7_77_0_HCLK/A VGND VGND VPWR VPWR _23194_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18411__A _18411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18237__B1 _18176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23058_ _23058_/A VGND VGND VPWR VPWR HADDR[26] sky130_fd_sc_hd__inv_2
XANTENNA__22033__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14900_ _14897_/X _14898_/X _14900_/C VGND VGND VPWR VPWR _14901_/C sky130_fd_sc_hd__and3_4
XANTENNA__13555__A _12773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22009_ _21836_/X _22003_/X _12763_/B _22007_/X VGND VGND VPWR VPWR _23530_/D sky130_fd_sc_hd__o22a_4
XFILLER_62_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15880_ _13530_/A _15864_/X _15880_/C VGND VGND VPWR VPWR _15912_/B sky130_fd_sc_hd__or3_4
XFILLER_23_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21792__B1 _23647_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14831_ _14658_/A _14761_/B VGND VGND VPWR VPWR _14831_/X sky130_fd_sc_hd__or2_4
XANTENNA__24325__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17550_ _16452_/Y _17024_/X _17031_/X _17659_/B VGND VGND VPWR VPWR _17551_/B sky130_fd_sc_hd__o22a_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14762_ _12250_/A _14762_/B _14761_/X VGND VGND VPWR VPWR _14762_/X sky130_fd_sc_hd__and3_4
X_11974_ _16138_/A VGND VGND VPWR VPWR _16568_/A sky130_fd_sc_hd__buf_2
XANTENNA__16015__A2 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16501_ _16481_/X _16432_/B VGND VGND VPWR VPWR _16502_/C sky130_fd_sc_hd__or2_4
XANTENNA__17212__A1 _12680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13713_ _15487_/A _13713_/B VGND VGND VPWR VPWR _13713_/X sky130_fd_sc_hd__or2_4
X_17481_ _11876_/X _17481_/B VGND VGND VPWR VPWR _17481_/X sky130_fd_sc_hd__and2_4
XFILLER_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14693_ _14693_/A _14691_/X _14692_/X VGND VGND VPWR VPWR _14697_/B sky130_fd_sc_hd__and3_4
XANTENNA__14386__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16432_ _16409_/A _16432_/B VGND VGND VPWR VPWR _16432_/X sky130_fd_sc_hd__or2_4
XANTENNA__11803__A _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19220_ _24311_/Q _19131_/X _19219_/Y VGND VGND VPWR VPWR _19220_/X sky130_fd_sc_hd__o21a_4
XFILLER_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24475__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13644_ _12503_/A _13733_/B VGND VGND VPWR VPWR _13644_/X sky130_fd_sc_hd__or2_4
XANTENNA__19398__A1_N _19396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12618__B _12618_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19151_ _19151_/A _19151_/B VGND VGND VPWR VPWR _19151_/X sky130_fd_sc_hd__and2_4
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _16316_/A _16300_/B VGND VGND VPWR VPWR _16363_/X sky130_fd_sc_hd__or2_4
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21847__B2 _21846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _13574_/X VGND VGND VPWR VPWR _16832_/A sky130_fd_sc_hd__inv_2
X_18102_ _17963_/X _18073_/Y _18033_/X _18101_/X VGND VGND VPWR VPWR _18102_/X sky130_fd_sc_hd__o22a_4
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ _11708_/A _15253_/B VGND VGND VPWR VPWR _15317_/B sky130_fd_sc_hd__or2_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19082_ _18957_/X VGND VGND VPWR VPWR _19082_/X sky130_fd_sc_hd__buf_2
X_12526_ _12473_/A VGND VGND VPWR VPWR _13974_/A sky130_fd_sc_hd__buf_2
X_16294_ _11904_/X _16294_/B VGND VGND VPWR VPWR _16294_/X sky130_fd_sc_hd__or2_4
XFILLER_12_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22108__A _20415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18033_ _18032_/X VGND VGND VPWR VPWR _18033_/X sky130_fd_sc_hd__buf_2
X_15245_ _14248_/A _15173_/B VGND VGND VPWR VPWR _15246_/C sky130_fd_sc_hd__or2_4
X_12457_ _12885_/A _23755_/Q VGND VGND VPWR VPWR _12458_/C sky130_fd_sc_hd__or2_4
XFILLER_145_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12634__A _12634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16106__A _15969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21075__A2 _21073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15176_ _14988_/A _15176_/B VGND VGND VPWR VPWR _15176_/X sky130_fd_sc_hd__or2_4
X_12388_ _15887_/A _12384_/X _12388_/C VGND VGND VPWR VPWR _12396_/B sky130_fd_sc_hd__or3_4
XFILLER_113_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20283__B1 _24468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11563__A2 IRQ[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14127_ _14127_/A _23935_/Q VGND VGND VPWR VPWR _14129_/B sky130_fd_sc_hd__or2_4
X_19984_ _24499_/Q VGND VGND VPWR VPWR _19984_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18935_ _18928_/A VGND VGND VPWR VPWR _18935_/X sky130_fd_sc_hd__buf_2
X_14058_ _11753_/A _14054_/X _14057_/X VGND VGND VPWR VPWR _14058_/X sky130_fd_sc_hd__or3_4
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13465__A _13441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13009_ _12537_/A _23944_/Q VGND VGND VPWR VPWR _13009_/X sky130_fd_sc_hd__or2_4
XANTENNA__19976__B1 _17014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18866_ _15784_/X _18863_/X _24420_/Q _18864_/X VGND VGND VPWR VPWR _24420_/D sky130_fd_sc_hd__o22a_4
XFILLER_94_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17817_ _17817_/A VGND VGND VPWR VPWR _17817_/X sky130_fd_sc_hd__buf_2
XANTENNA__14265__A1 _14263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18797_ _18790_/A VGND VGND VPWR VPWR _18797_/X sky130_fd_sc_hd__buf_2
XFILLER_82_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15680__A _12279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20338__A1 _20302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17748_ _17748_/A _17321_/X VGND VGND VPWR VPWR _17748_/X sky130_fd_sc_hd__and2_4
XANTENNA__20338__B2 _20225_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20298__A _20298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17679_ _17679_/A _17699_/A VGND VGND VPWR VPWR _17683_/A sky130_fd_sc_hd__or2_4
XFILLER_39_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14296__A _14296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19418_ _19406_/X VGND VGND VPWR VPWR _19418_/X sky130_fd_sc_hd__buf_2
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20690_ _20535_/X _20690_/B VGND VGND VPWR VPWR _20690_/X sky130_fd_sc_hd__or2_4
X_19349_ _19347_/X _18242_/X _19347_/X _20526_/A VGND VGND VPWR VPWR _19349_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19900__B1 _16927_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22360_ _22354_/Y _22359_/X _22095_/X _22359_/X VGND VGND VPWR VPWR _23316_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14743__B _14743_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21311_ _21311_/A VGND VGND VPWR VPWR _21311_/X sky130_fd_sc_hd__buf_2
X_22291_ _22291_/A VGND VGND VPWR VPWR _22291_/X sky130_fd_sc_hd__buf_2
XANTENNA__12544__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24030_ _23880_/CLK _24030_/D VGND VGND VPWR VPWR _24030_/Q sky130_fd_sc_hd__dfxtp_4
X_21242_ _21233_/Y _21240_/X _21241_/X _21240_/X VGND VGND VPWR VPWR _23956_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22263__B2 _22262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12751__A1 _13307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21173_ _21152_/A VGND VGND VPWR VPWR _21173_/X sky130_fd_sc_hd__buf_2
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18231__A _18562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20124_ _20124_/A _20124_/B VGND VGND VPWR VPWR _20125_/B sky130_fd_sc_hd__or2_4
XANTENNA__22015__B2 _22014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20055_ _19961_/X VGND VGND VPWR VPWR _20055_/X sky130_fd_sc_hd__buf_2
XANTENNA__24288__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16245__A2 _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22318__A2 _22315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16686__A _16687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23814_ _23397_/CLK _21497_/X VGND VGND VPWR VPWR _23814_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _23908_/CLK _23745_/D VGND VGND VPWR VPWR _23745_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _24216_/Q _20895_/X _20956_/Y VGND VGND VPWR VPWR _20958_/A sky130_fd_sc_hd__o21a_4
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12719__A _12279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18942__A1 _16866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__A _11623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11689_/X VGND VGND VPWR VPWR _13399_/A sky130_fd_sc_hd__buf_2
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23676_ _23675_/CLK _23676_/D VGND VGND VPWR VPWR _14366_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _24251_/Q _20661_/X _20887_/X VGND VGND VPWR VPWR _20888_/X sky130_fd_sc_hd__o21a_4
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22627_ _22468_/X _22622_/X _14362_/B _22626_/X VGND VGND VPWR VPWR _23164_/D sky130_fd_sc_hd__o22a_4
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18406__A _18406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13360_ _13375_/A _23302_/Q VGND VGND VPWR VPWR _13361_/C sky130_fd_sc_hd__or2_4
XFILLER_158_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22558_ _22558_/A VGND VGND VPWR VPWR _22558_/X sky130_fd_sc_hd__buf_2
XFILLER_166_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12311_ _12311_/A _12399_/B VGND VGND VPWR VPWR _12312_/C sky130_fd_sc_hd__or2_4
XFILLER_158_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21509_ _21297_/X _21506_/X _13930_/B _21503_/X VGND VGND VPWR VPWR _23805_/D sky130_fd_sc_hd__o22a_4
X_13291_ _13303_/A VGND VGND VPWR VPWR _13319_/A sky130_fd_sc_hd__buf_2
X_22489_ _22489_/A VGND VGND VPWR VPWR _22505_/A sky130_fd_sc_hd__inv_2
XFILLER_6_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12454__A _12454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15030_ _13642_/A _23477_/Q VGND VGND VPWR VPWR _15030_/X sky130_fd_sc_hd__or2_4
XANTENNA__21057__A2 _21052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21767__A _21767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12242_ _12294_/A VGND VGND VPWR VPWR _12258_/A sky130_fd_sc_hd__buf_2
X_24228_ _24134_/CLK _19415_/X HRESETn VGND VGND VPWR VPWR _24228_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22254__B2 _22248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15765__A _11689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24159_ _24271_/CLK _24159_/D HRESETn VGND VGND VPWR VPWR _24159_/Q sky130_fd_sc_hd__dfrtp_4
X_12173_ _12166_/A _12173_/B VGND VGND VPWR VPWR _12173_/X sky130_fd_sc_hd__or2_4
XFILLER_174_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22006__B2 _22000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16981_ _16981_/A _16980_/X VGND VGND VPWR VPWR _16981_/X sky130_fd_sc_hd__or2_4
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22557__A2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18720_ _16940_/Y _18717_/X _16939_/X _18719_/X VGND VGND VPWR VPWR _18720_/Y sky130_fd_sc_hd__a22oi_4
X_15932_ _15932_/A _13580_/Y _15932_/C VGND VGND VPWR VPWR _15933_/A sky130_fd_sc_hd__and3_4
XFILLER_118_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22598__A _22598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_6_0_HCLK clkbuf_7_6_0_HCLK/A VGND VGND VPWR VPWR _24357_/CLK sky130_fd_sc_hd__clkbuf_1
X_15863_ _15887_/A _15859_/X _15863_/C VGND VGND VPWR VPWR _15863_/X sky130_fd_sc_hd__or3_4
X_18651_ _18483_/A _18651_/B VGND VGND VPWR VPWR _18651_/Y sky130_fd_sc_hd__nor2_4
XFILLER_49_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22309__A2 _22308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14814_ _14667_/A _14812_/X _14813_/X VGND VGND VPWR VPWR _14814_/X sky130_fd_sc_hd__and3_4
X_17602_ _17522_/X _17601_/X _17515_/X _17524_/X VGND VGND VPWR VPWR _17603_/B sky130_fd_sc_hd__a211o_4
X_15794_ _13324_/A _15792_/X _15793_/X VGND VGND VPWR VPWR _15795_/C sky130_fd_sc_hd__and3_4
XFILLER_18_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18582_ _17436_/A _18581_/X VGND VGND VPWR VPWR _18582_/X sky130_fd_sc_hd__or2_4
XANTENNA__21517__B1 _15177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17533_ _13262_/X _17522_/B VGND VGND VPWR VPWR _17533_/Y sky130_fd_sc_hd__nand2_4
X_14745_ _12469_/A _14743_/X _14744_/X VGND VGND VPWR VPWR _14745_/X sky130_fd_sc_hd__and3_4
X_11957_ _11951_/X _11957_/B _11957_/C VGND VGND VPWR VPWR _11964_/B sky130_fd_sc_hd__and3_4
XFILLER_45_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12629__A _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18933__A1 _17272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17464_ _17046_/A _17463_/X _17418_/A VGND VGND VPWR VPWR _17464_/X sky130_fd_sc_hd__o21a_4
X_14676_ _14676_/A _14674_/X _14676_/C VGND VGND VPWR VPWR _14676_/X sky130_fd_sc_hd__and3_4
X_11888_ _11888_/A VGND VGND VPWR VPWR _13455_/A sky130_fd_sc_hd__buf_2
XANTENNA__20740__A1 _20662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16415_ _16401_/X _16415_/B VGND VGND VPWR VPWR _16415_/X sky130_fd_sc_hd__or2_4
X_19203_ _19141_/B VGND VGND VPWR VPWR _19203_/Y sky130_fd_sc_hd__inv_2
X_13627_ _13627_/A VGND VGND VPWR VPWR _13628_/A sky130_fd_sc_hd__buf_2
X_17395_ _17609_/D VGND VGND VPWR VPWR _17396_/D sky130_fd_sc_hd__inv_2
XANTENNA__14844__A _14843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16346_ _13383_/A _16328_/X _16345_/X VGND VGND VPWR VPWR _16346_/X sky130_fd_sc_hd__or3_4
X_19134_ _19134_/A _19133_/X VGND VGND VPWR VPWR _19215_/A sky130_fd_sc_hd__and2_4
X_13558_ _13546_/A _13470_/B VGND VGND VPWR VPWR _13558_/X sky130_fd_sc_hd__or2_4
XANTENNA__21296__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12509_ _13042_/A VGND VGND VPWR VPWR _12510_/A sky130_fd_sc_hd__buf_2
X_19065_ _19063_/Y _19064_/Y _11528_/B VGND VGND VPWR VPWR _19065_/X sky130_fd_sc_hd__o21a_4
X_16277_ _11971_/X _16276_/X VGND VGND VPWR VPWR _16277_/X sky130_fd_sc_hd__and2_4
XFILLER_145_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13489_ _12923_/A VGND VGND VPWR VPWR _13532_/A sky130_fd_sc_hd__buf_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21048__A2 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18016_ _17663_/X _18015_/X _17663_/X _18015_/X VGND VGND VPWR VPWR _18016_/X sky130_fd_sc_hd__a2bb2o_4
X_15228_ _14771_/A _15226_/X _15227_/X VGND VGND VPWR VPWR _15228_/X sky130_fd_sc_hd__and3_4
XANTENNA__22245__B2 _22241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21677__A _21677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15675__A _13145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15159_ _15294_/A _15223_/B VGND VGND VPWR VPWR _15159_/X sky130_fd_sc_hd__or2_4
XFILLER_153_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17121__B1 _17120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19967_ _19966_/X VGND VGND VPWR VPWR _19967_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13195__A _13230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11708__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18918_ _13262_/X _18913_/X _19032_/A _18914_/X VGND VGND VPWR VPWR _24391_/D sky130_fd_sc_hd__o22a_4
X_19898_ _19889_/A _19898_/B VGND VGND VPWR VPWR _19898_/X sky130_fd_sc_hd__or2_4
XFILLER_110_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18849_ _18840_/A VGND VGND VPWR VPWR _18849_/X sky130_fd_sc_hd__buf_2
XANTENNA__24310__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22301__A _22294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13923__A _13923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21860_ _20770_/A VGND VGND VPWR VPWR _21860_/X sky130_fd_sc_hd__buf_2
XANTENNA__21508__B1 _13766_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20811_ _20754_/X _20810_/X _24318_/Q _20761_/X VGND VGND VPWR VPWR _20812_/B sky130_fd_sc_hd__o22a_4
XFILLER_70_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21791_ _21791_/A VGND VGND VPWR VPWR _21791_/X sky130_fd_sc_hd__buf_2
XANTENNA__18924__A1 _15916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22720__A2 _22715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23530_ _23531_/CLK _23530_/D VGND VGND VPWR VPWR _12763_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20742_ _20535_/X _20741_/X VGND VGND VPWR VPWR _20742_/X sky130_fd_sc_hd__or2_4
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23461_ _23397_/CLK _23461_/D VGND VGND VPWR VPWR _13518_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20673_ _20845_/A _20669_/X _20673_/C VGND VGND VPWR VPWR _20673_/X sky130_fd_sc_hd__and3_4
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14754__A _12294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22412_ _20336_/A VGND VGND VPWR VPWR _22412_/X sky130_fd_sc_hd__buf_2
XFILLER_149_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23392_ _23392_/CLK _22257_/X VGND VGND VPWR VPWR _14062_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_104_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22343_ _14117_/B VGND VGND VPWR VPWR _22343_/X sky130_fd_sc_hd__buf_2
XFILLER_148_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21039__A2 _21038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21587__A _20892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22236__B2 _22234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22274_ _22273_/X VGND VGND VPWR VPWR _22275_/A sky130_fd_sc_hd__buf_2
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24170__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24013_ _24077_/CLK _21150_/X VGND VGND VPWR VPWR _24013_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_151_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21225_ _20892_/X _21219_/X _23963_/Q _21223_/X VGND VGND VPWR VPWR _21225_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15585__A _14647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21156_ _20559_/X _21155_/X _24009_/Q _21152_/X VGND VGND VPWR VPWR _21156_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20107_ _19906_/X _20106_/X _19325_/X _17738_/X VGND VGND VPWR VPWR _20107_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__11618__A _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21087_ _21086_/X VGND VGND VPWR VPWR _21087_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21211__A2 _21205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20038_ _20016_/X _17686_/A _20022_/X _20037_/X VGND VGND VPWR VPWR _20038_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12860_ _12860_/A _23785_/Q VGND VGND VPWR VPWR _12861_/C sky130_fd_sc_hd__or2_4
XFILLER_100_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11811_ _15378_/A VGND VGND VPWR VPWR _11812_/A sky130_fd_sc_hd__buf_2
X_12791_ _12773_/X _12789_/X _12790_/X VGND VGND VPWR VPWR _12791_/X sky130_fd_sc_hd__and3_4
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12449__A _12863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21989_ _21706_/A _21656_/B _21706_/C _21030_/A VGND VGND VPWR VPWR _21990_/A sky130_fd_sc_hd__or4_4
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18915__A1 _17156_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22711__A2 _22708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14530_ _11781_/A _14522_/X _14530_/C VGND VGND VPWR VPWR _14546_/B sky130_fd_sc_hd__and3_4
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23728_ _23728_/CLK _21668_/X VGND VGND VPWR VPWR _16445_/B sky130_fd_sc_hd__dfxtp_4
X_11742_ _16056_/A VGND VGND VPWR VPWR _11742_/X sky130_fd_sc_hd__buf_2
XFILLER_109_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _12428_/A _14459_/X _14460_/X VGND VGND VPWR VPWR _14461_/X sky130_fd_sc_hd__and3_4
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23659_ _23558_/CLK _21775_/X VGND VGND VPWR VPWR _12672_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A VGND VGND VPWR VPWR _11674_/A sky130_fd_sc_hd__buf_2
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _16231_/A _24013_/Q VGND VGND VPWR VPWR _16201_/C sky130_fd_sc_hd__or2_4
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13379_/A _23654_/Q VGND VGND VPWR VPWR _13412_/X sky130_fd_sc_hd__or2_4
XFILLER_128_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17180_ _17137_/X _17168_/X _17112_/X _17179_/X VGND VGND VPWR VPWR _17180_/X sky130_fd_sc_hd__o22a_4
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22475__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14392_ _14511_/A _14392_/B VGND VGND VPWR VPWR _14392_/X sky130_fd_sc_hd__or2_4
XANTENNA__23268__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16131_ _11867_/X _16104_/X _16111_/X _16120_/X _16130_/X VGND VGND VPWR VPWR _16131_/X
+ sky130_fd_sc_hd__a32o_4
X_13343_ _13343_/A VGND VGND VPWR VPWR _13376_/A sky130_fd_sc_hd__buf_2
XANTENNA__17975__A _17974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22592__A2_N _22591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16062_ _16062_/A _15989_/B VGND VGND VPWR VPWR _16063_/C sky130_fd_sc_hd__or2_4
XFILLER_155_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13274_ _12561_/A _13274_/B VGND VGND VPWR VPWR _13274_/X sky130_fd_sc_hd__or2_4
XANTENNA__17694__B _17493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15013_ _11930_/A _15009_/X _15013_/C VGND VGND VPWR VPWR _15014_/B sky130_fd_sc_hd__or3_4
X_12225_ _11935_/A _12225_/B _12224_/X VGND VGND VPWR VPWR _12225_/X sky130_fd_sc_hd__or3_4
XANTENNA__12912__A _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19821_ _19820_/X VGND VGND VPWR VPWR _19821_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21450__A2 _21448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12156_ _12156_/A _23859_/Q VGND VGND VPWR VPWR _12156_/X sky130_fd_sc_hd__or2_4
XFILLER_116_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24139__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12631__B _12500_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_46_0_HCLK clkbuf_6_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19752_ _19749_/X _19752_/B _19883_/A _19752_/D VGND VGND VPWR VPWR _19752_/X sky130_fd_sc_hd__or4_4
X_16964_ _17718_/A VGND VGND VPWR VPWR _16964_/Y sky130_fd_sc_hd__inv_2
X_12087_ _12059_/X _23859_/Q VGND VGND VPWR VPWR _12087_/X sky130_fd_sc_hd__or2_4
XFILLER_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18703_ _18628_/X _17321_/X _18702_/Y VGND VGND VPWR VPWR _18703_/X sky130_fd_sc_hd__o21a_4
X_15915_ _15849_/X VGND VGND VPWR VPWR _15915_/Y sky130_fd_sc_hd__inv_2
X_19683_ _19683_/A _19683_/B VGND VGND VPWR VPWR _19683_/X sky130_fd_sc_hd__or2_4
XFILLER_76_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16895_ _16888_/X _16890_/X _16895_/C _16895_/D VGND VGND VPWR VPWR _16896_/D sky130_fd_sc_hd__and4_4
XANTENNA__13691__A2 _11629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14839__A _14647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18634_ _17109_/X _18599_/B _18538_/X _18601_/Y VGND VGND VPWR VPWR _18634_/X sky130_fd_sc_hd__o22a_4
XFILLER_92_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15846_ _12911_/A _15842_/X _15846_/C VGND VGND VPWR VPWR _15846_/X sky130_fd_sc_hd__or3_4
XANTENNA__21960__A _21960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18565_ _18565_/A _17612_/Y VGND VGND VPWR VPWR _18565_/X sky130_fd_sc_hd__and2_4
XFILLER_64_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12989_ _12854_/A _23528_/Q VGND VGND VPWR VPWR _12990_/C sky130_fd_sc_hd__or2_4
X_15777_ _15770_/A _15704_/B VGND VGND VPWR VPWR _15779_/B sky130_fd_sc_hd__or2_4
XFILLER_75_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22702__A2 _22701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_HCLK clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17516_ _18282_/B _17515_/X VGND VGND VPWR VPWR _17517_/A sky130_fd_sc_hd__or2_4
X_14728_ _13607_/A _14728_/B VGND VGND VPWR VPWR _14729_/C sky130_fd_sc_hd__or2_4
X_18496_ _17717_/X _17764_/X _17717_/X _17764_/X VGND VGND VPWR VPWR _18496_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17447_ _17396_/B _17445_/Y _17446_/X VGND VGND VPWR VPWR _17447_/X sky130_fd_sc_hd__o21a_4
X_14659_ _14680_/A _14659_/B _14659_/C VGND VGND VPWR VPWR _14660_/C sky130_fd_sc_hd__and3_4
XANTENNA__14574__A _14574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17378_ _17378_/A VGND VGND VPWR VPWR _17378_/X sky130_fd_sc_hd__buf_2
XANTENNA__24193__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19117_ _18987_/A _19115_/X _19116_/Y _19106_/X VGND VGND VPWR VPWR _19117_/X sky130_fd_sc_hd__o22a_4
X_16329_ _16316_/A _16270_/B VGND VGND VPWR VPWR _16331_/B sky130_fd_sc_hd__or2_4
XANTENNA__17885__A _18562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17893__A1 _16943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22218__B2 _22212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19048_ _24388_/Q VGND VGND VPWR VPWR _19048_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12822__A _13556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21010_ _19791_/Y _20873_/X _22737_/A _20697_/X VGND VGND VPWR VPWR _21010_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22961_ _22961_/A _22961_/B VGND VGND VPWR VPWR _22963_/B sky130_fd_sc_hd__nand2_4
XANTENNA__22031__A _21991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14749__A _14331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21912_ _21843_/X _21909_/X _23591_/Q _21906_/X VGND VGND VPWR VPWR _21912_/X sky130_fd_sc_hd__o22a_4
XFILLER_56_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22892_ _22876_/X _22832_/X _17353_/Y _22877_/X VGND VGND VPWR VPWR _22892_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21843_ _20596_/A VGND VGND VPWR VPWR _21843_/X sky130_fd_sc_hd__buf_2
XFILLER_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19340__A _19340_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21774_ _21774_/A VGND VGND VPWR VPWR _21774_/X sky130_fd_sc_hd__buf_2
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20486__A _20486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19570__A1 _19469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21139__A2_N _21138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23513_ _23391_/CLK _23513_/D VGND VGND VPWR VPWR _23513_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23410__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20725_ _20257_/X VGND VGND VPWR VPWR _20930_/A sky130_fd_sc_hd__buf_2
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24493_ _24306_/CLK _24493_/D HRESETn VGND VGND VPWR VPWR _20012_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14484__A _12372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11901__A _12854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23444_ _23476_/CLK _22178_/X VGND VGND VPWR VPWR _11828_/B sky130_fd_sc_hd__dfxtp_4
X_20656_ _20857_/A _20655_/X VGND VGND VPWR VPWR _20656_/Y sky130_fd_sc_hd__nand2_4
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19322__A1 _23086_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20468__B1 _20306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23375_ _23760_/CLK _22286_/X VGND VGND VPWR VPWR _16251_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_164_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20587_ _20539_/X _20586_/X _19148_/A _20549_/X VGND VGND VPWR VPWR _20587_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22326_ _22326_/A VGND VGND VPWR VPWR _22326_/X sky130_fd_sc_hd__buf_2
XANTENNA__17884__A1 _17875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21680__A2 _21677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22209__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13828__A _11932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22257_ _22144_/X _22251_/X _14062_/B _22255_/X VGND VGND VPWR VPWR _22257_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12732__A _12298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12010_ _11939_/X _12010_/B _12010_/C VGND VGND VPWR VPWR _12010_/X sky130_fd_sc_hd__or3_4
X_21208_ _20596_/X _21205_/X _23975_/Q _21202_/X VGND VGND VPWR VPWR _23975_/D sky130_fd_sc_hd__o22a_4
XFILLER_133_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21432__A2 _21427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22188_ _22110_/X _22187_/X _23438_/Q _22184_/X VGND VGND VPWR VPWR _22188_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21139_ _21132_/Y _21138_/X _20299_/X _21138_/X VGND VGND VPWR VPWR _24020_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23037__A _22912_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13961_ _13957_/A _23776_/Q VGND VGND VPWR VPWR _13962_/C sky130_fd_sc_hd__or2_4
XFILLER_101_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21196__B2 _21195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13563__A _13563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12912_ _12912_/A _12911_/X VGND VGND VPWR VPWR _12912_/X sky130_fd_sc_hd__and2_4
X_15700_ _13338_/A _15700_/B _15699_/X VGND VGND VPWR VPWR _15700_/X sky130_fd_sc_hd__or3_4
X_16680_ _16677_/A _23666_/Q VGND VGND VPWR VPWR _16681_/C sky130_fd_sc_hd__or2_4
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13892_ _14385_/A _13889_/X _13891_/X VGND VGND VPWR VPWR _13893_/C sky130_fd_sc_hd__and3_4
XANTENNA__20099__C _20098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15631_ _13886_/A _15629_/X _15631_/C VGND VGND VPWR VPWR _15632_/C sky130_fd_sc_hd__and3_4
X_12843_ _12753_/Y _12842_/X VGND VGND VPWR VPWR _12846_/A sky130_fd_sc_hd__and2_4
XANTENNA__12179__A _11671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18350_ _18333_/X _18338_/Y _18344_/X _18348_/X _18349_/Y VGND VGND VPWR VPWR _18350_/X
+ sky130_fd_sc_hd__a32o_4
X_15562_ _14420_/A _15562_/B VGND VGND VPWR VPWR _15562_/X sky130_fd_sc_hd__or2_4
X_12774_ _12759_/A _12774_/B VGND VGND VPWR VPWR _12774_/X sky130_fd_sc_hd__or2_4
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20396__A _20396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22696__B2 _22691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14513_/A _14513_/B _14513_/C VGND VGND VPWR VPWR _14514_/C sky130_fd_sc_hd__or3_4
X_17301_ _17301_/A _17300_/X VGND VGND VPWR VPWR _17301_/Y sky130_fd_sc_hd__nand2_4
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _13256_/A VGND VGND VPWR VPWR _12370_/A sky130_fd_sc_hd__buf_2
X_15493_ _13753_/A _15493_/B VGND VGND VPWR VPWR _15493_/X sky130_fd_sc_hd__or2_4
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18281_ _18407_/A _17515_/X VGND VGND VPWR VPWR _18281_/Y sky130_fd_sc_hd__nor2_4
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20171__A2 IRQ[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _15393_/A _14500_/B VGND VGND VPWR VPWR _14445_/C sky130_fd_sc_hd__or2_4
X_17232_ _17130_/X VGND VGND VPWR VPWR _17233_/A sky130_fd_sc_hd__buf_2
XANTENNA__22448__B2 _22445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _13923_/A VGND VGND VPWR VPWR _12410_/A sky130_fd_sc_hd__buf_2
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20459__B1 _20714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17163_ _17162_/Y _17144_/X _12982_/X _17146_/X VGND VGND VPWR VPWR _17163_/X sky130_fd_sc_hd__o22a_4
X_14375_ _14375_/A VGND VGND VPWR VPWR _14540_/A sky130_fd_sc_hd__buf_2
XFILLER_35_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _11513_/Y _11544_/X _24407_/Q _11586_/X VGND VGND VPWR VPWR _11587_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21120__B2 _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16114_ _16101_/A VGND VGND VPWR VPWR _16147_/A sky130_fd_sc_hd__buf_2
X_13326_ _13320_/A _24102_/Q VGND VGND VPWR VPWR _13326_/X sky130_fd_sc_hd__or2_4
XANTENNA__21671__A2 _21670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17094_ _18008_/A VGND VGND VPWR VPWR _17094_/Y sky130_fd_sc_hd__inv_2
X_16045_ _16057_/A _23694_/Q VGND VGND VPWR VPWR _16047_/B sky130_fd_sc_hd__or2_4
XFILLER_142_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13257_ _13235_/A _13255_/X _13257_/C VGND VGND VPWR VPWR _13258_/C sky130_fd_sc_hd__and3_4
XANTENNA__12642__A _12587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12208_ _12571_/A _12208_/B _12207_/X VGND VGND VPWR VPWR _12208_/X sky130_fd_sc_hd__or3_4
XFILLER_9_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13188_ _12851_/A _13188_/B _13187_/X VGND VGND VPWR VPWR _13189_/C sky130_fd_sc_hd__and3_4
XANTENNA__22620__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19804_ _19516_/X _19793_/X _19803_/X VGND VGND VPWR VPWR _19804_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15953__A _13330_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12139_ _12127_/A _23699_/Q VGND VGND VPWR VPWR _12141_/B sky130_fd_sc_hd__or2_4
XANTENNA__19425__A _19428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17996_ _17996_/A VGND VGND VPWR VPWR _17996_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19735_ _20512_/B _19573_/X _19734_/X _19638_/X VGND VGND VPWR VPWR _19735_/X sky130_fd_sc_hd__a211o_4
X_16947_ _24159_/Q VGND VGND VPWR VPWR _16997_/A sky130_fd_sc_hd__inv_2
XFILLER_84_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14569__A _14448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13473__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19666_ _19662_/X _19828_/C _19546_/A VGND VGND VPWR VPWR _19666_/Y sky130_fd_sc_hd__o21ai_4
X_16878_ _16878_/A _16874_/Y _16876_/X _16877_/X VGND VGND VPWR VPWR _16878_/X sky130_fd_sc_hd__and4_4
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23433__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18617_ _24138_/Q _22935_/B _16976_/X VGND VGND VPWR VPWR _22943_/B sky130_fd_sc_hd__o21a_4
XANTENNA__16602__A2 _11632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15829_ _12891_/A _15829_/B VGND VGND VPWR VPWR _15829_/X sky130_fd_sc_hd__or2_4
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19597_ _19589_/X _19724_/A _19596_/X VGND VGND VPWR VPWR _19597_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14613__A1 _11854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14613__B2 _14612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18548_ _18506_/A _18540_/Y _18541_/X _18543_/X _18547_/Y VGND VGND VPWR VPWR _18548_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18479_ _16980_/X VGND VGND VPWR VPWR _18479_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22439__A1 _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20510_ _20510_/A VGND VGND VPWR VPWR _20510_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21490_ _21263_/X _21485_/X _12565_/B _21489_/X VGND VGND VPWR VPWR _21490_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22439__B2 _22433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20441_ _20441_/A VGND VGND VPWR VPWR _20441_/X sky130_fd_sc_hd__buf_2
XFILLER_14_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18504__A _18032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23160_ _23194_/CLK _23160_/D VGND VGND VPWR VPWR _23160_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_134_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20372_ _17957_/X _20260_/X _20341_/X _20371_/Y VGND VGND VPWR VPWR _20372_/X sky130_fd_sc_hd__a211o_4
XFILLER_173_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14751__B _14751_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22111_ _22123_/A VGND VGND VPWR VPWR _22111_/X sky130_fd_sc_hd__buf_2
XFILLER_134_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20870__B1 HRDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13648__A _11878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23091_ _16901_/A VGND VGND VPWR VPWR HSIZE[0] sky130_fd_sc_hd__buf_2
XFILLER_133_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24373__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22042_ _22057_/A VGND VGND VPWR VPWR _22042_/X sky130_fd_sc_hd__buf_2
XANTENNA__21865__A _20819_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21414__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22611__B2 _22605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15863__A _15887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19335__A _20200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23993_ _24057_/CLK _23993_/D VGND VGND VPWR VPWR _14721_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14479__A _14292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21178__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13383__A _13383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22944_ _18613_/X _22930_/Y _19319_/X _22943_/X VGND VGND VPWR VPWR _22945_/C sky130_fd_sc_hd__a211o_4
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22875_ _19909_/X VGND VGND VPWR VPWR _22875_/X sky130_fd_sc_hd__buf_2
XFILLER_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21826_ _20441_/A VGND VGND VPWR VPWR _21826_/X sky130_fd_sc_hd__buf_2
XANTENNA__22678__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21757_ _21756_/X VGND VGND VPWR VPWR _21791_/A sky130_fd_sc_hd__buf_2
XANTENNA__12727__A _12727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21350__B2 _21345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15103__A _15103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20708_ _20325_/X VGND VGND VPWR VPWR _20708_/X sky130_fd_sc_hd__buf_2
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _12890_/A _12465_/X _12490_/C VGND VGND VPWR VPWR _12490_/X sky130_fd_sc_hd__or3_4
X_24476_ _23126_/CLK _18621_/X HRESETn VGND VGND VPWR VPWR _24476_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21688_ _21674_/A VGND VGND VPWR VPWR _21688_/X sky130_fd_sc_hd__buf_2
XANTENNA__20944__A HRDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23427_ _23523_/CLK _22203_/X VGND VGND VPWR VPWR _15830_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20639_ _20639_/A VGND VGND VPWR VPWR _20639_/X sky130_fd_sc_hd__buf_2
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24484__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21102__B2 _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14160_ _14988_/A VGND VGND VPWR VPWR _14267_/A sky130_fd_sc_hd__buf_2
XANTENNA__22850__A1 _15048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21653__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23358_ _23518_/CLK _22310_/X VGND VGND VPWR VPWR _13605_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13111_ _13103_/A _13109_/X _13111_/C VGND VGND VPWR VPWR _13115_/B sky130_fd_sc_hd__and3_4
XANTENNA__13558__A _13546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22309_ _22146_/X _22308_/X _23359_/Q _22305_/X VGND VGND VPWR VPWR _23359_/D sky130_fd_sc_hd__o22a_4
XFILLER_153_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14091_ _14138_/A _23519_/Q VGND VGND VPWR VPWR _14092_/C sky130_fd_sc_hd__or2_4
Xclkbuf_7_111_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR _23557_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12462__A _12881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23289_ _23290_/CLK _22399_/X VGND VGND VPWR VPWR _14717_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13042_ _13042_/A _23720_/Q VGND VGND VPWR VPWR _13044_/B sky130_fd_sc_hd__or2_4
XFILLER_4_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22602__B2 _22598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15773__A _11689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17850_ _17823_/A VGND VGND VPWR VPWR _17850_/X sky130_fd_sc_hd__buf_2
XFILLER_26_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16801_ _16606_/A _16801_/B _16800_/X VGND VGND VPWR VPWR _16801_/X sky130_fd_sc_hd__or3_4
XANTENNA__23456__CLK _23456_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17781_ _17657_/Y _17779_/X _17959_/A VGND VGND VPWR VPWR _17781_/X sky130_fd_sc_hd__a21bo_4
XFILLER_94_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14993_ _14155_/A VGND VGND VPWR VPWR _14994_/A sky130_fd_sc_hd__buf_2
XANTENNA__13293__A _13304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11806__A _16647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19520_ _20672_/A _19518_/X _19519_/X HRDATA[14] VGND VGND VPWR VPWR _19520_/Y sky130_fd_sc_hd__a22oi_4
X_16732_ _16732_/A _16730_/X _16731_/X VGND VGND VPWR VPWR _16733_/C sky130_fd_sc_hd__and3_4
X_13944_ _11813_/A _13944_/B _13943_/X VGND VGND VPWR VPWR _13945_/C sky130_fd_sc_hd__or3_4
XFILLER_75_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20916__A1 _20894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20916__B2 _20861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19451_ _19767_/A VGND VGND VPWR VPWR _19507_/A sky130_fd_sc_hd__inv_2
X_16663_ _16646_/A _16661_/X _16663_/C VGND VGND VPWR VPWR _16667_/B sky130_fd_sc_hd__and3_4
X_13875_ _13888_/A VGND VGND VPWR VPWR _14386_/A sky130_fd_sc_hd__buf_2
X_18402_ _18402_/A _18368_/X VGND VGND VPWR VPWR _18402_/X sky130_fd_sc_hd__and2_4
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12826_ _13343_/A _12824_/X _12826_/C VGND VGND VPWR VPWR _12826_/X sky130_fd_sc_hd__and3_4
X_15614_ _13885_/A _15540_/B VGND VGND VPWR VPWR _15615_/C sky130_fd_sc_hd__or2_4
X_19382_ _19377_/X _18776_/Y _19381_/X _24245_/Q VGND VGND VPWR VPWR _19382_/X sky130_fd_sc_hd__a2bb2o_4
X_16594_ _16594_/A _23826_/Q VGND VGND VPWR VPWR _16594_/X sky130_fd_sc_hd__or2_4
XFILLER_163_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18333_ _18405_/A _17508_/X VGND VGND VPWR VPWR _18333_/X sky130_fd_sc_hd__or2_4
X_12757_ _13067_/A VGND VGND VPWR VPWR _12758_/A sky130_fd_sc_hd__buf_2
X_15545_ _13687_/A _15543_/X _15544_/X VGND VGND VPWR VPWR _15545_/X sky130_fd_sc_hd__and3_4
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11708_ _11708_/A VGND VGND VPWR VPWR _13866_/A sky130_fd_sc_hd__buf_2
XANTENNA__15013__A _11930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15476_ _13063_/A _15472_/X _15475_/X VGND VGND VPWR VPWR _15476_/X sky130_fd_sc_hd__or3_4
X_18264_ _18264_/A VGND VGND VPWR VPWR _18264_/Y sky130_fd_sc_hd__inv_2
X_12688_ _11881_/A _12688_/B _12687_/X VGND VGND VPWR VPWR _12692_/B sky130_fd_sc_hd__and3_4
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ _14431_/A _14427_/B _14426_/X VGND VGND VPWR VPWR _14427_/X sky130_fd_sc_hd__and3_4
X_17215_ _16242_/X _17115_/X _14413_/Y _17116_/X VGND VGND VPWR VPWR _17215_/X sky130_fd_sc_hd__o22a_4
X_11639_ _11639_/A VGND VGND VPWR VPWR _11640_/B sky130_fd_sc_hd__inv_2
X_18195_ _18378_/A _17486_/Y VGND VGND VPWR VPWR _18196_/D sky130_fd_sc_hd__and2_4
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21644__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22841__A1 _15915_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17146_ _17146_/A VGND VGND VPWR VPWR _17146_/X sky130_fd_sc_hd__buf_2
X_14358_ _11681_/A _14347_/X _14357_/X VGND VGND VPWR VPWR _14358_/X sky130_fd_sc_hd__and3_4
XFILLER_171_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13468__A _13468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13309_ _13309_/A _13309_/B VGND VGND VPWR VPWR _13311_/B sky130_fd_sc_hd__or2_4
XFILLER_143_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17077_ _17077_/A VGND VGND VPWR VPWR _17077_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12372__A _12372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14289_ _15402_/A _22346_/A VGND VGND VPWR VPWR _14289_/X sky130_fd_sc_hd__or2_4
XFILLER_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24231__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16028_ _16062_/A _23790_/Q VGND VGND VPWR VPWR _16029_/C sky130_fd_sc_hd__or2_4
XFILLER_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19470__B1 _18027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18273__B2 _18272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_16_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__16823__A2 _16821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17979_ _17976_/X _17978_/X _17882_/X VGND VGND VPWR VPWR _17979_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__14299__A _13823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19718_ _19705_/X _19787_/A _19603_/X _19717_/Y VGND VGND VPWR VPWR _19718_/X sky130_fd_sc_hd__a211o_4
X_20990_ _20990_/A VGND VGND VPWR VPWR _20990_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19649_ _19649_/A _19649_/B VGND VGND VPWR VPWR _19657_/C sky130_fd_sc_hd__nor2_4
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17403__A _13945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13931__A _14385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22660_ _22440_/X _22658_/X _13025_/B _22655_/X VGND VGND VPWR VPWR _22660_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14746__B _23385_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21611_ _21602_/Y _21610_/X _21526_/X _21610_/X VGND VGND VPWR VPWR _21611_/X sky130_fd_sc_hd__a2bb2o_4
X_22591_ _22598_/A VGND VGND VPWR VPWR _22591_/X sky130_fd_sc_hd__buf_2
XANTENNA__12547__A _12911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16019__A _16047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21332__B2 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24330_ _24342_/CLK _19182_/X HRESETn VGND VGND VPWR VPWR _19151_/A sky130_fd_sc_hd__dfrtp_4
X_21542_ _21542_/A VGND VGND VPWR VPWR _21542_/X sky130_fd_sc_hd__buf_2
XFILLER_21_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15858__A _15851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24261_ _24127_/CLK _24261_/D HRESETn VGND VGND VPWR VPWR _24261_/Q sky130_fd_sc_hd__dfrtp_4
X_21473_ _21506_/A VGND VGND VPWR VPWR _21489_/A sky130_fd_sc_hd__inv_2
XANTENNA__11601__D _18782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23212_ _23728_/CLK _23212_/D VGND VGND VPWR VPWR _12344_/B sky130_fd_sc_hd__dfxtp_4
X_20424_ _20490_/A VGND VGND VPWR VPWR _20425_/A sky130_fd_sc_hd__buf_2
XFILLER_162_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21635__A2 _21634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24192_ _24182_/CLK _19838_/X HRESETn VGND VGND VPWR VPWR _16901_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13378__A _13378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23143_ _24039_/CLK _23143_/D VGND VGND VPWR VPWR _13237_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_49_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20355_ _17892_/X _20260_/X _20341_/X _20354_/Y VGND VGND VPWR VPWR _20355_/X sky130_fd_sc_hd__a211o_4
XFILLER_84_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18888__B _18888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23074_ _17650_/X _23079_/B VGND VGND VPWR VPWR _23074_/X sky130_fd_sc_hd__or2_4
XANTENNA__23479__CLK _23864_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20286_ _20264_/X VGND VGND VPWR VPWR _20287_/A sky130_fd_sc_hd__inv_2
XFILLER_103_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21399__B2 _21395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17067__A2 _11595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22025_ _21862_/X _22024_/X _23519_/Q _22021_/X VGND VGND VPWR VPWR _22025_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15593__A _15620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22899__A1 _12112_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23976_ _24073_/CLK _21207_/X VGND VGND VPWR VPWR _23976_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_152_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11990_ _11990_/A _24084_/Q VGND VGND VPWR VPWR _11990_/X sky130_fd_sc_hd__or2_4
XFILLER_60_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22927_ _22908_/X _18627_/X _22909_/X _22926_/X VGND VGND VPWR VPWR _22927_/X sky130_fd_sc_hd__a211o_4
XFILLER_17_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20374__A2 _20365_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21571__B2 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13841__A _13658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13660_ _11879_/A _13658_/X _13659_/X VGND VGND VPWR VPWR _13661_/C sky130_fd_sc_hd__and3_4
X_22858_ _17518_/Y _22847_/X _22853_/X _22857_/X VGND VGND VPWR VPWR _22859_/A sky130_fd_sc_hd__a211o_4
XFILLER_71_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_36_0_HCLK clkbuf_7_37_0_HCLK/A VGND VGND VPWR VPWR _23889_/CLK sky130_fd_sc_hd__clkbuf_1
X_12611_ _12632_/A _12611_/B VGND VGND VPWR VPWR _12611_/X sky130_fd_sc_hd__or2_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21809_ _21834_/A VGND VGND VPWR VPWR _21809_/X sky130_fd_sc_hd__buf_2
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13591_ _13591_/A VGND VGND VPWR VPWR _13965_/A sky130_fd_sc_hd__buf_2
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_99_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR _23908_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_12_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22789_ _22766_/Y _22788_/B VGND VGND VPWR VPWR _22789_/Y sky130_fd_sc_hd__nand2_4
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15330_ _15330_/A _15324_/X _15329_/X VGND VGND VPWR VPWR _15331_/C sky130_fd_sc_hd__or3_4
X_12542_ _12895_/A _12647_/B VGND VGND VPWR VPWR _12543_/C sky130_fd_sc_hd__or2_4
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23050__A _18101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15261_ _15257_/A _23768_/Q VGND VGND VPWR VPWR _15262_/C sky130_fd_sc_hd__or2_4
XANTENNA__23076__A1 _19953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12473_ _12473_/A VGND VGND VPWR VPWR _12474_/A sky130_fd_sc_hd__buf_2
X_24459_ _23347_/CLK _18802_/X HRESETn VGND VGND VPWR VPWR _11554_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16750__A1 _12027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17000_ _16999_/X VGND VGND VPWR VPWR _17000_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24254__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14212_ _14635_/A _14209_/X _14212_/C VGND VGND VPWR VPWR _14212_/X sky130_fd_sc_hd__and3_4
XFILLER_172_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21626__A2 _21620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15487__B _15487_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15192_ _14769_/A _15188_/X _15192_/C VGND VGND VPWR VPWR _15202_/B sky130_fd_sc_hd__or3_4
XANTENNA__14391__B _14391_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_HCLK clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_3_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13288__A _13318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14143_ _12287_/A _14143_/B _14142_/X VGND VGND VPWR VPWR _14143_/X sky130_fd_sc_hd__or3_4
XANTENNA__12192__A _13042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18951_ _24404_/Q _18953_/B _18950_/A _11544_/C _18950_/Y VGND VGND VPWR VPWR _24372_/D
+ sky130_fd_sc_hd__a32o_4
X_14074_ _14074_/A _14069_/X _14073_/X VGND VGND VPWR VPWR _14074_/X sky130_fd_sc_hd__or3_4
XANTENNA__16599__A _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13025_ _12905_/A _13025_/B VGND VGND VPWR VPWR _13027_/B sky130_fd_sc_hd__or2_4
XFILLER_106_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17902_ _16997_/B VGND VGND VPWR VPWR _17902_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12920__A _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22051__A2 _22046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18882_ _15380_/A _18877_/X _24408_/Q _18878_/X VGND VGND VPWR VPWR _18882_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20062__A1 _20040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17833_ _17833_/A VGND VGND VPWR VPWR _17833_/X sky130_fd_sc_hd__buf_2
XFILLER_120_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17764_ _17720_/X _17724_/X _17762_/X _17720_/B _17763_/Y VGND VGND VPWR VPWR _17764_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_66_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14976_ _14976_/A _23222_/Q VGND VGND VPWR VPWR _14976_/X sky130_fd_sc_hd__or2_4
XANTENNA__21011__B1 _20262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19503_ _19546_/A _19537_/B VGND VGND VPWR VPWR _19503_/X sky130_fd_sc_hd__and2_4
XFILLER_35_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16715_ _11941_/A _16776_/B VGND VGND VPWR VPWR _16715_/X sky130_fd_sc_hd__or2_4
X_13927_ _14335_/A _13927_/B _13927_/C VGND VGND VPWR VPWR _13927_/X sky130_fd_sc_hd__or3_4
X_17695_ _16986_/A _17501_/X VGND VGND VPWR VPWR _17772_/A sky130_fd_sc_hd__and2_4
XFILLER_63_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21562__B2 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19434_ _19433_/X _18727_/X _19433_/X _24214_/Q VGND VGND VPWR VPWR _19434_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16646_ _16646_/A _16644_/X _16645_/X VGND VGND VPWR VPWR _16646_/X sky130_fd_sc_hd__and3_4
XFILLER_62_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13858_ _15447_/A _13933_/B VGND VGND VPWR VPWR _13859_/C sky130_fd_sc_hd__or2_4
XFILLER_16_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12809_ _12759_/A _12809_/B VGND VGND VPWR VPWR _12809_/X sky130_fd_sc_hd__or2_4
XFILLER_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19365_ _19372_/A VGND VGND VPWR VPWR _19365_/X sky130_fd_sc_hd__buf_2
XANTENNA__12367__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16577_ _16592_/A _16577_/B _16577_/C VGND VGND VPWR VPWR _16577_/X sky130_fd_sc_hd__or3_4
XANTENNA__21314__B2 _21239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13789_ _13591_/A VGND VGND VPWR VPWR _13954_/A sky130_fd_sc_hd__buf_2
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18316_ _17856_/X _18046_/Y _17985_/X _18048_/X VGND VGND VPWR VPWR _18316_/X sky130_fd_sc_hd__o22a_4
X_15528_ _12186_/A _15524_/X _15528_/C VGND VGND VPWR VPWR _15528_/X sky130_fd_sc_hd__or3_4
X_19296_ _24289_/Q _19237_/X _19295_/Y VGND VGND VPWR VPWR _19296_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24335__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20584__A _20270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18247_ _16985_/X VGND VGND VPWR VPWR _18248_/C sky130_fd_sc_hd__inv_2
X_15459_ _12592_/A _23746_/Q VGND VGND VPWR VPWR _15460_/C sky130_fd_sc_hd__or2_4
XANTENNA__21078__B1 _14884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18178_ _18150_/X _18156_/Y _18163_/X _18175_/X _18177_/Y VGND VGND VPWR VPWR _18178_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13198__A _13052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17129_ _12097_/X VGND VGND VPWR VPWR _17160_/A sky130_fd_sc_hd__buf_2
XANTENNA__22290__A2 _22287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20140_ _11555_/X VGND VGND VPWR VPWR _20140_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13926__A _13720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20071_ _20071_/A VGND VGND VPWR VPWR _20071_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20589__C1 _20588_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23771__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20053__A1 _20040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23830_ _23862_/CLK _23830_/D VGND VGND VPWR VPWR _14959_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_100_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24127__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23761_ _23761_/CLK _23761_/D VGND VGND VPWR VPWR _23761_/Q sky130_fd_sc_hd__dfxtp_4
X_20973_ _21017_/A _20973_/B VGND VGND VPWR VPWR _20973_/Y sky130_fd_sc_hd__nor2_4
XPHY_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22712_ _22705_/A VGND VGND VPWR VPWR _22712_/X sky130_fd_sc_hd__buf_2
XANTENNA__13661__A _11933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23692_ _24012_/CLK _21723_/X VGND VGND VPWR VPWR _23692_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22643_ _22672_/A VGND VGND VPWR VPWR _22658_/A sky130_fd_sc_hd__buf_2
XANTENNA__12277__A _12273_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21856__A2 _21851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22574_ _22464_/X _22572_/X _13721_/B _22569_/X VGND VGND VPWR VPWR _22574_/X sky130_fd_sc_hd__o22a_4
XFILLER_142_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24313_ _24292_/CLK _19216_/X HRESETn VGND VGND VPWR VPWR _19134_/A sky130_fd_sc_hd__dfrtp_4
X_21525_ _21524_/X VGND VGND VPWR VPWR _21525_/X sky130_fd_sc_hd__buf_2
XANTENNA__15588__A _15606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24244_ _24471_/CLK _19387_/X HRESETn VGND VGND VPWR VPWR _24244_/Q sky130_fd_sc_hd__dfrtp_4
X_21456_ _21292_/X _21455_/X _23839_/Q _21452_/X VGND VGND VPWR VPWR _23839_/D sky130_fd_sc_hd__o22a_4
XFILLER_5_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20407_ _20754_/A _20406_/X _19156_/A _20761_/A VGND VGND VPWR VPWR _20407_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24175_ _24184_/CLK _24175_/D HRESETn VGND VGND VPWR VPWR _24175_/Q sky130_fd_sc_hd__dfrtp_4
X_21387_ _21261_/X _21384_/X _12314_/B _21381_/X VGND VGND VPWR VPWR _21387_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22281__A2 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23126_ _23126_/CLK _22684_/X VGND VGND VPWR VPWR _14958_/B sky130_fd_sc_hd__dfxtp_4
X_20338_ _20302_/X _20337_/X _24115_/Q _20225_/X VGND VGND VPWR VPWR _24115_/D sky130_fd_sc_hd__o22a_4
XFILLER_107_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23057_ _23036_/X _17660_/A _23048_/X _23056_/X VGND VGND VPWR VPWR _23058_/A sky130_fd_sc_hd__a211o_4
XANTENNA__17308__A _14412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22033__A2 _22031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20269_ _20269_/A VGND VGND VPWR VPWR _20269_/X sky130_fd_sc_hd__buf_2
XANTENNA__20044__A1 _20040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22008_ _21833_/X _22003_/X _12584_/B _22007_/X VGND VGND VPWR VPWR _23531_/D sky130_fd_sc_hd__o22a_4
XFILLER_76_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21792__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14830_ _14691_/A _14760_/B VGND VGND VPWR VPWR _14832_/B sky130_fd_sc_hd__or2_4
XANTENNA__20669__A HRDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11973_ _16130_/A VGND VGND VPWR VPWR _11973_/X sky130_fd_sc_hd__buf_2
X_14761_ _13637_/A _14761_/B VGND VGND VPWR VPWR _14761_/X sky130_fd_sc_hd__or2_4
XFILLER_5_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23959_ _23416_/CLK _23959_/D VGND VGND VPWR VPWR _15156_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_44_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16500_ _16479_/X _16431_/B VGND VGND VPWR VPWR _16500_/X sky130_fd_sc_hd__or2_4
XFILLER_72_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13571__A _13342_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16015__A3 _15980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13712_ _12600_/A VGND VGND VPWR VPWR _15487_/A sky130_fd_sc_hd__buf_2
XFILLER_45_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14692_ _14679_/A _14598_/B VGND VGND VPWR VPWR _14692_/X sky130_fd_sc_hd__or2_4
X_17480_ _12574_/X VGND VGND VPWR VPWR _17480_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22884__A _22884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16431_ _16402_/X _16431_/B VGND VGND VPWR VPWR _16431_/X sky130_fd_sc_hd__or2_4
XFILLER_60_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13643_ _13652_/A _13732_/B VGND VGND VPWR VPWR _13643_/X sky130_fd_sc_hd__or2_4
XANTENNA__12187__A _13045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19150_ _24329_/Q _19185_/A VGND VGND VPWR VPWR _19151_/B sky130_fd_sc_hd__and2_4
XANTENNA__21847__A2 _21839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16362_ _13399_/A VGND VGND VPWR VPWR _16362_/X sky130_fd_sc_hd__buf_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13574_ _13126_/X _13265_/Y _13269_/A _13573_/Y VGND VGND VPWR VPWR _13574_/X sky130_fd_sc_hd__a211o_4
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18101_ _18074_/X _18080_/Y _18093_/X _18099_/X _18100_/Y VGND VGND VPWR VPWR _18101_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _13483_/A _12459_/X _12490_/X _12516_/X _12524_/X VGND VGND VPWR VPWR _12525_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23644__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15313_ _13951_/X _11627_/A _15282_/X _11604_/A _15312_/X VGND VGND VPWR VPWR _15382_/A
+ sky130_fd_sc_hd__a32o_4
X_16293_ _11890_/X _16293_/B VGND VGND VPWR VPWR _16293_/X sky130_fd_sc_hd__or2_4
X_19081_ _19068_/X _19080_/X _19068_/X _19075_/A VGND VGND VPWR VPWR _24351_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12915__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18032_ _16939_/X VGND VGND VPWR VPWR _18032_/X sky130_fd_sc_hd__buf_2
XFILLER_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12456_ _12876_/A VGND VGND VPWR VPWR _12885_/A sky130_fd_sc_hd__buf_2
XFILLER_145_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15244_ _14254_/A _15172_/B VGND VGND VPWR VPWR _15246_/B sky130_fd_sc_hd__or2_4
XFILLER_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15175_ _14301_/A _15175_/B _15175_/C VGND VGND VPWR VPWR _15175_/X sky130_fd_sc_hd__or3_4
X_12387_ _12387_/A _12387_/B _12387_/C VGND VGND VPWR VPWR _12388_/C sky130_fd_sc_hd__and3_4
XFILLER_99_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14126_ _14905_/A VGND VGND VPWR VPWR _14127_/A sky130_fd_sc_hd__buf_2
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19983_ _19961_/X VGND VGND VPWR VPWR _19983_/X sky130_fd_sc_hd__buf_2
XFILLER_158_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18934_ _18896_/A VGND VGND VPWR VPWR _18934_/X sky130_fd_sc_hd__buf_2
XFILLER_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14057_ _11698_/A _14055_/X _14057_/C VGND VGND VPWR VPWR _14057_/X sky130_fd_sc_hd__and3_4
XANTENNA__12650__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13008_ _12911_/A _13008_/B _13007_/X VGND VGND VPWR VPWR _13008_/X sky130_fd_sc_hd__or3_4
XANTENNA__19976__A1 _16943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21232__B1 _23957_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18865_ _13567_/X _18863_/X _24421_/Q _18864_/X VGND VGND VPWR VPWR _18865_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21783__B2 _21781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19433__A _19428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17816_ _17233_/A VGND VGND VPWR VPWR _17816_/X sky130_fd_sc_hd__buf_2
X_18796_ _18796_/A VGND VGND VPWR VPWR _18796_/X sky130_fd_sc_hd__buf_2
XANTENNA__14265__A2 _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17747_ _17743_/A _17298_/X _17743_/X VGND VGND VPWR VPWR _17747_/X sky130_fd_sc_hd__a21bo_4
X_14959_ _14919_/A _14959_/B VGND VGND VPWR VPWR _14959_/X sky130_fd_sc_hd__or2_4
XANTENNA__14577__A _13596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13481__A _12515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21535__B2 _21525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17678_ _18190_/A _17464_/X VGND VGND VPWR VPWR _17699_/A sky130_fd_sc_hd__and2_4
X_19417_ _19414_/X _18457_/Y _19414_/X _24226_/Q VGND VGND VPWR VPWR _19417_/X sky130_fd_sc_hd__a2bb2o_4
X_16629_ _16682_/A _16623_/X _16629_/C VGND VGND VPWR VPWR _16629_/X sky130_fd_sc_hd__or3_4
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12097__A _12105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19348_ _19347_/X _18212_/X _19347_/X _24267_/Q VGND VGND VPWR VPWR _19348_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_82_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR _23511_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_149_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19279_ _19247_/B VGND VGND VPWR VPWR _19279_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12825__A _12801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21310_ _21309_/X _21305_/X _23928_/Q _21300_/X VGND VGND VPWR VPWR _23928_/D sky130_fd_sc_hd__o22a_4
X_22290_ _22115_/X _22287_/X _12204_/B _22284_/X VGND VGND VPWR VPWR _22290_/X sky130_fd_sc_hd__o22a_4
X_21241_ _21526_/A VGND VGND VPWR VPWR _21241_/X sky130_fd_sc_hd__buf_2
XANTENNA__22263__A2 _22258_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21172_ _20841_/X _21169_/X _23997_/Q _21166_/X VGND VGND VPWR VPWR _23997_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13656__A _13656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20123_ _20120_/X _20122_/Y _20110_/Y VGND VGND VPWR VPWR _20123_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__22015__A2 _22010_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12560__A _12569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20054_ _20053_/X VGND VGND VPWR VPWR _20054_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20577__A2 _19773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19343__A _19340_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20489__A _20257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23813_ _23557_/CLK _23813_/D VGND VGND VPWR VPWR _13477_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_27_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22723__B1 _23103_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13391__A _13413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _23744_/CLK _23744_/D VGND VGND VPWR VPWR _23744_/Q sky130_fd_sc_hd__dfxtp_4
X_20956_ _20977_/A _20955_/X VGND VGND VPWR VPWR _20956_/Y sky130_fd_sc_hd__nand2_4
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__A1 _11984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23675_/CLK _23675_/D VGND VGND VPWR VPWR _14436_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _20639_/A _20875_/X _20779_/X _20886_/Y VGND VGND VPWR VPWR _20887_/X sky130_fd_sc_hd__a211o_4
XFILLER_41_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22626_ _22605_/A VGND VGND VPWR VPWR _22626_/X sky130_fd_sc_hd__buf_2
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22557_ _22435_/X _22551_/X _12774_/B _22555_/X VGND VGND VPWR VPWR _23210_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12735__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16207__A _13383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12310_ _13152_/A _12398_/B VGND VGND VPWR VPWR _12312_/B sky130_fd_sc_hd__or2_4
XANTENNA__15111__A _15080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21508_ _21295_/X _21506_/X _13766_/B _21503_/X VGND VGND VPWR VPWR _21508_/X sky130_fd_sc_hd__o22a_4
X_13290_ _13290_/A VGND VGND VPWR VPWR _13330_/A sky130_fd_sc_hd__buf_2
X_22488_ _22487_/X VGND VGND VPWR VPWR _22489_/A sky130_fd_sc_hd__buf_2
X_12241_ _13164_/A _12374_/B VGND VGND VPWR VPWR _12241_/X sky130_fd_sc_hd__or2_4
X_24227_ _24127_/CLK _19416_/X HRESETn VGND VGND VPWR VPWR _24227_/Q sky130_fd_sc_hd__dfrtp_4
X_21439_ _21263_/X _21434_/X _12549_/B _21438_/X VGND VGND VPWR VPWR _21439_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22254__A2 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14950__A _11673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24158_ _24158_/CLK _20002_/Y HRESETn VGND VGND VPWR VPWR _16948_/A sky130_fd_sc_hd__dfrtp_4
X_12172_ _12122_/A _12172_/B _12172_/C VGND VGND VPWR VPWR _12172_/X sky130_fd_sc_hd__and3_4
X_23109_ _23557_/CLK _23109_/D VGND VGND VPWR VPWR _13476_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13566__A _13566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22006__A2 _22003_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12470__A _12470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16980_ _16964_/Y _16979_/X VGND VGND VPWR VPWR _16980_/X sky130_fd_sc_hd__or2_4
X_24089_ _24057_/CLK _20939_/X VGND VGND VPWR VPWR _14751_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_122_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15931_ _13272_/X _13585_/X _12987_/X _15931_/D VGND VGND VPWR VPWR _15932_/C sky130_fd_sc_hd__or4_4
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15781__A _13123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21765__B2 _21760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18650_ _17301_/A _18648_/X VGND VGND VPWR VPWR _18650_/X sky130_fd_sc_hd__or2_4
X_15862_ _13521_/X _15862_/B _15861_/X VGND VGND VPWR VPWR _15863_/C sky130_fd_sc_hd__and3_4
XFILLER_114_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17601_ _17495_/X _17504_/A _17508_/B VGND VGND VPWR VPWR _17601_/X sky130_fd_sc_hd__a21o_4
X_14813_ _14820_/A _14737_/B VGND VGND VPWR VPWR _14813_/X sky130_fd_sc_hd__or2_4
X_18581_ _17109_/X _17635_/D _18538_/X _18418_/A VGND VGND VPWR VPWR _18581_/X sky130_fd_sc_hd__o22a_4
X_15793_ _12848_/A _15854_/B VGND VGND VPWR VPWR _15793_/X sky130_fd_sc_hd__or2_4
XFILLER_40_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21517__B2 _21482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11814__A _12978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17532_ _17509_/Y _17530_/Y _17531_/X VGND VGND VPWR VPWR _17532_/X sky130_fd_sc_hd__o21a_4
XFILLER_83_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21007__B _21007_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14744_ _13655_/A _14744_/B VGND VGND VPWR VPWR _14744_/X sky130_fd_sc_hd__or2_4
X_11956_ _12103_/A _24020_/Q VGND VGND VPWR VPWR _11957_/C sky130_fd_sc_hd__or2_4
XFILLER_33_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22190__B2 _22184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17463_ _16702_/A _17481_/B VGND VGND VPWR VPWR _17463_/X sky130_fd_sc_hd__and2_4
X_11887_ _11887_/A VGND VGND VPWR VPWR _11888_/A sky130_fd_sc_hd__buf_2
XFILLER_72_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14675_ _14675_/A _14591_/B VGND VGND VPWR VPWR _14676_/C sky130_fd_sc_hd__or2_4
X_19202_ _19141_/A _19141_/B _19201_/Y VGND VGND VPWR VPWR _19202_/X sky130_fd_sc_hd__o21a_4
X_16414_ _13467_/A _16412_/X _16413_/X VGND VGND VPWR VPWR _16414_/X sky130_fd_sc_hd__and3_4
X_13626_ _15405_/A _13620_/X _13626_/C VGND VGND VPWR VPWR _13626_/X sky130_fd_sc_hd__or3_4
XFILLER_20_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17394_ _17394_/A _17393_/X VGND VGND VPWR VPWR _17609_/D sky130_fd_sc_hd__or2_4
XFILLER_125_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19133_ _24312_/Q _19219_/A VGND VGND VPWR VPWR _19133_/X sky130_fd_sc_hd__and2_4
XANTENNA__21023__A _22169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16345_ _11784_/X _16337_/X _16344_/X VGND VGND VPWR VPWR _16345_/X sky130_fd_sc_hd__and3_4
X_13557_ _13543_/X _13469_/B VGND VGND VPWR VPWR _13559_/B sky130_fd_sc_hd__or2_4
XANTENNA__12645__A _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15021__A _13965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12508_ _12903_/A _12500_/X _12507_/X VGND VGND VPWR VPWR _12508_/X sky130_fd_sc_hd__and3_4
X_19064_ _11526_/X VGND VGND VPWR VPWR _19064_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13488_ _13531_/A _23269_/Q VGND VGND VPWR VPWR _13488_/X sky130_fd_sc_hd__or2_4
X_16276_ _15978_/A _16272_/X _16275_/X VGND VGND VPWR VPWR _16276_/X sky130_fd_sc_hd__or3_4
XFILLER_139_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18015_ _17664_/Y _18014_/X _17661_/X VGND VGND VPWR VPWR _18015_/X sky130_fd_sc_hd__o21a_4
XFILLER_173_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12439_ _12848_/A _12584_/B VGND VGND VPWR VPWR _12439_/X sky130_fd_sc_hd__or2_4
XFILLER_145_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15227_ _14196_/A _15227_/B VGND VGND VPWR VPWR _15227_/X sky130_fd_sc_hd__or2_4
XANTENNA__22245__A2 _22244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18449__B2 _18448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19428__A _19428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15158_ _15267_/A _15222_/B VGND VGND VPWR VPWR _15158_/X sky130_fd_sc_hd__or2_4
XANTENNA__17121__A1 _14845_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14109_ _14140_/A _23679_/Q VGND VGND VPWR VPWR _14112_/B sky130_fd_sc_hd__or2_4
XANTENNA__12380__A _13530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19887__A2_N _19886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19966_ _17793_/X _19966_/B _19966_/C _19966_/D VGND VGND VPWR VPWR _19966_/X sky130_fd_sc_hd__or4_4
X_15089_ _15096_/A _24053_/Q VGND VGND VPWR VPWR _15090_/C sky130_fd_sc_hd__or2_4
X_18917_ _13266_/X _18913_/X _24392_/Q _18914_/X VGND VGND VPWR VPWR _24392_/D sky130_fd_sc_hd__o22a_4
XFILLER_84_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19897_ _19607_/X _19896_/X _16936_/X _19571_/X VGND VGND VPWR VPWR _19897_/X sky130_fd_sc_hd__o22a_4
XFILLER_171_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16787__A _16053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18848_ _16523_/B _18840_/X _24432_/Q _18843_/X VGND VGND VPWR VPWR _18848_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16937__D _17087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18779_ _16915_/A VGND VGND VPWR VPWR _18779_/X sky130_fd_sc_hd__buf_2
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21508__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11724__A _12362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20810_ _20755_/X _20809_/X _11524_/A _20708_/X VGND VGND VPWR VPWR _20810_/X sky130_fd_sc_hd__o22a_4
X_21790_ _21575_/X _21784_/X _23648_/Q _21788_/X VGND VGND VPWR VPWR _23648_/D sky130_fd_sc_hd__o22a_4
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14100__A _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12539__B _12646_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22181__B2 _22177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20741_ _24257_/Q _20661_/X _20740_/X VGND VGND VPWR VPWR _20741_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19610__B HRDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23460_ _23588_/CLK _23460_/D VGND VGND VPWR VPWR _15682_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_11_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17411__A _17153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20672_ _20672_/A _20844_/B VGND VGND VPWR VPWR _20673_/C sky130_fd_sc_hd__or2_4
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22411_ _22404_/Y _22409_/X _22410_/X _22409_/X VGND VGND VPWR VPWR _22411_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23391_ _23391_/CLK _23391_/D VGND VGND VPWR VPWR _23391_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21692__B1 _23711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22342_ _22342_/A VGND VGND VPWR VPWR _23328_/D sky130_fd_sc_hd__buf_2
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20772__A _20772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24315__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14174__A1 _14302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22236__A2 _22230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22273_ _22090_/A _21656_/B _22637_/C _21236_/D VGND VGND VPWR VPWR _22273_/X sky130_fd_sc_hd__or4_4
X_24012_ _24012_/CLK _21151_/X VGND VGND VPWR VPWR _24012_/Q sky130_fd_sc_hd__dfxtp_4
X_21224_ _20860_/X _21219_/X _23964_/Q _21223_/X VGND VGND VPWR VPWR _23964_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21155_ _21155_/A VGND VGND VPWR VPWR _21155_/X sky130_fd_sc_hd__buf_2
XFILLER_105_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18860__A1 _13266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12290__A _12858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19397__A1_N _19396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20106_ _19979_/X _20104_/X _20105_/X _18622_/Y _19952_/Y VGND VGND VPWR VPWR _20106_/X
+ sky130_fd_sc_hd__a32o_4
X_21086_ _21101_/A VGND VGND VPWR VPWR _21086_/X sky130_fd_sc_hd__buf_2
XANTENNA__21747__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20037_ _18305_/X _20031_/X _20036_/Y _20018_/X VGND VGND VPWR VPWR _20037_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21108__A _21101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11810_ _11673_/A VGND VGND VPWR VPWR _15378_/A sky130_fd_sc_hd__inv_2
XANTENNA__15106__A _15106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12790_ _12801_/A _12790_/B VGND VGND VPWR VPWR _12790_/X sky130_fd_sc_hd__or2_4
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _23540_/Q VGND VGND VPWR VPWR _21988_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12449__B _23371_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _16465_/A VGND VGND VPWR VPWR _16056_/A sky130_fd_sc_hd__buf_2
XFILLER_27_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23727_ _23246_/CLK _23727_/D VGND VGND VPWR VPWR _16303_/B sky130_fd_sc_hd__dfxtp_4
X_20939_ _20894_/X _20938_/X _14751_/B _20861_/X VGND VGND VPWR VPWR _20939_/X sky130_fd_sc_hd__o22a_4
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20666__B _20665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14460_ _12455_/A _14460_/B VGND VGND VPWR VPWR _14460_/X sky130_fd_sc_hd__or2_4
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11664_/A VGND VGND VPWR VPWR _11673_/A sky130_fd_sc_hd__buf_2
X_23658_ _23723_/CLK _21776_/X VGND VGND VPWR VPWR _23658_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ _13378_/A _23238_/Q VGND VGND VPWR VPWR _13411_/X sky130_fd_sc_hd__or2_4
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22609_ _22437_/X _22608_/X _12935_/B _22605_/X VGND VGND VPWR VPWR _22609_/X sky130_fd_sc_hd__o22a_4
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _14510_/A _14391_/B VGND VGND VPWR VPWR _14393_/B sky130_fd_sc_hd__or2_4
X_23589_ _23241_/CLK _23589_/D VGND VGND VPWR VPWR _13447_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16130_ _16130_/A _16129_/X VGND VGND VPWR VPWR _16130_/X sky130_fd_sc_hd__and2_4
X_13342_ _13341_/X VGND VGND VPWR VPWR _13342_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16061_ _16061_/A _15988_/B VGND VGND VPWR VPWR _16061_/X sky130_fd_sc_hd__or2_4
X_13273_ _12559_/A _13273_/B VGND VGND VPWR VPWR _13273_/X sky130_fd_sc_hd__or2_4
XANTENNA__15776__A _12766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18152__A _18407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12224_ _12698_/A _12216_/X _12224_/C VGND VGND VPWR VPWR _12224_/X sky130_fd_sc_hd__and3_4
XFILLER_6_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15012_ _12467_/A _15010_/X _15011_/X VGND VGND VPWR VPWR _15013_/C sky130_fd_sc_hd__and3_4
XFILLER_155_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19820_ _19471_/X _19815_/X _19819_/Y _16915_/C _19512_/X VGND VGND VPWR VPWR _19820_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21986__B2 _21950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11809__A _16053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12155_ _11717_/X _12155_/B VGND VGND VPWR VPWR _12155_/X sky130_fd_sc_hd__or2_4
XANTENNA__18851__A1 _16381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19751_ _19539_/A _19532_/A _19588_/C VGND VGND VPWR VPWR _19752_/D sky130_fd_sc_hd__or3_4
X_16963_ _24143_/Q VGND VGND VPWR VPWR _16981_/A sky130_fd_sc_hd__inv_2
X_12086_ _12051_/A _12155_/B VGND VGND VPWR VPWR _12086_/X sky130_fd_sc_hd__or2_4
X_18702_ _17748_/X VGND VGND VPWR VPWR _18702_/Y sky130_fd_sc_hd__inv_2
X_15914_ _15849_/X _15913_/Y VGND VGND VPWR VPWR _15914_/X sky130_fd_sc_hd__or2_4
X_19682_ _19682_/A _19808_/A VGND VGND VPWR VPWR _19683_/B sky130_fd_sc_hd__or2_4
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16894_ _16824_/A _16893_/X _16824_/A _16893_/X VGND VGND VPWR VPWR _16895_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18633_ _17738_/X _18632_/Y _24137_/Q _18632_/A VGND VGND VPWR VPWR _18633_/X sky130_fd_sc_hd__o22a_4
XFILLER_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15845_ _12870_/A _15845_/B _15845_/C VGND VGND VPWR VPWR _15846_/C sky130_fd_sc_hd__and3_4
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15016__A _13952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18564_ _18518_/X _17412_/A _18519_/X VGND VGND VPWR VPWR _18564_/X sky130_fd_sc_hd__a21o_4
X_15776_ _12766_/X _15774_/X _15776_/C VGND VGND VPWR VPWR _15776_/X sky130_fd_sc_hd__and3_4
X_12988_ _12852_/A _12988_/B VGND VGND VPWR VPWR _12990_/B sky130_fd_sc_hd__or2_4
XANTENNA__20857__A _20857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17515_ _17165_/Y _17515_/B VGND VGND VPWR VPWR _17515_/X sky130_fd_sc_hd__and2_4
XFILLER_166_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14727_ _13990_/A _14727_/B VGND VGND VPWR VPWR _14727_/X sky130_fd_sc_hd__or2_4
X_18495_ _18477_/X _18482_/Y _18373_/X _18494_/X VGND VGND VPWR VPWR _18495_/X sky130_fd_sc_hd__o22a_4
X_11939_ _16138_/A VGND VGND VPWR VPWR _11939_/X sky130_fd_sc_hd__buf_2
XANTENNA__21910__A1 _21838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14855__A _13662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21910__B2 _21906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17446_ _17170_/Y _17446_/B VGND VGND VPWR VPWR _17446_/X sky130_fd_sc_hd__or2_4
X_14658_ _14658_/A _23546_/Q VGND VGND VPWR VPWR _14659_/C sky130_fd_sc_hd__or2_4
XFILLER_21_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17590__A1 _17120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13609_ _15423_/A _13713_/B VGND VGND VPWR VPWR _13609_/X sky130_fd_sc_hd__or2_4
XFILLER_20_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17377_ _17360_/A VGND VGND VPWR VPWR _17493_/A sky130_fd_sc_hd__buf_2
XFILLER_174_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12375__A _12923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14589_ _14310_/A _14585_/X _14588_/X VGND VGND VPWR VPWR _14589_/X sky130_fd_sc_hd__or3_4
X_19116_ _24376_/Q VGND VGND VPWR VPWR _19116_/Y sky130_fd_sc_hd__inv_2
X_16328_ _11684_/X _16328_/B _16328_/C VGND VGND VPWR VPWR _16328_/X sky130_fd_sc_hd__and3_4
XANTENNA__21688__A _21674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19047_ _11530_/A _11530_/B _19041_/Y VGND VGND VPWR VPWR _19047_/Y sky130_fd_sc_hd__a21oi_4
X_16259_ _16282_/A _16259_/B VGND VGND VPWR VPWR _16259_/X sky130_fd_sc_hd__or2_4
XANTENNA__22218__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14590__A _12530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24488__CLK _24294_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21977__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15656__A1 _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19605__B _19788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19949_ _11648_/X _11598_/X _18834_/C _19948_/X VGND VGND VPWR VPWR _19949_/X sky130_fd_sc_hd__or4_4
XANTENNA__22312__A _22291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21729__B2 _21724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13934__A _13720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22960_ _19438_/A VGND VGND VPWR VPWR _22961_/A sky130_fd_sc_hd__buf_2
XANTENNA__17406__A _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16310__A _13367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21911_ _21841_/X _21909_/X _23592_/Q _21906_/X VGND VGND VPWR VPWR _21911_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22891_ _22897_/A _22891_/B VGND VGND VPWR VPWR HWDATA[27] sky130_fd_sc_hd__nor2_4
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21842_ _21841_/X _21839_/X _23624_/Q _21834_/X VGND VGND VPWR VPWR _21842_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20767__A _20857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21773_ _21546_/X _21770_/X _23660_/Q _21767_/X VGND VGND VPWR VPWR _21773_/X sky130_fd_sc_hd__o22a_4
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21901__B2 _21899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20724_ _20778_/A _20724_/B VGND VGND VPWR VPWR _20724_/X sky130_fd_sc_hd__or2_4
XFILLER_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19570__A2 _19569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24396__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23512_ _23098_/CLK _23512_/D VGND VGND VPWR VPWR _23512_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24492_ _24277_/CLK _24492_/D HRESETn VGND VGND VPWR VPWR _20017_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_51_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23443_ _23475_/CLK _23443_/D VGND VGND VPWR VPWR _12159_/B sky130_fd_sc_hd__dfxtp_4
X_20655_ _20466_/X _20643_/Y _20653_/X _20654_/Y _20481_/X VGND VGND VPWR VPWR _20655_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_52_0_HCLK clkbuf_6_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23705__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23374_ _23501_/CLK _23374_/D VGND VGND VPWR VPWR _23374_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_109_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21598__A _21313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20586_ _20540_/X _20585_/X _24359_/Q _20547_/X VGND VGND VPWR VPWR _20586_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22325_ _16782_/B VGND VGND VPWR VPWR _23345_/D sky130_fd_sc_hd__buf_2
XANTENNA__22209__A2 _22208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22256_ _22141_/X _22251_/X _15562_/B _22255_/X VGND VGND VPWR VPWR _23393_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20007__A _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21207_ _20575_/X _21205_/X _23976_/Q _21202_/X VGND VGND VPWR VPWR _21207_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21968__B2 _21964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11629__A _11629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22187_ _22194_/A VGND VGND VPWR VPWR _22187_/X sky130_fd_sc_hd__buf_2
X_21138_ _21137_/X VGND VGND VPWR VPWR _21138_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_5_0_HCLK_A clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17316__A _14845_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21069_ _20841_/X _21066_/X _24061_/Q _21063_/X VGND VGND VPWR VPWR _24061_/D sky130_fd_sc_hd__o22a_4
XFILLER_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13960_ _13983_/A _23200_/Q VGND VGND VPWR VPWR _13960_/X sky130_fd_sc_hd__or2_4
XFILLER_24_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21196__A2 _21191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22393__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12911_ _12911_/A _12907_/X _12911_/C VGND VGND VPWR VPWR _12911_/X sky130_fd_sc_hd__or3_4
XANTENNA__24201__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13891_ _14507_/A _13811_/B VGND VGND VPWR VPWR _13891_/X sky130_fd_sc_hd__or2_4
XFILLER_47_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15630_ _15642_/A _15563_/B VGND VGND VPWR VPWR _15631_/C sky130_fd_sc_hd__or2_4
X_12842_ _13566_/A _12808_/X _12841_/X VGND VGND VPWR VPWR _12842_/X sky130_fd_sc_hd__and3_4
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18349__B1 _18176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22145__B2 _22142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15561_ _14418_/X _15559_/X _15560_/X VGND VGND VPWR VPWR _15561_/X sky130_fd_sc_hd__and3_4
XFILLER_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12773_ _12944_/A VGND VGND VPWR VPWR _12773_/X sky130_fd_sc_hd__buf_2
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22696__A2 _22694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _14844_/X _17300_/B VGND VGND VPWR VPWR _17300_/X sky130_fd_sc_hd__and2_4
X_14512_ _14512_/A _14512_/B _14512_/C VGND VGND VPWR VPWR _14513_/C sky130_fd_sc_hd__and3_4
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _12362_/A VGND VGND VPWR VPWR _13256_/A sky130_fd_sc_hd__buf_2
XFILLER_30_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18280_ _18406_/A _18280_/B VGND VGND VPWR VPWR _18283_/B sky130_fd_sc_hd__and2_4
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _12597_/A _15488_/X _15491_/X VGND VGND VPWR VPWR _15492_/X sky130_fd_sc_hd__or3_4
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17838_/A VGND VGND VPWR VPWR _17231_/X sky130_fd_sc_hd__buf_2
X_14443_ _14304_/A _14499_/B VGND VGND VPWR VPWR _14445_/B sky130_fd_sc_hd__or2_4
XFILLER_35_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11655_ _15595_/A VGND VGND VPWR VPWR _13923_/A sky130_fd_sc_hd__buf_2
XANTENNA__22448__A2 _22438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17162_ _17161_/X VGND VGND VPWR VPWR _17162_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14374_ _13229_/A _14358_/X _14373_/X VGND VGND VPWR VPWR _14412_/B sky130_fd_sc_hd__or3_4
X_11586_ _11549_/X _11559_/X _20111_/D _11585_/X VGND VGND VPWR VPWR _11586_/X sky130_fd_sc_hd__or4_4
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16113_ _16142_/A _16199_/B VGND VGND VPWR VPWR _16116_/B sky130_fd_sc_hd__or2_4
X_13325_ _13319_/A _23494_/Q VGND VGND VPWR VPWR _13325_/X sky130_fd_sc_hd__or2_4
X_17093_ _17092_/X VGND VGND VPWR VPWR _18008_/A sky130_fd_sc_hd__buf_2
XANTENNA__12923__A _12923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16044_ _11759_/X _16040_/X _16044_/C VGND VGND VPWR VPWR _16044_/X sky130_fd_sc_hd__or3_4
X_13256_ _13256_/A _23655_/Q VGND VGND VPWR VPWR _13257_/C sky130_fd_sc_hd__or2_4
XANTENNA__13738__B _13738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21959__B2 _21957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12207_ _12691_/A _12204_/X _12207_/C VGND VGND VPWR VPWR _12207_/X sky130_fd_sc_hd__and3_4
X_13187_ _12747_/A _23879_/Q VGND VGND VPWR VPWR _13187_/X sky130_fd_sc_hd__or2_4
XFILLER_151_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12138_ _12138_/A _12138_/B _12137_/X VGND VGND VPWR VPWR _12138_/X sky130_fd_sc_hd__or3_4
X_19803_ _19895_/A _19803_/B _19803_/C _19803_/D VGND VGND VPWR VPWR _19803_/X sky130_fd_sc_hd__or4_4
XFILLER_151_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22132__A _20632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17995_ _17986_/X _17993_/X _17988_/X _17994_/X VGND VGND VPWR VPWR _17996_/A sky130_fd_sc_hd__o22a_4
XFILLER_96_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13754__A _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19734_ _19474_/X HRDATA[5] VGND VGND VPWR VPWR _19734_/X sky130_fd_sc_hd__and2_4
X_16946_ _24160_/Q VGND VGND VPWR VPWR _17655_/A sky130_fd_sc_hd__inv_2
XANTENNA__17226__A _18538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12069_ _16742_/A _23603_/Q VGND VGND VPWR VPWR _12070_/C sky130_fd_sc_hd__or2_4
XANTENNA__16130__A _16130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18588__B1 _17792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22384__B2 _22380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19665_ _19665_/A _19665_/B VGND VGND VPWR VPWR _19828_/C sky130_fd_sc_hd__and2_4
XFILLER_38_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16877_ _14266_/B _16848_/X _14266_/B _16848_/X VGND VGND VPWR VPWR _16877_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20934__A2 _20231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18616_ _16975_/X VGND VGND VPWR VPWR _22935_/B sky130_fd_sc_hd__inv_2
X_15828_ _12440_/A _15826_/X _15827_/X VGND VGND VPWR VPWR _15828_/X sky130_fd_sc_hd__and3_4
X_19596_ _19546_/A _19681_/A _19678_/B VGND VGND VPWR VPWR _19596_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22136__B2 _22130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24160__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18547_ _18547_/A VGND VGND VPWR VPWR _18547_/Y sky130_fd_sc_hd__inv_2
X_15759_ _12780_/X _15759_/B VGND VGND VPWR VPWR _15759_/X sky130_fd_sc_hd__or2_4
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14585__A _14280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18057__A _18538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18478_ _18478_/A _18365_/X VGND VGND VPWR VPWR _18478_/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17429_ _14262_/X _17429_/B VGND VGND VPWR VPWR _17429_/X sky130_fd_sc_hd__or2_4
XANTENNA__22439__A2 _22438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20440_ _22110_/A VGND VGND VPWR VPWR _20441_/A sky130_fd_sc_hd__buf_2
XANTENNA__18512__B1 _18467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20371_ _20342_/X _20371_/B VGND VGND VPWR VPWR _20371_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13929__A _13916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12833__A _12833_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16305__A _11917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22110_ _22110_/A VGND VGND VPWR VPWR _22110_/X sky130_fd_sc_hd__buf_2
XFILLER_173_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23090_ VGND VGND VPWR VPWR _23090_/HI HTRANS[0] sky130_fd_sc_hd__conb_1
XANTENNA__12552__B _12657_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22041_ _22041_/A VGND VGND VPWR VPWR _22057_/A sky130_fd_sc_hd__inv_2
XFILLER_47_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18815__A1 _17169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22611__A2 _22608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22042__A _22057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13664__A _14331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16040__A _16056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23992_ _23290_/CLK _21179_/X VGND VGND VPWR VPWR _23992_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21178__A2 _21176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22977__A _22908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22375__B2 _22373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21881__A _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22943_ _22931_/A _22943_/B VGND VGND VPWR VPWR _22943_/X sky130_fd_sc_hd__and2_4
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22874_ _22874_/A VGND VGND VPWR VPWR HWDATA[23] sky130_fd_sc_hd__inv_2
XFILLER_44_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21825_ _21824_/X _21815_/X _16282_/B _21822_/X VGND VGND VPWR VPWR _21825_/X sky130_fd_sc_hd__o22a_4
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21756_ _22487_/A _21134_/D VGND VGND VPWR VPWR _21756_/X sky130_fd_sc_hd__or2_4
XANTENNA__21886__B1 _23605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21350__A2 _21348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20707_ _20644_/X _20706_/X _24290_/Q _20519_/X VGND VGND VPWR VPWR _20707_/X sky130_fd_sc_hd__o22a_4
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21687_ _21570_/X _21684_/X _23714_/Q _21681_/X VGND VGND VPWR VPWR _23714_/D sky130_fd_sc_hd__o22a_4
XFILLER_106_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24475_ _24471_/CLK _24475_/D HRESETn VGND VGND VPWR VPWR _24475_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23426_ _23523_/CLK _23426_/D VGND VGND VPWR VPWR _15497_/B sky130_fd_sc_hd__dfxtp_4
X_20638_ _20638_/A VGND VGND VPWR VPWR _20639_/A sky130_fd_sc_hd__buf_2
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21102__A2 _21097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13839__A _12504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23357_ _23518_/CLK _23357_/D VGND VGND VPWR VPWR _13876_/B sky130_fd_sc_hd__dfxtp_4
X_20569_ _18299_/X _20469_/X _20514_/X _20568_/Y VGND VGND VPWR VPWR _20569_/X sky130_fd_sc_hd__a211o_4
XFILLER_4_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13110_ _13085_/A _13110_/B VGND VGND VPWR VPWR _13111_/C sky130_fd_sc_hd__or2_4
X_22308_ _22275_/A VGND VGND VPWR VPWR _22308_/X sky130_fd_sc_hd__buf_2
XFILLER_124_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14090_ _12218_/A VGND VGND VPWR VPWR _14138_/A sky130_fd_sc_hd__buf_2
XFILLER_153_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23288_ _23290_/CLK _23288_/D VGND VGND VPWR VPWR _15264_/B sky130_fd_sc_hd__dfxtp_4
X_13041_ _12492_/A _13041_/B _13041_/C VGND VGND VPWR VPWR _13045_/B sky130_fd_sc_hd__and3_4
X_22239_ _22113_/X _22237_/X _16142_/B _22234_/X VGND VGND VPWR VPWR _22239_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18806__A1 _12980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22602__A2 _22601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_59_0_HCLK clkbuf_7_59_0_HCLK/A VGND VGND VPWR VPWR _24012_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23048__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16800_ _16759_/A _16798_/X _16799_/X VGND VGND VPWR VPWR _16800_/X sky130_fd_sc_hd__and3_4
XANTENNA__17046__A _17046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17780_ _17780_/A _17263_/Y VGND VGND VPWR VPWR _17959_/A sky130_fd_sc_hd__or2_4
X_14992_ _14988_/A _15059_/B VGND VGND VPWR VPWR _14992_/X sky130_fd_sc_hd__or2_4
XFILLER_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21791__A _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16731_ _12041_/A _16799_/B VGND VGND VPWR VPWR _16731_/X sky130_fd_sc_hd__or2_4
X_13943_ _13894_/A _13935_/X _13943_/C VGND VGND VPWR VPWR _13943_/X sky130_fd_sc_hd__and3_4
XFILLER_74_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19450_ _19450_/A VGND VGND VPWR VPWR _19767_/A sky130_fd_sc_hd__buf_2
X_16662_ _16662_/A _23858_/Q VGND VGND VPWR VPWR _16663_/C sky130_fd_sc_hd__or2_4
XFILLER_62_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13874_ _15318_/A VGND VGND VPWR VPWR _13888_/A sky130_fd_sc_hd__buf_2
X_18401_ _18307_/X _18398_/X _24485_/Q _18400_/X VGND VGND VPWR VPWR _24485_/D sky130_fd_sc_hd__a2bb2o_4
X_15613_ _15641_/A _15539_/B VGND VGND VPWR VPWR _15615_/B sky130_fd_sc_hd__or2_4
X_12825_ _12801_/A _12825_/B VGND VGND VPWR VPWR _12826_/C sky130_fd_sc_hd__or2_4
X_19381_ _19377_/A VGND VGND VPWR VPWR _19381_/X sky130_fd_sc_hd__buf_2
X_16593_ _16593_/A _23122_/Q VGND VGND VPWR VPWR _16593_/X sky130_fd_sc_hd__or2_4
XANTENNA__20200__A _20200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18332_ _18248_/X _23001_/B _18248_/X _23001_/B VGND VGND VPWR VPWR _18332_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15544_ _14421_/A _15602_/B VGND VGND VPWR VPWR _15544_/X sky130_fd_sc_hd__or2_4
XFILLER_163_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12756_ _13052_/A VGND VGND VPWR VPWR _13067_/A sky130_fd_sc_hd__buf_2
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17545__A1 _17452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12637__B _12514_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _15325_/A VGND VGND VPWR VPWR _11708_/A sky130_fd_sc_hd__buf_2
X_18263_ _18131_/X _18262_/X _18200_/X _17978_/X VGND VGND VPWR VPWR _18264_/A sky130_fd_sc_hd__o22a_4
X_15475_ _13051_/A _15473_/X _15474_/X VGND VGND VPWR VPWR _15475_/X sky130_fd_sc_hd__and3_4
XFILLER_124_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12687_ _12687_/A _12763_/B VGND VGND VPWR VPWR _12687_/X sky130_fd_sc_hd__or2_4
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _17145_/Y _17197_/X _13947_/X _17198_/X VGND VGND VPWR VPWR _17214_/X sky130_fd_sc_hd__o22a_4
X_14426_ _14430_/A _14488_/B VGND VGND VPWR VPWR _14426_/X sky130_fd_sc_hd__or2_4
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11638_ _11638_/A _11637_/X VGND VGND VPWR VPWR _11639_/A sky130_fd_sc_hd__and2_4
X_18194_ _18377_/A _17487_/X VGND VGND VPWR VPWR _18196_/C sky130_fd_sc_hd__nor2_4
XANTENNA__22127__A _20595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13749__A _13229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17145_ _12419_/X VGND VGND VPWR VPWR _17145_/Y sky130_fd_sc_hd__inv_2
X_14357_ _14522_/A _14351_/X _14356_/X VGND VGND VPWR VPWR _14357_/X sky130_fd_sc_hd__or3_4
XANTENNA__12653__A _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11569_ _11566_/X _11569_/B VGND VGND VPWR VPWR _11570_/B sky130_fd_sc_hd__or2_4
X_13308_ _13483_/A _13282_/X _13289_/X _13299_/X _13307_/X VGND VGND VPWR VPWR _13308_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_144_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17076_ _11644_/X _16921_/A _16918_/X VGND VGND VPWR VPWR _18772_/A sky130_fd_sc_hd__o21a_4
X_14288_ _12470_/A _14288_/B _14288_/C VGND VGND VPWR VPWR _14292_/B sky130_fd_sc_hd__and3_4
X_16027_ _16061_/A _23214_/Q VGND VGND VPWR VPWR _16027_/X sky130_fd_sc_hd__or2_4
X_13239_ _13223_/A _13237_/X _13238_/X VGND VGND VPWR VPWR _13239_/X sky130_fd_sc_hd__and3_4
XFILLER_131_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18273__A2 _18254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19470__B2 _19469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24123__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17978_ _17977_/X _17936_/X _17880_/X VGND VGND VPWR VPWR _17978_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14299__B _14363_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19717_ _19716_/X VGND VGND VPWR VPWR _19717_/Y sky130_fd_sc_hd__inv_2
X_16929_ _16927_/Y _17087_/A VGND VGND VPWR VPWR _16929_/X sky130_fd_sc_hd__or2_4
XFILLER_66_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19648_ _19647_/Y _19660_/A _19687_/D _19644_/Y VGND VGND VPWR VPWR _19649_/B sky130_fd_sc_hd__o22a_4
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22109__B2 _22106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19579_ _24173_/Q _19457_/A HRDATA[25] _19454_/A VGND VGND VPWR VPWR _19579_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21610_ _21617_/A VGND VGND VPWR VPWR _21610_/X sky130_fd_sc_hd__buf_2
XANTENNA__11732__A _11705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22590_ _22605_/A VGND VGND VPWR VPWR _22598_/A sky130_fd_sc_hd__buf_2
XANTENNA__21332__A2 _21327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21541_ _20441_/A VGND VGND VPWR VPWR _21541_/X sky130_fd_sc_hd__buf_2
XFILLER_166_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24260_ _24127_/CLK _24260_/D HRESETn VGND VGND VPWR VPWR _20654_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_18_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21472_ _21471_/X VGND VGND VPWR VPWR _21506_/A sky130_fd_sc_hd__buf_2
XFILLER_147_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23211_ _24012_/CLK _23211_/D VGND VGND VPWR VPWR _12599_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13659__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20423_ _20251_/X _20422_/X _20235_/X VGND VGND VPWR VPWR _20423_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21096__B2 _21094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24191_ _23383_/CLK _19847_/X HRESETn VGND VGND VPWR VPWR _17296_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12563__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23142_ _24102_/CLK _22663_/X VGND VGND VPWR VPWR _13316_/B sky130_fd_sc_hd__dfxtp_4
X_20354_ _20342_/X _20353_/X VGND VGND VPWR VPWR _20354_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__20780__A _20233_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23073_ _23078_/A _23073_/B VGND VGND VPWR VPWR _23075_/B sky130_fd_sc_hd__or2_4
X_20285_ _20273_/X _20284_/X _19257_/Y _20273_/X VGND VGND VPWR VPWR _20285_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21399__A2 _21398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22596__B2 _22591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22024_ _21991_/A VGND VGND VPWR VPWR _22024_/X sky130_fd_sc_hd__buf_2
XFILLER_142_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13394__A _13385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11907__A _11941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23975_ _24039_/CLK _23975_/D VGND VGND VPWR VPWR _23975_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14002__B _23648_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21020__A1 _20305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21020__B2 _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22926_ _22929_/A _22926_/B _22925_/X VGND VGND VPWR VPWR _22926_/X sky130_fd_sc_hd__and3_4
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21571__A2 _21566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22857_ _17327_/Y _22848_/X _22849_/X VGND VGND VPWR VPWR _22857_/X sky130_fd_sc_hd__o21a_4
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12738__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12610_ _12610_/A VGND VGND VPWR VPWR _12632_/A sky130_fd_sc_hd__buf_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15114__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21808_ _21808_/A VGND VGND VPWR VPWR _21834_/A sky130_fd_sc_hd__inv_2
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13590_ _12466_/A VGND VGND VPWR VPWR _13591_/A sky130_fd_sc_hd__buf_2
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22788_ _22766_/Y _22788_/B VGND VGND VPWR VPWR _22792_/B sky130_fd_sc_hd__or2_4
XANTENNA__12457__B _23755_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22520__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12541_ _12906_/A VGND VGND VPWR VPWR _12895_/A sky130_fd_sc_hd__buf_2
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21739_ _21572_/X _21734_/X _23681_/Q _21738_/X VGND VGND VPWR VPWR _23681_/D sky130_fd_sc_hd__o22a_4
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15260_ _14140_/A _15260_/B VGND VGND VPWR VPWR _15262_/B sky130_fd_sc_hd__or2_4
X_12472_ _12472_/A VGND VGND VPWR VPWR _12869_/A sky130_fd_sc_hd__buf_2
X_24458_ _23347_/CLK _18805_/X HRESETn VGND VGND VPWR VPWR _24458_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16750__A2 _11632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14211_ _14248_/A _23455_/Q VGND VGND VPWR VPWR _14212_/C sky130_fd_sc_hd__or2_4
Xclkbuf_5_22_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13569__A _13485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23409_ _23409_/CLK _23409_/D VGND VGND VPWR VPWR _16798_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_138_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15191_ _14191_/A _15191_/B _15191_/C VGND VGND VPWR VPWR _15192_/C sky130_fd_sc_hd__and3_4
XANTENNA__12473__A _12473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24389_ _24419_/CLK _18922_/X HRESETn VGND VGND VPWR VPWR _24389_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__20834__A1 _18590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ _12426_/A _14140_/X _14142_/C VGND VGND VPWR VPWR _14142_/X sky130_fd_sc_hd__and3_4
XANTENNA__20690__A _20535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22036__B1 _14850_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15784__A _15783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18950_ _18950_/A VGND VGND VPWR VPWR _18950_/Y sky130_fd_sc_hd__inv_2
X_14073_ _14073_/A _14071_/X _14073_/C VGND VGND VPWR VPWR _14073_/X sky130_fd_sc_hd__and3_4
XFILLER_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13024_ _12881_/A _13024_/B _13024_/C VGND VGND VPWR VPWR _13024_/X sky130_fd_sc_hd__or3_4
X_17901_ _17009_/A VGND VGND VPWR VPWR _17903_/A sky130_fd_sc_hd__buf_2
X_18881_ _14844_/X _18877_/X _24409_/Q _18878_/X VGND VGND VPWR VPWR _18881_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17832_ _17849_/A VGND VGND VPWR VPWR _17833_/A sky130_fd_sc_hd__buf_2
XFILLER_86_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23573__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17763_ _17720_/A _17723_/Y VGND VGND VPWR VPWR _17763_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19703__B HRDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14975_ _14916_/X _14973_/X _14975_/C VGND VGND VPWR VPWR _14975_/X sky130_fd_sc_hd__and3_4
XANTENNA__15008__B _23573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22410__A _20298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19502_ _19823_/A VGND VGND VPWR VPWR _19546_/A sky130_fd_sc_hd__buf_2
X_16714_ _16711_/A _16774_/B VGND VGND VPWR VPWR _16714_/X sky130_fd_sc_hd__or2_4
XFILLER_47_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13926_ _13720_/A _13924_/X _13926_/C VGND VGND VPWR VPWR _13927_/C sky130_fd_sc_hd__and3_4
X_17694_ _17905_/A _17493_/X VGND VGND VPWR VPWR _17694_/X sky130_fd_sc_hd__or2_4
XFILLER_48_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21562__A2 _21554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19433_ _19428_/A VGND VGND VPWR VPWR _19433_/X sky130_fd_sc_hd__buf_2
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16645_ _16658_/A _24018_/Q VGND VGND VPWR VPWR _16645_/X sky130_fd_sc_hd__or2_4
X_13857_ _15446_/A _23709_/Q VGND VGND VPWR VPWR _13859_/B sky130_fd_sc_hd__or2_4
XANTENNA__15024__A _13953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12808_ _13530_/A _12788_/X _12807_/X VGND VGND VPWR VPWR _12808_/X sky130_fd_sc_hd__or3_4
X_19364_ _19362_/X _18529_/X _19362_/X _20765_/A VGND VGND VPWR VPWR _24256_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16576_ _16556_/A _16576_/B _16576_/C VGND VGND VPWR VPWR _16577_/C sky130_fd_sc_hd__and3_4
X_13788_ _13788_/A VGND VGND VPWR VPWR _15398_/A sky130_fd_sc_hd__buf_2
XANTENNA__21314__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22511__B2 _22505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18315_ _18315_/A VGND VGND VPWR VPWR _18315_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15527_ _12236_/A _15525_/X _15527_/C VGND VGND VPWR VPWR _15528_/C sky130_fd_sc_hd__and3_4
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12739_ _13332_/A _12836_/B VGND VGND VPWR VPWR _12739_/X sky130_fd_sc_hd__or2_4
X_19295_ _19295_/A VGND VGND VPWR VPWR _19295_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18335__A _18335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18246_ _17681_/A _16989_/B _18217_/C VGND VGND VPWR VPWR _23020_/B sky130_fd_sc_hd__a21o_4
X_15458_ _15477_/A _15458_/B VGND VGND VPWR VPWR _15458_/X sky130_fd_sc_hd__or2_4
XANTENNA__15678__B _23940_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14409_ _13756_/A _14409_/B _14408_/X VGND VGND VPWR VPWR _14410_/C sky130_fd_sc_hd__or3_4
XANTENNA__21078__B2 _21042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18177_ _17490_/C _18175_/B _18176_/X VGND VGND VPWR VPWR _18177_/Y sky130_fd_sc_hd__a21oi_4
X_15389_ _15389_/A _15389_/B VGND VGND VPWR VPWR _15389_/X sky130_fd_sc_hd__and2_4
X_17128_ _17128_/A VGND VGND VPWR VPWR _17128_/X sky130_fd_sc_hd__buf_2
XFILLER_116_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15694__A _13277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17059_ _11644_/X _16915_/A _16921_/A _11645_/X VGND VGND VPWR VPWR _17059_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22578__B2 _22576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20070_ _19956_/A VGND VGND VPWR VPWR _20070_/X sky130_fd_sc_hd__buf_2
XANTENNA__20589__B1 _20538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_42_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR _24078_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__11727__A _11727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21250__B2 _21240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13942__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17414__A _17414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23760_ _23760_/CLK _23760_/D VGND VGND VPWR VPWR _16391_/B sky130_fd_sc_hd__dfxtp_4
X_20972_ _20343_/A _20971_/X _24311_/Q _20352_/A VGND VGND VPWR VPWR _20973_/B sky130_fd_sc_hd__o22a_4
XANTENNA__14757__B _14827_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22711_ _20596_/A _22708_/X _23111_/Q _22705_/X VGND VGND VPWR VPWR _23111_/D sky130_fd_sc_hd__o22a_4
XPHY_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23691_ _23558_/CLK _21725_/X VGND VGND VPWR VPWR _12500_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12558__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22642_ _22636_/Y _22641_/X _22410_/X _22641_/X VGND VGND VPWR VPWR _22642_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20775__A HRDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22502__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15869__A _13546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22573_ _22461_/X _22572_/X _23199_/Q _22569_/X VGND VGND VPWR VPWR _23199_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20513__B1 _20306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14773__A _14773_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24312_ _24287_/CLK _24312_/D HRESETn VGND VGND VPWR VPWR _24312_/Q sky130_fd_sc_hd__dfrtp_4
X_21524_ _21549_/A VGND VGND VPWR VPWR _21524_/X sky130_fd_sc_hd__buf_2
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21069__B2 _21063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24243_ _24471_/CLK _24243_/D HRESETn VGND VGND VPWR VPWR _24243_/Q sky130_fd_sc_hd__dfrtp_4
X_21455_ _21455_/A VGND VGND VPWR VPWR _21455_/X sky130_fd_sc_hd__buf_2
XANTENNA__12293__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11557__A1 _24458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20406_ _20315_/X _20405_/X _24367_/Q _20325_/X VGND VGND VPWR VPWR _20406_/X sky130_fd_sc_hd__o22a_4
X_24174_ _23383_/CLK _19933_/X HRESETn VGND VGND VPWR VPWR _24174_/Q sky130_fd_sc_hd__dfrtp_4
X_21386_ _21259_/X _21384_/X _23885_/Q _21381_/X VGND VGND VPWR VPWR _21386_/X sky130_fd_sc_hd__o22a_4
XFILLER_135_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20337_ _21528_/A VGND VGND VPWR VPWR _20337_/X sky130_fd_sc_hd__buf_2
X_23125_ _23456_/CLK _22685_/X VGND VGND VPWR VPWR _23125_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_116_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23056_ _23051_/A _23056_/B _23056_/C VGND VGND VPWR VPWR _23056_/X sky130_fd_sc_hd__and3_4
XFILLER_1_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20268_ _20267_/X VGND VGND VPWR VPWR _20269_/A sky130_fd_sc_hd__buf_2
XFILLER_88_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22007_ _22007_/A VGND VGND VPWR VPWR _22007_/X sky130_fd_sc_hd__buf_2
XANTENNA__19985__A2 _19983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15109__A _15081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20199_ _20154_/Y _19959_/A _20198_/X VGND VGND VPWR VPWR _20200_/B sky130_fd_sc_hd__o21a_4
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21792__A2 _21791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22230__A _22244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17324__A _15382_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13852__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14760_ _13627_/A _14760_/B VGND VGND VPWR VPWR _14762_/B sky130_fd_sc_hd__or2_4
X_11972_ _11971_/X VGND VGND VPWR VPWR _16130_/A sky130_fd_sc_hd__buf_2
X_23958_ _23416_/CLK _21231_/X VGND VGND VPWR VPWR _23958_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13711_ _15486_/A _13605_/B VGND VGND VPWR VPWR _13711_/X sky130_fd_sc_hd__or2_4
XFILLER_17_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22909_ _22742_/A VGND VGND VPWR VPWR _22909_/X sky130_fd_sc_hd__buf_2
XANTENNA__17043__B _17481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13571__B _13417_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14691_ _14691_/A _14597_/B VGND VGND VPWR VPWR _14691_/X sky130_fd_sc_hd__or2_4
X_23889_ _23889_/CLK _23889_/D VGND VGND VPWR VPWR _23889_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_71_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16430_ _15998_/X _16428_/X _16429_/X VGND VGND VPWR VPWR _16434_/B sky130_fd_sc_hd__and3_4
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24221__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13642_ _13642_/A VGND VGND VPWR VPWR _13652_/A sky130_fd_sc_hd__buf_2
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16361_ _11784_/X _16353_/X _16360_/X VGND VGND VPWR VPWR _16361_/X sky130_fd_sc_hd__and3_4
XANTENNA__15779__A _11701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20504__B1 _20714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _13272_/X _13573_/B VGND VGND VPWR VPWR _13573_/Y sky130_fd_sc_hd__nor2_4
XFILLER_158_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18155__A _18283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18100_ _18099_/A _18098_/X _18009_/X VGND VGND VPWR VPWR _18100_/Y sky130_fd_sc_hd__a21oi_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ _14302_/A _15289_/X _15296_/X _15303_/X _15311_/X VGND VGND VPWR VPWR _15312_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12524_ _12882_/A _12524_/B VGND VGND VPWR VPWR _12524_/X sky130_fd_sc_hd__and2_4
X_19080_ _19074_/X _19077_/X _19078_/Y _19079_/X VGND VGND VPWR VPWR _19080_/X sky130_fd_sc_hd__o22a_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _16159_/A _16292_/B _16291_/X VGND VGND VPWR VPWR _16292_/X sky130_fd_sc_hd__or3_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18031_ _18030_/X VGND VGND VPWR VPWR _18031_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13299__A _12516_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15243_ _14191_/A _15243_/B _15243_/C VGND VGND VPWR VPWR _15247_/B sky130_fd_sc_hd__and3_4
XFILLER_172_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12455_ _12455_/A VGND VGND VPWR VPWR _12876_/A sky130_fd_sc_hd__buf_2
XFILLER_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19673__A1 _19576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15174_ _13593_/A _15172_/X _15174_/C VGND VGND VPWR VPWR _15175_/C sky130_fd_sc_hd__and3_4
XFILLER_158_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12386_ _12363_/X _24076_/Q VGND VGND VPWR VPWR _12387_/C sky130_fd_sc_hd__or2_4
XFILLER_125_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14125_ _11929_/A VGND VGND VPWR VPWR _14133_/A sky130_fd_sc_hd__buf_2
XANTENNA__21480__B2 _21475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12931__A _12977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19982_ _19981_/X VGND VGND VPWR VPWR _19982_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18933_ _17272_/X _18927_/X _19094_/A _18928_/X VGND VGND VPWR VPWR _24380_/D sky130_fd_sc_hd__o22a_4
X_14056_ _14056_/A _24064_/Q VGND VGND VPWR VPWR _14057_/C sky130_fd_sc_hd__or2_4
XFILLER_79_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13007_ _12570_/A _13007_/B _13007_/C VGND VGND VPWR VPWR _13007_/X sky130_fd_sc_hd__and3_4
Xclkbuf_6_29_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15019__A _15000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21232__B2 _21195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18864_ _18842_/A VGND VGND VPWR VPWR _18864_/X sky130_fd_sc_hd__buf_2
XFILLER_121_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21783__A2 _21777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17815_ _17814_/X VGND VGND VPWR VPWR _17815_/X sky130_fd_sc_hd__buf_2
X_18795_ _16523_/B _18787_/X _24464_/Q _18790_/X VGND VGND VPWR VPWR _24464_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13762__A _12587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23319__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17746_ _17746_/A _17744_/A VGND VGND VPWR VPWR _17746_/X sky130_fd_sc_hd__or2_4
XANTENNA__22360__A2_N _22359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14958_ _14922_/A _14958_/B VGND VGND VPWR VPWR _14958_/X sky130_fd_sc_hd__or2_4
XFILLER_78_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21535__A2 _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14577__B _14649_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22732__B2 _22726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13909_ _13720_/A _13907_/X _13908_/X VGND VGND VPWR VPWR _13910_/C sky130_fd_sc_hd__and3_4
X_17677_ _18190_/A _17464_/X VGND VGND VPWR VPWR _17679_/A sky130_fd_sc_hd__nor2_4
XANTENNA__12378__A _15894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14889_ _11618_/A _14889_/B _14888_/X VGND VGND VPWR VPWR _14893_/B sky130_fd_sc_hd__and3_4
XFILLER_74_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16628_ _16646_/A _16624_/X _16627_/X VGND VGND VPWR VPWR _16629_/C sky130_fd_sc_hd__and3_4
X_19416_ _19414_/X _18436_/Y _19414_/X _24227_/Q VGND VGND VPWR VPWR _19416_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20595__A _20595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15689__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16559_ _16554_/X _23570_/Q VGND VGND VPWR VPWR _16560_/C sky130_fd_sc_hd__or2_4
X_19347_ _19340_/A VGND VGND VPWR VPWR _19347_/X sky130_fd_sc_hd__buf_2
XFILLER_149_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14593__A _14307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18065__A _18064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19361__B1 _19358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19278_ _19247_/A _19247_/B _19277_/Y VGND VGND VPWR VPWR _24298_/D sky130_fd_sc_hd__o21a_4
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19410__A2_N _18309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18229_ _18229_/A VGND VGND VPWR VPWR _18229_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13002__A _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21240_ _21239_/X VGND VGND VPWR VPWR _21240_/X sky130_fd_sc_hd__buf_2
XFILLER_11_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22315__A _22275_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21171_ _20819_/X _21169_/X _23998_/Q _21166_/X VGND VGND VPWR VPWR _21171_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17409__A _17153_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12841__A _13416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20122_ _20121_/Y _11549_/X _11564_/X VGND VGND VPWR VPWR _20122_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__19416__B2 _24227_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19624__A _19624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20053_ _20040_/X _17906_/A _20046_/X _20052_/X VGND VGND VPWR VPWR _20053_/X sky130_fd_sc_hd__o22a_4
XFILLER_58_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22050__A _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14768__A _15321_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23812_ _23523_/CLK _23812_/D VGND VGND VPWR VPWR _23812_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24244__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22985__A _18448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22723__A1 _20801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22723__B2 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23743_ _23679_/CLK _21642_/X VGND VGND VPWR VPWR _23743_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12288__A _12288_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20955_ _20305_/X _20946_/Y _20953_/X _20954_/Y _20255_/A VGND VGND VPWR VPWR _20955_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ _24090_/CLK _21749_/X VGND VGND VPWR VPWR _14567_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20885_/X VGND VGND VPWR VPWR _20886_/Y sky130_fd_sc_hd__inv_2
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22625_ _22466_/X _22622_/X _13900_/B _22619_/X VGND VGND VPWR VPWR _23165_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15599__A _15625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11920__A _16148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22556_ _22432_/X _22551_/X _12599_/B _22555_/X VGND VGND VPWR VPWR _23211_/D sky130_fd_sc_hd__o22a_4
XFILLER_167_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21507_ _21292_/X _21506_/X _23807_/Q _21503_/X VGND VGND VPWR VPWR _23807_/D sky130_fd_sc_hd__o22a_4
XFILLER_5_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22487_ _22487_/A _22487_/B VGND VGND VPWR VPWR _22487_/X sky130_fd_sc_hd__or2_4
XANTENNA__14008__A _12188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12240_ _12240_/A VGND VGND VPWR VPWR _13164_/A sky130_fd_sc_hd__buf_2
X_24226_ _24134_/CLK _19417_/X HRESETn VGND VGND VPWR VPWR _24226_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21438_ _21438_/A VGND VGND VPWR VPWR _21438_/X sky130_fd_sc_hd__buf_2
XFILLER_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22225__A _22258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12171_ _11746_/X _24115_/Q VGND VGND VPWR VPWR _12172_/C sky130_fd_sc_hd__or2_4
X_21369_ _23892_/Q VGND VGND VPWR VPWR _21369_/Y sky130_fd_sc_hd__inv_2
X_24157_ _24158_/CLK _20006_/Y HRESETn VGND VGND VPWR VPWR _16949_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17319__A _15382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23108_ _23908_/CLK _23108_/D VGND VGND VPWR VPWR _23108_/Q sky130_fd_sc_hd__dfxtp_4
X_24088_ _23290_/CLK _24088_/D VGND VGND VPWR VPWR _24088_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_107_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15930_ _15391_/X _15919_/X _15787_/X _15929_/Y VGND VGND VPWR VPWR _15931_/D sky130_fd_sc_hd__o22a_4
XFILLER_89_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21214__B2 _21209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23039_ _18178_/X _23055_/B VGND VGND VPWR VPWR _23040_/C sky130_fd_sc_hd__or2_4
XANTENNA__19534__A _19705_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21765__A2 _21763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15861_ _13540_/X _15800_/B VGND VGND VPWR VPWR _15861_/X sky130_fd_sc_hd__or2_4
XFILLER_40_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17600_ _17461_/X _18165_/B _17600_/C _17600_/D VGND VGND VPWR VPWR _17639_/A sky130_fd_sc_hd__or4_4
XFILLER_92_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17054__A _17015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14812_ _14819_/A _14736_/B VGND VGND VPWR VPWR _14812_/X sky130_fd_sc_hd__or2_4
X_18580_ _18575_/X _18579_/Y _17006_/A _18578_/X VGND VGND VPWR VPWR _18580_/X sky130_fd_sc_hd__o22a_4
X_15792_ _12847_/A _15853_/B VGND VGND VPWR VPWR _15792_/X sky130_fd_sc_hd__or2_4
XFILLER_57_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21517__A2 _21513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22714__B2 _22712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17531_ _17173_/Y _18334_/B VGND VGND VPWR VPWR _17531_/X sky130_fd_sc_hd__or2_4
X_14743_ _13652_/A _14743_/B VGND VGND VPWR VPWR _14743_/X sky130_fd_sc_hd__or2_4
X_11955_ _12012_/A VGND VGND VPWR VPWR _12103_/A sky130_fd_sc_hd__buf_2
XANTENNA__12198__A _12198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22190__A2 _22187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19591__B1 HRDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17462_ _17461_/X VGND VGND VPWR VPWR _17490_/A sky130_fd_sc_hd__inv_2
X_14674_ _14674_/A _14590_/B VGND VGND VPWR VPWR _14674_/X sky130_fd_sc_hd__or2_4
X_11886_ _11886_/A VGND VGND VPWR VPWR _11887_/A sky130_fd_sc_hd__buf_2
X_16413_ _16413_/A _16413_/B VGND VGND VPWR VPWR _16413_/X sky130_fd_sc_hd__or2_4
X_19201_ _19142_/B VGND VGND VPWR VPWR _19201_/Y sky130_fd_sc_hd__inv_2
X_13625_ _15404_/A _13625_/B _13624_/X VGND VGND VPWR VPWR _13626_/C sky130_fd_sc_hd__and3_4
X_17393_ _15913_/Y _17448_/B VGND VGND VPWR VPWR _17393_/X sky130_fd_sc_hd__and2_4
X_19132_ _24311_/Q _19131_/X VGND VGND VPWR VPWR _19219_/A sky130_fd_sc_hd__and2_4
XFILLER_164_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16344_ _13407_/A _16340_/X _16343_/X VGND VGND VPWR VPWR _16344_/X sky130_fd_sc_hd__or3_4
XANTENNA__23761__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15302__A _13593_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13556_ _13556_/A _13556_/B _13556_/C VGND VGND VPWR VPWR _13564_/B sky130_fd_sc_hd__or3_4
XFILLER_125_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12507_ _12872_/A _12632_/B VGND VGND VPWR VPWR _12507_/X sky130_fd_sc_hd__or2_4
X_19063_ _19063_/A VGND VGND VPWR VPWR _19063_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16275_ _11882_/X _16273_/X _16274_/X VGND VGND VPWR VPWR _16275_/X sky130_fd_sc_hd__and3_4
XFILLER_173_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13487_ _12948_/A VGND VGND VPWR VPWR _13531_/A sky130_fd_sc_hd__buf_2
XFILLER_9_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18014_ _17671_/B _18014_/B VGND VGND VPWR VPWR _18014_/X sky130_fd_sc_hd__and2_4
X_15226_ _14225_/A _15162_/B VGND VGND VPWR VPWR _15226_/X sky130_fd_sc_hd__or2_4
X_12438_ _12854_/A VGND VGND VPWR VPWR _12848_/A sky130_fd_sc_hd__buf_2
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22135__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24117__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15157_ _14272_/A _15157_/B _15157_/C VGND VGND VPWR VPWR _15157_/X sky130_fd_sc_hd__and3_4
XANTENNA__21453__B2 _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12369_ _11712_/X _23692_/Q VGND VGND VPWR VPWR _12369_/X sky130_fd_sc_hd__or2_4
XFILLER_141_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14108_ _14108_/A VGND VGND VPWR VPWR _14140_/A sky130_fd_sc_hd__buf_2
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21974__A _21941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19965_ _17801_/X _19965_/B VGND VGND VPWR VPWR _19966_/D sky130_fd_sc_hd__and2_4
X_15088_ _15095_/A _23605_/Q VGND VGND VPWR VPWR _15090_/B sky130_fd_sc_hd__or2_4
XFILLER_113_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18916_ _12980_/X _18913_/X _19020_/A _18914_/X VGND VGND VPWR VPWR _24393_/D sky130_fd_sc_hd__o22a_4
X_14039_ _12581_/A _14039_/B VGND VGND VPWR VPWR _14040_/C sky130_fd_sc_hd__or2_4
XANTENNA__24267__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19896_ _19516_/X _19724_/A _19895_/X VGND VGND VPWR VPWR _19896_/X sky130_fd_sc_hd__o21a_4
XFILLER_171_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18847_ _17266_/X _18840_/X _24433_/Q _18843_/X VGND VGND VPWR VPWR _18847_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14588__A _15394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13492__A _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18778_ _18667_/X _18777_/X _24469_/Q _18667_/X VGND VGND VPWR VPWR _18778_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21508__A2 _21506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17729_ _17729_/A VGND VGND VPWR VPWR _17730_/A sky130_fd_sc_hd__inv_2
XFILLER_36_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22181__A2 _22180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20740_ _20662_/X _20724_/X _20537_/X _20739_/Y VGND VGND VPWR VPWR _20740_/X sky130_fd_sc_hd__a211o_4
X_20671_ _20671_/A VGND VGND VPWR VPWR _20844_/B sky130_fd_sc_hd__buf_2
XFILLER_91_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18137__A1 _17594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11740__A _13377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15212__A _14616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22410_ _20298_/A VGND VGND VPWR VPWR _22410_/X sky130_fd_sc_hd__buf_2
XFILLER_149_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23390_ _23582_/CLK _22260_/X VGND VGND VPWR VPWR _13760_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12555__B _12668_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22341_ _15539_/B VGND VGND VPWR VPWR _22341_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22272_ _11745_/B VGND VGND VPWR VPWR _22272_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22045__A _22041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24011_ _23558_/CLK _21153_/X VGND VGND VPWR VPWR _12632_/B sky130_fd_sc_hd__dfxtp_4
X_21223_ _21202_/A VGND VGND VPWR VPWR _21223_/X sky130_fd_sc_hd__buf_2
XANTENNA__13667__A _15406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17139__A _16085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12571__A _12571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21444__B2 _21438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21154_ _20531_/X _21148_/X _24010_/Q _21152_/X VGND VGND VPWR VPWR _24010_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24356__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20105_ _11639_/A _18645_/X VGND VGND VPWR VPWR _20105_/X sky130_fd_sc_hd__or2_4
XFILLER_63_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19354__A _19340_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21085_ _21118_/A VGND VGND VPWR VPWR _21101_/A sky130_fd_sc_hd__inv_2
XFILLER_144_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21747__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20036_ _20036_/A VGND VGND VPWR VPWR _20036_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_12_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14498__A _11681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11915__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11634__B _11633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21987_ _21885_/X _21960_/A _23541_/Q _21950_/A VGND VGND VPWR VPWR _23541_/D sky130_fd_sc_hd__o22a_4
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23726_ _23501_/CLK _21671_/X VGND VGND VPWR VPWR _23726_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23784__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _13377_/A VGND VGND VPWR VPWR _16465_/A sky130_fd_sc_hd__buf_2
XFILLER_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20938_/A VGND VGND VPWR VPWR _20938_/X sky130_fd_sc_hd__buf_2
XANTENNA__20183__A1 _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23657_ _23241_/CLK _23657_/D VGND VGND VPWR VPWR _12902_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _13417_/A VGND VGND VPWR VPWR _11671_/X sky130_fd_sc_hd__buf_2
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12746__A _13183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _20869_/A VGND VGND VPWR VPWR _20869_/X sky130_fd_sc_hd__buf_2
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13410_/A _13410_/B _13410_/C VGND VGND VPWR VPWR _13414_/B sky130_fd_sc_hd__and3_4
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22608_ _22608_/A VGND VGND VPWR VPWR _22608_/X sky130_fd_sc_hd__buf_2
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14390_ _14390_/A VGND VGND VPWR VPWR _14510_/A sky130_fd_sc_hd__buf_2
X_23588_ _23588_/CLK _21917_/X VGND VGND VPWR VPWR _15735_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13341_ _11858_/A _11631_/A _13308_/X _11607_/A _13340_/X VGND VGND VPWR VPWR _13341_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17887__B1 _18562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21683__B2 _21681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22539_ _22539_/A VGND VGND VPWR VPWR _22555_/A sky130_fd_sc_hd__inv_2
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16060_ _11759_/X _16056_/X _16060_/C VGND VGND VPWR VPWR _16068_/B sky130_fd_sc_hd__or3_4
X_13272_ _13269_/X _13271_/X VGND VGND VPWR VPWR _13272_/X sky130_fd_sc_hd__or2_4
XFILLER_108_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15011_ _12450_/X _23445_/Q VGND VGND VPWR VPWR _15011_/X sky130_fd_sc_hd__or2_4
X_12223_ _12721_/A _12223_/B VGND VGND VPWR VPWR _12224_/C sky130_fd_sc_hd__or2_4
X_24209_ _23126_/CLK _19570_/Y HRESETn VGND VGND VPWR VPWR _17251_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21435__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22632__B1 _23160_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12481__A _12194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18300__B2 _18299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21986__A2 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12154_ _11760_/X _12150_/X _12153_/X VGND VGND VPWR VPWR _12162_/B sky130_fd_sc_hd__or3_4
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21476__A2_N _21475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15792__A _12847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19750_ _19750_/A _19619_/A _19642_/A _19816_/B VGND VGND VPWR VPWR _19752_/B sky130_fd_sc_hd__or4_4
X_16962_ _16962_/A VGND VGND VPWR VPWR _16982_/A sky130_fd_sc_hd__inv_2
X_12085_ _12078_/X _12085_/B _12085_/C VGND VGND VPWR VPWR _12085_/X sky130_fd_sc_hd__or3_4
XFILLER_104_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18701_ _17755_/X VGND VGND VPWR VPWR _18701_/Y sky130_fd_sc_hd__inv_2
X_15913_ _15912_/X VGND VGND VPWR VPWR _15913_/Y sky130_fd_sc_hd__inv_2
X_19681_ _19681_/A _19681_/B VGND VGND VPWR VPWR _19808_/A sky130_fd_sc_hd__or2_4
X_16893_ _16533_/X _16823_/X _16822_/A VGND VGND VPWR VPWR _16893_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20946__B1 _20262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15844_ _12906_/A _15844_/B VGND VGND VPWR VPWR _15845_/C sky130_fd_sc_hd__or2_4
X_18632_ _18632_/A VGND VGND VPWR VPWR _18632_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14201__A _14201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15775_ _15743_/X _15702_/B VGND VGND VPWR VPWR _15776_/C sky130_fd_sc_hd__or2_4
XFILLER_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18563_ _17807_/X _18203_/Y _17870_/X _18562_/X VGND VGND VPWR VPWR _18563_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15016__B _23893_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12987_ _12684_/X _12986_/X VGND VGND VPWR VPWR _12987_/X sky130_fd_sc_hd__or2_4
X_17514_ _17513_/X VGND VGND VPWR VPWR _18282_/B sky130_fd_sc_hd__inv_2
X_14726_ _14331_/A _14722_/X _14726_/C VGND VGND VPWR VPWR _14726_/X sky130_fd_sc_hd__or3_4
X_11938_ _16129_/A VGND VGND VPWR VPWR _16138_/A sky130_fd_sc_hd__buf_2
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18494_ _18483_/X _18488_/Y _18490_/X _18492_/X _18493_/Y VGND VGND VPWR VPWR _18494_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_166_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21910__A2 _21909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17445_ _15651_/X _17445_/B VGND VGND VPWR VPWR _17445_/Y sky130_fd_sc_hd__nand2_4
X_14657_ _14657_/A _14570_/B VGND VGND VPWR VPWR _14659_/B sky130_fd_sc_hd__or2_4
XANTENNA__12656__A _12610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11869_ _11869_/A VGND VGND VPWR VPWR _15449_/A sky130_fd_sc_hd__buf_2
XFILLER_14_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13608_ _13823_/A VGND VGND VPWR VPWR _15423_/A sky130_fd_sc_hd__buf_2
X_17376_ _18415_/B VGND VGND VPWR VPWR _17396_/B sky130_fd_sc_hd__inv_2
XANTENNA__21123__B1 _24028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14588_ _15394_/A _14586_/X _14587_/X VGND VGND VPWR VPWR _14588_/X sky130_fd_sc_hd__and3_4
XFILLER_159_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16327_ _13414_/A _16323_/X _16326_/X VGND VGND VPWR VPWR _16328_/C sky130_fd_sc_hd__or3_4
X_19115_ _19114_/Y _11516_/X _11519_/B VGND VGND VPWR VPWR _19115_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15967__A _15967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13539_ _13539_/A _13462_/B VGND VGND VPWR VPWR _13539_/X sky130_fd_sc_hd__or2_4
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14871__A _12473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18343__A _18411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19046_ _19016_/A VGND VGND VPWR VPWR _19046_/X sky130_fd_sc_hd__buf_2
X_16258_ _16123_/A _16256_/X _16257_/X VGND VGND VPWR VPWR _16262_/B sky130_fd_sc_hd__and3_4
XFILLER_118_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14590__B _14590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13487__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15209_ _14630_/A _15205_/X _15209_/C VGND VGND VPWR VPWR _15217_/B sky130_fd_sc_hd__or3_4
XANTENNA__22623__B1 _23167_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16189_ _16216_/A _16189_/B VGND VGND VPWR VPWR _16189_/X sky130_fd_sc_hd__or2_4
XANTENNA__12391__A _11701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21977__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23657__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15656__A2 _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19948_ _17816_/X _18888_/X VGND VGND VPWR VPWR _19948_/X sky130_fd_sc_hd__or2_4
XFILLER_101_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21729__A2 _21727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21209__A _21202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19879_ _19849_/A _19839_/A _19879_/C _19879_/D VGND VGND VPWR VPWR _19879_/X sky130_fd_sc_hd__and4_4
XANTENNA__20113__A _20112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21910_ _21838_/X _21909_/X _23593_/Q _21906_/X VGND VGND VPWR VPWR _21910_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15207__A _14669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11735__A _11735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22890_ _16452_/Y _22885_/X _22875_/X _22889_/X VGND VGND VPWR VPWR _22891_/B sky130_fd_sc_hd__o22a_4
XANTENNA__14111__A _15257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21841_ _20575_/A VGND VGND VPWR VPWR _21841_/X sky130_fd_sc_hd__buf_2
XFILLER_82_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21772_ _21544_/X _21770_/X _16150_/B _21767_/X VGND VGND VPWR VPWR _21772_/X sky130_fd_sc_hd__o22a_4
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21901__A2 _21895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24500__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23511_ _23511_/CLK _22035_/X VGND VGND VPWR VPWR _15123_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20723_ _20664_/A _20721_/X _20722_/X VGND VGND VPWR VPWR _20724_/B sky130_fd_sc_hd__and3_4
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24491_ _24277_/CLK _24491_/D HRESETn VGND VGND VPWR VPWR _20023_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12566__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23442_ _23204_/CLK _22182_/X VGND VGND VPWR VPWR _16665_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21114__B1 _15465_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20654_ _20654_/A VGND VGND VPWR VPWR _20654_/Y sky130_fd_sc_hd__inv_2
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_3_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__15877__A _13547_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23373_ _24045_/CLK _23373_/D VGND VGND VPWR VPWR _23373_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21665__B2 _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20585_ _20490_/X _20583_/Y _24295_/Q _20584_/X VGND VGND VPWR VPWR _20585_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22324_ _23346_/Q VGND VGND VPWR VPWR _23346_/D sky130_fd_sc_hd__buf_2
XFILLER_104_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13397__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21417__B2 _21381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22255_ _22226_/A VGND VGND VPWR VPWR _22255_/X sky130_fd_sc_hd__buf_2
XFILLER_118_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21968__A2 _21967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21206_ _20559_/X _21205_/X _23977_/Q _21202_/X VGND VGND VPWR VPWR _23977_/D sky130_fd_sc_hd__o22a_4
XFILLER_133_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22186_ _22108_/X _22180_/X _16290_/B _22184_/X VGND VGND VPWR VPWR _23439_/D sky130_fd_sc_hd__o22a_4
XFILLER_79_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21137_ _21152_/A VGND VGND VPWR VPWR _21137_/X sky130_fd_sc_hd__buf_2
XFILLER_120_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21068_ _20819_/X _21066_/X _24062_/Q _21063_/X VGND VGND VPWR VPWR _24062_/D sky130_fd_sc_hd__o22a_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22393__A2 _22390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ _12870_/A _12908_/X _12909_/X VGND VGND VPWR VPWR _12911_/C sky130_fd_sc_hd__and3_4
XFILLER_24_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20019_ _18185_/X _20007_/X _20017_/Y _20018_/X VGND VGND VPWR VPWR _20019_/X sky130_fd_sc_hd__o22a_4
XFILLER_58_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14021__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13890_ _13877_/A VGND VGND VPWR VPWR _14507_/A sky130_fd_sc_hd__buf_2
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20958__A _20958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12841_ _13416_/A _12823_/X _12840_/X VGND VGND VPWR VPWR _12841_/X sky130_fd_sc_hd__or3_4
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22145__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13860__A _14331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15560_ _12304_/A _15560_/B VGND VGND VPWR VPWR _15560_/X sky130_fd_sc_hd__or2_4
XANTENNA__17332__A _15252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12772_ _12976_/A VGND VGND VPWR VPWR _13563_/A sky130_fd_sc_hd__buf_2
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13830__A1 _14480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14511_/A _14440_/B VGND VGND VPWR VPWR _14512_/C sky130_fd_sc_hd__or2_4
XFILLER_42_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23709_ _23646_/CLK _23709_/D VGND VGND VPWR VPWR _23709_/Q sky130_fd_sc_hd__dfxtp_4
X_11723_ _14658_/A VGND VGND VPWR VPWR _12362_/A sky130_fd_sc_hd__buf_2
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _12621_/X _15491_/B _15491_/C VGND VGND VPWR VPWR _15491_/X sky130_fd_sc_hd__and3_4
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_19_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR _24240_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12476__A _14325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17230_ _17836_/A VGND VGND VPWR VPWR _17230_/X sky130_fd_sc_hd__buf_2
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _12546_/A _14442_/B _14441_/X VGND VGND VPWR VPWR _14442_/X sky130_fd_sc_hd__or3_4
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11654_/A VGND VGND VPWR VPWR _15595_/A sky130_fd_sc_hd__buf_2
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20459__A2 _20445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17161_ _14084_/X VGND VGND VPWR VPWR _17161_/X sky130_fd_sc_hd__buf_2
XANTENNA__15787__A _15717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14373_ _12616_/A _14365_/X _14373_/C VGND VGND VPWR VPWR _14373_/X sky130_fd_sc_hd__and3_4
XFILLER_7_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ _11572_/X _11574_/X _20119_/A _11585_/D VGND VGND VPWR VPWR _11585_/X sky130_fd_sc_hd__or4_4
XFILLER_128_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16112_ _16112_/A VGND VGND VPWR VPWR _16142_/A sky130_fd_sc_hd__buf_2
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _13324_/A VGND VGND VPWR VPWR _13327_/A sky130_fd_sc_hd__buf_2
XFILLER_156_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17092_ _17090_/X _17091_/X _17912_/A VGND VGND VPWR VPWR _17092_/X sky130_fd_sc_hd__or3_4
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16043_ _16035_/A _16041_/X _16042_/X VGND VGND VPWR VPWR _16044_/C sky130_fd_sc_hd__and3_4
XFILLER_157_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13255_ _13248_/A _13179_/B VGND VGND VPWR VPWR _13255_/X sky130_fd_sc_hd__or2_4
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21959__A2 _21953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13100__A _13100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12206_ _12687_/A _23756_/Q VGND VGND VPWR VPWR _12207_/C sky130_fd_sc_hd__or2_4
X_13186_ _11887_/A _23719_/Q VGND VGND VPWR VPWR _13188_/B sky130_fd_sc_hd__or2_4
XFILLER_124_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22413__A _22462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19802_ _19819_/A _19801_/X VGND VGND VPWR VPWR _19803_/D sky130_fd_sc_hd__and2_4
X_12137_ _11834_/A _12135_/X _12136_/X VGND VGND VPWR VPWR _12137_/X sky130_fd_sc_hd__and3_4
XFILLER_150_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16411__A _16159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17994_ _17922_/X _17861_/X _17815_/X _17851_/X VGND VGND VPWR VPWR _17994_/X sky130_fd_sc_hd__o22a_4
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19733_ HRDATA[21] VGND VGND VPWR VPWR _20512_/B sky130_fd_sc_hd__buf_2
XANTENNA__21029__A _21081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16945_ _16945_/A VGND VGND VPWR VPWR _16945_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12068_ _16741_/A _23955_/Q VGND VGND VPWR VPWR _12070_/B sky130_fd_sc_hd__or2_4
XANTENNA__20919__B1 HRDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22384__A2 _22383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19722__A HRDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19664_ _19663_/Y VGND VGND VPWR VPWR _19665_/A sky130_fd_sc_hd__buf_2
X_16876_ _14417_/X _16875_/X _14417_/X _16875_/X VGND VGND VPWR VPWR _16876_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24329__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18615_ _18577_/X VGND VGND VPWR VPWR _18615_/Y sky130_fd_sc_hd__inv_2
X_15827_ _12860_/A _15827_/B VGND VGND VPWR VPWR _15827_/X sky130_fd_sc_hd__or2_4
XANTENNA__24305__CLK _24306_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19595_ _19681_/B VGND VGND VPWR VPWR _19678_/B sky130_fd_sc_hd__inv_2
XANTENNA__22136__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17242__A _12077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14613__A3 _14582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15758_ _11755_/X _15758_/B _15757_/X VGND VGND VPWR VPWR _15758_/X sky130_fd_sc_hd__or3_4
X_18546_ _17432_/X _18544_/X _17792_/X _18545_/X VGND VGND VPWR VPWR _18547_/A sky130_fd_sc_hd__a211o_4
XFILLER_80_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14709_ _13596_/A _14779_/B VGND VGND VPWR VPWR _14709_/X sky130_fd_sc_hd__or2_4
X_15689_ _12722_/A _15687_/X _15689_/C VGND VGND VPWR VPWR _15689_/X sky130_fd_sc_hd__and3_4
X_18477_ _16941_/X VGND VGND VPWR VPWR _18477_/X sky130_fd_sc_hd__buf_2
XANTENNA__18760__A1 _18757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17428_ _17425_/Y _17354_/X _17028_/X _17427_/X VGND VGND VPWR VPWR _17429_/B sky130_fd_sc_hd__o22a_4
XFILLER_20_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15697__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21647__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17359_ _16902_/A _17378_/A _17358_/Y VGND VGND VPWR VPWR _17360_/B sky130_fd_sc_hd__o21a_4
XANTENNA__18512__A1 _18413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20370_ _20343_/X _20369_/X _19158_/A _20352_/X VGND VGND VPWR VPWR _20371_/B sky130_fd_sc_hd__o22a_4
XFILLER_146_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19029_ _24359_/Q VGND VGND VPWR VPWR _19029_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14106__A _14003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13010__A _13010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20607__C1 _20606_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22040_ _22039_/X VGND VGND VPWR VPWR _22041_/A sky130_fd_sc_hd__buf_2
XFILLER_138_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22072__B2 _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20622__A2 _20621_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13945__A _11668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23991_ _23991_/CLK _23991_/D VGND VGND VPWR VPWR _15211_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22375__A2 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22942_ _22929_/A _24138_/Q VGND VGND VPWR VPWR _22942_/X sky130_fd_sc_hd__or2_4
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22873_ _12320_/Y _22846_/X _22799_/X _22872_/X VGND VGND VPWR VPWR _22874_/A sky130_fd_sc_hd__a211o_4
XFILLER_3_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14776__A _15076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13680__A _12300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17152__A _13781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21824_ _21824_/A VGND VGND VPWR VPWR _21824_/X sky130_fd_sc_hd__buf_2
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21755_ _23668_/Q VGND VGND VPWR VPWR _21755_/Y sky130_fd_sc_hd__inv_2
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21886__B2 _21809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12296__A _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20706_ _20703_/X _20705_/X _24386_/Q _20647_/X VGND VGND VPWR VPWR _20706_/X sky130_fd_sc_hd__o22a_4
XFILLER_93_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24474_ _23126_/CLK _18668_/X HRESETn VGND VGND VPWR VPWR _24474_/Q sky130_fd_sc_hd__dfrtp_4
X_21686_ _21568_/X _21684_/X _15843_/B _21681_/X VGND VGND VPWR VPWR _21686_/X sky130_fd_sc_hd__o22a_4
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21402__A _21388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23425_ _23617_/CLK _22206_/X VGND VGND VPWR VPWR _15563_/B sky130_fd_sc_hd__dfxtp_4
X_20637_ _20226_/X VGND VGND VPWR VPWR _20857_/A sky130_fd_sc_hd__buf_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15400__A _15400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23356_ _23772_/CLK _22313_/X VGND VGND VPWR VPWR _14343_/B sky130_fd_sc_hd__dfxtp_4
X_20568_ _20388_/A _20567_/X VGND VGND VPWR VPWR _20568_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__20018__A _19950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22307_ _22144_/X _22301_/X _23360_/Q _22305_/X VGND VGND VPWR VPWR _23360_/D sky130_fd_sc_hd__o22a_4
X_23287_ _23383_/CLK _22401_/X VGND VGND VPWR VPWR _15136_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_124_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20499_ _20315_/X _20498_/X _19004_/A _20325_/X VGND VGND VPWR VPWR _20499_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18711__A _17974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13040_ _12540_/A _13110_/B VGND VGND VPWR VPWR _13041_/C sky130_fd_sc_hd__or2_4
XFILLER_124_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22238_ _22110_/X _22237_/X _23406_/Q _22234_/X VGND VGND VPWR VPWR _23406_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22063__B2 _22057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13855__A _15444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17327__A _15185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22169_ _22169_/A VGND VGND VPWR VPWR _22169_/X sky130_fd_sc_hd__buf_2
XFILLER_152_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23202__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24328__CLK _24342_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14991_ _14991_/A _14987_/X _14991_/C VGND VGND VPWR VPWR _14991_/X sky130_fd_sc_hd__or3_4
XANTENNA__24493__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13942_ _12596_/A _13942_/B _13942_/C VGND VGND VPWR VPWR _13943_/C sky130_fd_sc_hd__or3_4
XFILLER_8_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16730_ _16704_/A _16798_/B VGND VGND VPWR VPWR _16730_/X sky130_fd_sc_hd__or2_4
XANTENNA__24422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16661_ _16654_/A _16661_/B VGND VGND VPWR VPWR _16661_/X sky130_fd_sc_hd__or2_4
XFILLER_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13873_ _15325_/A VGND VGND VPWR VPWR _15318_/A sky130_fd_sc_hd__buf_2
XANTENNA__14686__A _14657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18400_ _18399_/X VGND VGND VPWR VPWR _18400_/X sky130_fd_sc_hd__buf_2
XFILLER_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13590__A _12466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15612_ _15612_/A _15612_/B _15612_/C VGND VGND VPWR VPWR _15612_/X sky130_fd_sc_hd__and3_4
X_12824_ _12800_/A _12824_/B VGND VGND VPWR VPWR _12824_/X sky130_fd_sc_hd__or2_4
XANTENNA__24478__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19380_ _19377_/X _18741_/X _19377_/X _24246_/Q VGND VGND VPWR VPWR _19380_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16592_ _16592_/A _16592_/B _16592_/C VGND VGND VPWR VPWR _16592_/X sky130_fd_sc_hd__or3_4
XFILLER_43_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18331_ _16958_/A _18248_/C _16986_/X VGND VGND VPWR VPWR _23001_/B sky130_fd_sc_hd__o21a_4
X_15543_ _12213_/A _15601_/B VGND VGND VPWR VPWR _15543_/X sky130_fd_sc_hd__or2_4
X_12755_ _12975_/A VGND VGND VPWR VPWR _13562_/A sky130_fd_sc_hd__buf_2
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18742__B2 _18741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11706_/A VGND VGND VPWR VPWR _15325_/A sky130_fd_sc_hd__buf_2
X_18262_ _17856_/X _17930_/Y _17985_/X _17940_/Y VGND VGND VPWR VPWR _18262_/X sky130_fd_sc_hd__o22a_4
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _12626_/A _15474_/B VGND VGND VPWR VPWR _15474_/X sky130_fd_sc_hd__or2_4
X_12686_ _12568_/A _12759_/B VGND VGND VPWR VPWR _12688_/B sky130_fd_sc_hd__or2_4
XANTENNA__22408__A _22433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _12435_/A _14487_/B VGND VGND VPWR VPWR _14427_/B sky130_fd_sc_hd__or2_4
X_17213_ _17114_/X _17211_/X _17119_/X _17212_/X VGND VGND VPWR VPWR _17213_/X sky130_fd_sc_hd__o22a_4
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21629__B2 _21624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11637_ _24405_/Q _11587_/X NMI _11636_/Y VGND VGND VPWR VPWR _11637_/X sky130_fd_sc_hd__a211o_4
X_18193_ _18037_/X _17487_/B VGND VGND VPWR VPWR _18196_/B sky130_fd_sc_hd__nor2_4
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12934__A _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15310__A _15029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17144_ _17144_/A VGND VGND VPWR VPWR _17144_/X sky130_fd_sc_hd__buf_2
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _14383_/A _14356_/B _14355_/X VGND VGND VPWR VPWR _14356_/X sky130_fd_sc_hd__and3_4
X_11568_ _24448_/Q IRQ[11] _11567_/X VGND VGND VPWR VPWR _11569_/B sky130_fd_sc_hd__a21o_4
XFILLER_144_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13307_ _13307_/A _13306_/X VGND VGND VPWR VPWR _13307_/X sky130_fd_sc_hd__and2_4
X_17075_ _17074_/X VGND VGND VPWR VPWR _17075_/X sky130_fd_sc_hd__buf_2
XFILLER_128_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14287_ _15400_/A _23996_/Q VGND VGND VPWR VPWR _14288_/C sky130_fd_sc_hd__or2_4
X_16026_ _11693_/X _16019_/X _16026_/C VGND VGND VPWR VPWR _16026_/X sky130_fd_sc_hd__or3_4
X_13238_ _13200_/X _23847_/Q VGND VGND VPWR VPWR _13238_/X sky130_fd_sc_hd__or2_4
XANTENNA__22054__B2 _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21801__A1 _21594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13169_ _13301_/A _23847_/Q VGND VGND VPWR VPWR _13169_/X sky130_fd_sc_hd__or2_4
XANTENNA__21801__B2 _21795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16141__A _16110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17977_ _17876_/X VGND VGND VPWR VPWR _17977_/X sky130_fd_sc_hd__buf_2
XFILLER_46_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19758__B1 _20917_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19452__A _17005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19716_ _19647_/Y _19709_/X _19684_/X _19714_/X _19715_/X VGND VGND VPWR VPWR _19716_/X
+ sky130_fd_sc_hd__a32o_4
X_16928_ _17038_/B VGND VGND VPWR VPWR _17087_/A sky130_fd_sc_hd__inv_2
XANTENNA__24163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19647_ _19888_/B VGND VGND VPWR VPWR _19647_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16859_ _12986_/B _16832_/X _12986_/B _16832_/X VGND VGND VPWR VPWR _16884_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22109__A2 _22099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18068__A _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14596__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19578_ _19899_/B VGND VGND VPWR VPWR _19578_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18529_ _17720_/X _18528_/X _17720_/X _18528_/X VGND VGND VPWR VPWR _18529_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21868__B2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13005__A _12510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21540_ _21539_/X _21530_/X _16257_/B _21537_/X VGND VGND VPWR VPWR _23791_/D sky130_fd_sc_hd__o22a_4
XFILLER_61_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_65_0_HCLK clkbuf_7_65_0_HCLK/A VGND VGND VPWR VPWR _24248_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21471_ _21806_/A _21370_/B _21134_/C _21134_/D VGND VGND VPWR VPWR _21471_/X sky130_fd_sc_hd__or4_4
XFILLER_140_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12844__A _12753_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23210_ _23531_/CLK _23210_/D VGND VGND VPWR VPWR _12774_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21096__A2 _21090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23995__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20422_ _20380_/A _20422_/B VGND VGND VPWR VPWR _20422_/X sky130_fd_sc_hd__and2_4
XANTENNA__22293__B2 _22291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24190_ _23862_/CLK _19855_/Y HRESETn VGND VGND VPWR VPWR _21028_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_147_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23141_ _23397_/CLK _23141_/D VGND VGND VPWR VPWR _13462_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20353_ _20343_/X _20351_/X _19159_/A _20352_/X VGND VGND VPWR VPWR _20353_/X sky130_fd_sc_hd__o22a_4
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18531__A _18399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23072_ _23071_/X VGND VGND VPWR VPWR HADDR[29] sky130_fd_sc_hd__inv_2
X_20284_ _20277_/X _20283_/X _24404_/Q _18894_/B VGND VGND VPWR VPWR _20284_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22053__A _22060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22596__A2 _22594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22023_ _21860_/X _22017_/X _23520_/Q _22021_/X VGND VGND VPWR VPWR _23520_/D sky130_fd_sc_hd__o22a_4
XFILLER_103_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22988__A _22987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21892__A _21899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15890__A _13542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23974_ _24102_/CLK _23974_/D VGND VGND VPWR VPWR _23974_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22925_ _18681_/X _22930_/A VGND VGND VPWR VPWR _22925_/X sky130_fd_sc_hd__or2_4
XANTENNA__21020__A2 _21011_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20301__A _20772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11923__A _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22856_ _22856_/A VGND VGND VPWR VPWR HWDATA[17] sky130_fd_sc_hd__inv_2
XFILLER_169_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21807_ _21806_/X VGND VGND VPWR VPWR _21808_/A sky130_fd_sc_hd__buf_2
XANTENNA__21859__B2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22787_ _22787_/A _22788_/B _22793_/A VGND VGND VPWR VPWR _24122_/D sky130_fd_sc_hd__and3_4
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17032__D _17087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12540_ _12540_/A VGND VGND VPWR VPWR _12906_/A sky130_fd_sc_hd__buf_2
X_21738_ _21724_/A VGND VGND VPWR VPWR _21738_/X sky130_fd_sc_hd__buf_2
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12471_ _12492_/A VGND VGND VPWR VPWR _12472_/A sky130_fd_sc_hd__buf_2
XFILLER_12_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24457_ _23347_/CLK _24457_/D HRESETn VGND VGND VPWR VPWR _11556_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12754__A _12945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21669_ _21539_/X _21663_/X _16303_/B _21667_/X VGND VGND VPWR VPWR _23727_/D sky130_fd_sc_hd__o22a_4
XFILLER_138_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14210_ _13868_/A VGND VGND VPWR VPWR _14248_/A sky130_fd_sc_hd__buf_2
X_23408_ _24080_/CLK _23408_/D VGND VGND VPWR VPWR _16431_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15130__A _15257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15190_ _14665_/A _23735_/Q VGND VGND VPWR VPWR _15191_/C sky130_fd_sc_hd__or2_4
XFILLER_165_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24388_ _24388_/CLK _24388_/D HRESETn VGND VGND VPWR VPWR _24388_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_126_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14141_ _11898_/A _24063_/Q VGND VGND VPWR VPWR _14142_/C sky130_fd_sc_hd__or2_4
X_23339_ _23241_/CLK _23339_/D VGND VGND VPWR VPWR _23339_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22036__B2 _22000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14072_ _12329_/A _23872_/Q VGND VGND VPWR VPWR _14073_/C sky130_fd_sc_hd__or2_4
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24150__CLK _24302_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13023_ _12493_/A _13021_/X _13022_/X VGND VGND VPWR VPWR _13024_/C sky130_fd_sc_hd__and3_4
XFILLER_140_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17900_ _17900_/A VGND VGND VPWR VPWR _17900_/X sky130_fd_sc_hd__buf_2
XFILLER_156_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18880_ _17290_/X _18877_/X _24410_/Q _18878_/X VGND VGND VPWR VPWR _24410_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17831_ _12077_/X VGND VGND VPWR VPWR _17849_/A sky130_fd_sc_hd__buf_2
XFILLER_86_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17762_ _17729_/A _17762_/B _17762_/C VGND VGND VPWR VPWR _17762_/X sky130_fd_sc_hd__and3_4
XANTENNA__21547__B1 _23788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14974_ _14970_/A _14895_/B VGND VGND VPWR VPWR _14975_/C sky130_fd_sc_hd__or2_4
XFILLER_59_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19501_ _19504_/B _19548_/B _19537_/B VGND VGND VPWR VPWR _19558_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__17215__A1 _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16713_ _16713_/A _16711_/X _16713_/C VGND VGND VPWR VPWR _16717_/B sky130_fd_sc_hd__and3_4
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13925_ _13937_/A _13842_/B VGND VGND VPWR VPWR _13926_/C sky130_fd_sc_hd__or2_4
X_17693_ _16986_/A _17501_/X VGND VGND VPWR VPWR _17693_/X sky130_fd_sc_hd__or2_4
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12929__A _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17766__A2 _17368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19432_ _19428_/X _18719_/X _19428_/X _24215_/Q VGND VGND VPWR VPWR _19432_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15305__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13856_ _11878_/A _13856_/B _13855_/X VGND VGND VPWR VPWR _13856_/X sky130_fd_sc_hd__and3_4
X_16644_ _16676_/A _23698_/Q VGND VGND VPWR VPWR _16644_/X sky130_fd_sc_hd__or2_4
XFILLER_63_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12807_ _13400_/A _12799_/X _12807_/C VGND VGND VPWR VPWR _12807_/X sky130_fd_sc_hd__and3_4
XANTENNA__11552__B IRQ[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19363_ _19362_/X _18496_/X _19362_/X _24257_/Q VGND VGND VPWR VPWR _24257_/D sky130_fd_sc_hd__a2bb2o_4
X_16575_ _16539_/X _24082_/Q VGND VGND VPWR VPWR _16576_/C sky130_fd_sc_hd__or2_4
X_13787_ _14991_/A VGND VGND VPWR VPWR _13788_/A sky130_fd_sc_hd__buf_2
XFILLER_163_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22511__A2 _22508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18314_ _18314_/A _18311_/Y _18312_/Y _18313_/X VGND VGND VPWR VPWR _18315_/A sky130_fd_sc_hd__or4_4
X_12738_ _12738_/A _12735_/X _12738_/C VGND VGND VPWR VPWR _12738_/X sky130_fd_sc_hd__and3_4
X_15526_ _12258_/A _23745_/Q VGND VGND VPWR VPWR _15527_/C sky130_fd_sc_hd__or2_4
X_19294_ _24290_/Q _19295_/A _19293_/Y VGND VGND VPWR VPWR _24290_/D sky130_fd_sc_hd__o21a_4
XFILLER_128_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21042__A _21042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15457_ _15457_/A VGND VGND VPWR VPWR _15477_/A sky130_fd_sc_hd__buf_2
X_18245_ _18145_/X _18243_/X _20027_/A _18244_/X VGND VGND VPWR VPWR _24490_/D sky130_fd_sc_hd__a2bb2o_4
X_12669_ _12943_/A _12669_/B VGND VGND VPWR VPWR _12669_/X sky130_fd_sc_hd__or2_4
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ _13743_/A _14406_/X _14407_/X VGND VGND VPWR VPWR _14408_/X sky130_fd_sc_hd__and3_4
XANTENNA__21078__A2 _21073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18176_ _18176_/A VGND VGND VPWR VPWR _18176_/X sky130_fd_sc_hd__buf_2
X_15388_ _14705_/X _14848_/Y _15386_/X _14704_/X _15387_/X VGND VGND VPWR VPWR _15388_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__12383__B _23980_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11566__A2 IRQ[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17127_ _12061_/A VGND VGND VPWR VPWR _17128_/A sky130_fd_sc_hd__buf_2
X_14339_ _14517_/A _14339_/B VGND VGND VPWR VPWR _14340_/C sky130_fd_sc_hd__or2_4
XFILLER_144_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18494__A3 _18490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17058_ _17017_/B VGND VGND VPWR VPWR _17090_/A sky130_fd_sc_hd__inv_2
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22027__B2 _22021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16009_ _13443_/A VGND VGND VPWR VPWR _16009_/X sky130_fd_sc_hd__buf_2
XANTENNA__13495__A _12949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20589__A1 _18325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_HCLK clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__21786__B1 _15837_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21250__A2 _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22601__A _22608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20971_ _20344_/A _20970_/X _11514_/A _20269_/A VGND VGND VPWR VPWR _20971_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12839__A _13563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22710_ _20575_/A _22708_/X _13109_/B _22705_/X VGND VGND VPWR VPWR _23112_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11743__A _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15215__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19910__A _23083_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23690_ _23723_/CLK _21726_/X VGND VGND VPWR VPWR _23690_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22641_ _22648_/A VGND VGND VPWR VPWR _22641_/X sky130_fd_sc_hd__buf_2
XANTENNA__22502__A2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24023__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15869__B _15869_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22572_ _22539_/A VGND VGND VPWR VPWR _22572_/X sky130_fd_sc_hd__buf_2
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24311_ _24287_/CLK _19220_/X HRESETn VGND VGND VPWR VPWR _24311_/Q sky130_fd_sc_hd__dfrtp_4
X_21523_ _21523_/A VGND VGND VPWR VPWR _21549_/A sky130_fd_sc_hd__inv_2
XFILLER_22_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17390__B1 _17028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21069__A2 _21066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24242_ _24240_/CLK _19390_/X HRESETn VGND VGND VPWR VPWR _24242_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22266__B2 _22262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21454_ _21290_/X _21448_/X _23840_/Q _21452_/X VGND VGND VPWR VPWR _23840_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20791__A _20264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24173__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11557__A2 IRQ[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20405_ _20273_/A _20404_/Y _19252_/A _20323_/X VGND VGND VPWR VPWR _20405_/X sky130_fd_sc_hd__o22a_4
XFILLER_162_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19357__A _19324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24173_ _23383_/CLK _19934_/X HRESETn VGND VGND VPWR VPWR _24173_/Q sky130_fd_sc_hd__dfrtp_4
X_21385_ _21256_/X _21384_/X _16010_/B _21381_/X VGND VGND VPWR VPWR _21385_/X sky130_fd_sc_hd__o22a_4
XFILLER_162_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23124_ _23764_/CLK _23124_/D VGND VGND VPWR VPWR _23124_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22018__B2 _22014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20336_ _20336_/A VGND VGND VPWR VPWR _21528_/A sky130_fd_sc_hd__buf_2
XFILLER_162_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11918__A _11917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23055_ _18062_/X _23055_/B VGND VGND VPWR VPWR _23056_/C sky130_fd_sc_hd__or2_4
X_20267_ _18889_/B _20095_/X VGND VGND VPWR VPWR _20267_/X sky130_fd_sc_hd__or2_4
XFILLER_115_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22006_ _21831_/X _22003_/X _23532_/Q _22000_/X VGND VGND VPWR VPWR _23532_/D sky130_fd_sc_hd__o22a_4
XFILLER_163_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20198_ _20150_/A _20197_/X VGND VGND VPWR VPWR _20198_/X sky130_fd_sc_hd__or2_4
XFILLER_89_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11971_ _13453_/A VGND VGND VPWR VPWR _11971_/X sky130_fd_sc_hd__buf_2
X_23957_ _23617_/CLK _23957_/D VGND VGND VPWR VPWR _23957_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12749__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20031__A _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13710_ _13710_/A VGND VGND VPWR VPWR _15486_/A sky130_fd_sc_hd__buf_2
XFILLER_16_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22908_ _22908_/A VGND VGND VPWR VPWR _22908_/X sky130_fd_sc_hd__buf_2
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14690_ _15616_/A _14685_/X _14690_/C VGND VGND VPWR VPWR _14698_/B sky130_fd_sc_hd__or3_4
X_23888_ _23728_/CLK _21382_/X VGND VGND VPWR VPWR _16446_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13641_ _12186_/A _13641_/B _13641_/C VGND VGND VPWR VPWR _13641_/X sky130_fd_sc_hd__or3_4
X_22839_ _22845_/A _22839_/B VGND VGND VPWR VPWR HWDATA[13] sky130_fd_sc_hd__nor2_4
XFILLER_71_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14964__A _15369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16360_ _13407_/A _16356_/X _16359_/X VGND VGND VPWR VPWR _16360_/X sky130_fd_sc_hd__or3_4
XANTENNA__17340__A _15118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _13582_/A _13570_/Y _13581_/A VGND VGND VPWR VPWR _13573_/B sky130_fd_sc_hd__o21ai_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15311_ _13853_/A _15310_/X VGND VGND VPWR VPWR _15311_/X sky130_fd_sc_hd__and2_4
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _12881_/A _12523_/B _12523_/C VGND VGND VPWR VPWR _12524_/B sky130_fd_sc_hd__or3_4
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16291_ _15952_/A _16289_/X _16290_/X VGND VGND VPWR VPWR _16291_/X sky130_fd_sc_hd__and3_4
XANTENNA__12484__A _12484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18030_ _18022_/X _17964_/B _18025_/Y _18027_/X _23054_/B VGND VGND VPWR VPWR _18030_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_9_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15242_ _14200_/A _15170_/B VGND VGND VPWR VPWR _15243_/C sky130_fd_sc_hd__or2_4
X_12454_ _12454_/A VGND VGND VPWR VPWR _12455_/A sky130_fd_sc_hd__buf_2
XANTENNA__22257__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11548__A2 IRQ[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15795__A _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15173_ _12484_/A _15173_/B VGND VGND VPWR VPWR _15174_/C sky130_fd_sc_hd__or2_4
XFILLER_153_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12385_ _12407_/A _23628_/Q VGND VGND VPWR VPWR _12387_/B sky130_fd_sc_hd__or2_4
XFILLER_138_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14124_ _13981_/A VGND VGND VPWR VPWR _15281_/A sky130_fd_sc_hd__buf_2
XANTENNA__22009__B2 _22007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21480__A2 _21478_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19981_ _18670_/X _19328_/Y _19956_/X _19980_/X VGND VGND VPWR VPWR _19981_/X sky130_fd_sc_hd__o22a_4
XFILLER_125_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18932_ _13945_/X _18927_/X _19090_/A _18928_/X VGND VGND VPWR VPWR _24381_/D sky130_fd_sc_hd__o22a_4
X_14055_ _14075_/A _23616_/Q VGND VGND VPWR VPWR _14055_/X sky130_fd_sc_hd__or2_4
XFILLER_106_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13006_ _12513_/A _13006_/B VGND VGND VPWR VPWR _13007_/C sky130_fd_sc_hd__or2_4
XANTENNA__21232__A2 _21198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11547__B IRQ[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15019__B _23605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18863_ _18838_/X VGND VGND VPWR VPWR _18863_/X sky130_fd_sc_hd__buf_2
XFILLER_79_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22421__A _22421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17814_ _17836_/A VGND VGND VPWR VPWR _17814_/X sky130_fd_sc_hd__buf_2
XFILLER_95_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18794_ _17266_/X _18787_/X _24465_/Q _18790_/X VGND VGND VPWR VPWR _18794_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21037__A _21033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17745_ _17758_/A VGND VGND VPWR VPWR _17746_/A sky130_fd_sc_hd__inv_2
XFILLER_36_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14957_ _14783_/X _14953_/X _14956_/X VGND VGND VPWR VPWR _14957_/X sky130_fd_sc_hd__or3_4
XANTENNA__12659__A _12659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18936__A1 _14548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22732__A2 _22729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13908_ _13706_/A _13819_/B VGND VGND VPWR VPWR _13908_/X sky130_fd_sc_hd__or2_4
X_17676_ _17676_/A _17482_/X VGND VGND VPWR VPWR _17770_/A sky130_fd_sc_hd__or2_4
XFILLER_39_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14888_ _14881_/A _14959_/B VGND VGND VPWR VPWR _14888_/X sky130_fd_sc_hd__or2_4
XFILLER_62_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_15_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_30_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19415_ _19411_/X _18404_/X _19414_/X _24228_/Q VGND VGND VPWR VPWR _19415_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16627_ _16658_/A _16627_/B VGND VGND VPWR VPWR _16627_/X sky130_fd_sc_hd__or2_4
X_13839_ _12504_/A _13839_/B VGND VGND VPWR VPWR _13840_/C sky130_fd_sc_hd__or2_4
XFILLER_44_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19346_ _19343_/X _18184_/X _19343_/X _24268_/Q VGND VGND VPWR VPWR _24268_/D sky130_fd_sc_hd__a2bb2o_4
X_16558_ _16558_/A _23346_/Q VGND VGND VPWR VPWR _16560_/B sky130_fd_sc_hd__or2_4
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22496__B2 _22491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24196__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15509_ _15502_/A _15509_/B VGND VGND VPWR VPWR _15509_/X sky130_fd_sc_hd__or2_4
X_19277_ _19248_/B VGND VGND VPWR VPWR _19277_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19900__A3 _19899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16489_ _13383_/A _16471_/X _16489_/C VGND VGND VPWR VPWR _16489_/X sky130_fd_sc_hd__or3_4
XFILLER_31_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18228_ _17873_/X _18227_/X _17848_/A _18052_/X VGND VGND VPWR VPWR _18229_/A sky130_fd_sc_hd__o22a_4
XFILLER_164_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18159_ _17933_/X _17989_/X _17824_/X _17993_/X VGND VGND VPWR VPWR _18159_/X sky130_fd_sc_hd__o22a_4
XFILLER_156_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21170_ _20801_/X _21169_/X _23999_/Q _21166_/X VGND VGND VPWR VPWR _23999_/D sky130_fd_sc_hd__o22a_4
XFILLER_117_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13937__B _24093_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20121_ _11570_/B VGND VGND VPWR VPWR _20121_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14114__A _14114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20052_ _18398_/X _20031_/X _20051_/Y _20042_/X VGND VGND VPWR VPWR _20052_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13953__A _13953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17425__A _14263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23811_ _23656_/CLK _23811_/D VGND VGND VPWR VPWR _15841_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13672__B _13761_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12569__A _12569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22723__A2 _22722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23742_ _23678_/CLK _21643_/X VGND VGND VPWR VPWR _13713_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20954_ _24248_/Q VGND VGND VPWR VPWR _20954_/Y sky130_fd_sc_hd__inv_2
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23413__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23673_ _23391_/CLK _21750_/X VGND VGND VPWR VPWR _14720_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _18643_/X _20675_/X _20780_/X _20884_/Y VGND VGND VPWR VPWR _20885_/X sky130_fd_sc_hd__a211o_4
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22624_ _22464_/X _22622_/X _13736_/B _22619_/X VGND VGND VPWR VPWR _22624_/X sky130_fd_sc_hd__o22a_4
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24379__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22555_ _22555_/A VGND VGND VPWR VPWR _22555_/X sky130_fd_sc_hd__buf_2
XANTENNA__22239__A1 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21506_ _21506_/A VGND VGND VPWR VPWR _21506_/X sky130_fd_sc_hd__buf_2
XANTENNA__22239__B2 _22234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22486_ _11845_/B VGND VGND VPWR VPWR _22486_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_35_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_35_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14008__B _23712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24225_ _24137_/CLK _24225_/D HRESETn VGND VGND VPWR VPWR _24225_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21437_ _21261_/X _21434_/X _12390_/B _21431_/X VGND VGND VPWR VPWR _23852_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16504__A _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24156_ _24495_/CLK _20011_/Y HRESETn VGND VGND VPWR VPWR _17669_/A sky130_fd_sc_hd__dfrtp_4
X_12170_ _12151_/A _23507_/Q VGND VGND VPWR VPWR _12172_/B sky130_fd_sc_hd__or2_4
XFILLER_163_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21368_ _21315_/X _21341_/A _23893_/Q _21331_/A VGND VGND VPWR VPWR _23893_/D sky130_fd_sc_hd__o22a_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23107_ _23523_/CLK _22717_/X VGND VGND VPWR VPWR _15840_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_123_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11648__A _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20319_ _24467_/Q VGND VGND VPWR VPWR _20320_/A sky130_fd_sc_hd__inv_2
X_24087_ _23544_/CLK _24087_/D VGND VGND VPWR VPWR _15170_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14024__A _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21299_ _20860_/A VGND VGND VPWR VPWR _21299_/X sky130_fd_sc_hd__buf_2
XANTENNA__21214__A2 _21212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23038_ _23043_/A _23038_/B VGND VGND VPWR VPWR _23038_/Y sky130_fd_sc_hd__nand2_4
XFILLER_118_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22411__B2 _22409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22241__A _22226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18091__A1 _17875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15860_ _13539_/A _15799_/B VGND VGND VPWR VPWR _15862_/B sky130_fd_sc_hd__or2_4
XFILLER_49_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14811_ _11674_/A _14794_/X _14811_/C VGND VGND VPWR VPWR _14811_/X sky130_fd_sc_hd__or3_4
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12479__A _12878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15791_ _12741_/A _15789_/X _15790_/X VGND VGND VPWR VPWR _15791_/X sky130_fd_sc_hd__and3_4
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18918__A1 _13262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22714__A2 _22708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17530_ _13567_/X _17530_/B VGND VGND VPWR VPWR _17530_/Y sky130_fd_sc_hd__nand2_4
XFILLER_123_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14742_ _11932_/A _14738_/X _14742_/C VGND VGND VPWR VPWR _14742_/X sky130_fd_sc_hd__or3_4
X_11954_ _11905_/X VGND VGND VPWR VPWR _12012_/A sky130_fd_sc_hd__buf_2
XANTENNA__23093__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23072__A _23071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17461_ _17459_/Y _17460_/X VGND VGND VPWR VPWR _17461_/X sky130_fd_sc_hd__or2_4
X_14673_ _14235_/A VGND VGND VPWR VPWR _14674_/A sky130_fd_sc_hd__buf_2
X_11885_ _16116_/A VGND VGND VPWR VPWR _16595_/A sky130_fd_sc_hd__buf_2
XFILLER_60_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14694__A _14657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19200_ _24321_/Q _19142_/B _19199_/Y VGND VGND VPWR VPWR _24321_/D sky130_fd_sc_hd__o21a_4
X_16412_ _16401_/X _16412_/B VGND VGND VPWR VPWR _16412_/X sky130_fd_sc_hd__or2_4
X_13624_ _12504_/A _13624_/B VGND VGND VPWR VPWR _13624_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_117_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR _23675_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17392_ _17391_/X VGND VGND VPWR VPWR _17394_/A sky130_fd_sc_hd__inv_2
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19131_ _24310_/Q _19131_/B VGND VGND VPWR VPWR _19131_/X sky130_fd_sc_hd__and2_4
X_13555_ _12773_/X _13555_/B _13555_/C VGND VGND VPWR VPWR _13556_/C sky130_fd_sc_hd__and3_4
X_16343_ _16465_/A _16341_/X _16343_/C VGND VGND VPWR VPWR _16343_/X sky130_fd_sc_hd__and3_4
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21150__B2 _21145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12506_ _12506_/A VGND VGND VPWR VPWR _12872_/A sky130_fd_sc_hd__buf_2
XANTENNA__13103__A _13103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16274_ _16099_/X _16274_/B VGND VGND VPWR VPWR _16274_/X sky130_fd_sc_hd__or2_4
X_19062_ _19052_/X _19061_/X _19052_/X _11528_/A VGND VGND VPWR VPWR _24354_/D sky130_fd_sc_hd__a2bb2o_4
X_13486_ _12659_/A VGND VGND VPWR VPWR _13528_/A sky130_fd_sc_hd__buf_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22416__A _20360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18013_ _17673_/X _18013_/B _18013_/C VGND VGND VPWR VPWR _18014_/B sky130_fd_sc_hd__or3_4
X_15225_ _14630_/A _15225_/B _15225_/C VGND VGND VPWR VPWR _15233_/B sky130_fd_sc_hd__or3_4
X_12437_ _12847_/A _12579_/B VGND VGND VPWR VPWR _12437_/X sky130_fd_sc_hd__or2_4
XANTENNA__12942__A _12942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16414__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15156_ _14148_/A _15156_/B VGND VGND VPWR VPWR _15157_/C sky130_fd_sc_hd__or2_4
X_12368_ _13251_/A VGND VGND VPWR VPWR _15894_/A sky130_fd_sc_hd__buf_2
XANTENNA__21453__A2 _21448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22650__B2 _22648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12661__B _12564_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14107_ _12287_/A _14107_/B _14107_/C VGND VGND VPWR VPWR _14107_/X sky130_fd_sc_hd__or3_4
XFILLER_5_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19964_ _18407_/A _19964_/B VGND VGND VPWR VPWR _19966_/C sky130_fd_sc_hd__nor2_4
X_15087_ _14073_/A _15085_/X _15087_/C VGND VGND VPWR VPWR _15087_/X sky130_fd_sc_hd__and3_4
X_12299_ _12299_/A VGND VGND VPWR VPWR _12300_/A sky130_fd_sc_hd__buf_2
XFILLER_99_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18915_ _17156_/A _18913_/X _24394_/Q _18914_/X VGND VGND VPWR VPWR _24394_/D sky130_fd_sc_hd__o22a_4
X_14038_ _11660_/A _23168_/Q VGND VGND VPWR VPWR _14038_/X sky130_fd_sc_hd__or2_4
XFILLER_136_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22402__B2 _22366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19895_ _19895_/A _19742_/A _19895_/C _19894_/X VGND VGND VPWR VPWR _19895_/X sky130_fd_sc_hd__or4_4
XANTENNA__22151__A _20840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14869__A _14114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13773__A _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18846_ _17255_/X _18840_/X _24434_/Q _18843_/X VGND VGND VPWR VPWR _24434_/D sky130_fd_sc_hd__o22a_4
XFILLER_171_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18777_ _16935_/A _18775_/X _17652_/X _18776_/Y VGND VGND VPWR VPWR _18777_/X sky130_fd_sc_hd__o22a_4
X_15989_ _15960_/A _15989_/B VGND VGND VPWR VPWR _15990_/C sky130_fd_sc_hd__or2_4
XANTENNA__18909__A1 _17139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17728_ _17730_/B _17727_/X VGND VGND VPWR VPWR _17762_/B sky130_fd_sc_hd__or2_4
X_17659_ _17659_/A _17659_/B VGND VGND VPWR VPWR _17659_/X sky130_fd_sc_hd__and2_4
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20670_ _20670_/A VGND VGND VPWR VPWR _20671_/A sky130_fd_sc_hd__buf_2
XFILLER_143_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19329_ _17037_/Y _19328_/A _17048_/A _19328_/Y VGND VGND VPWR VPWR _19330_/A sky130_fd_sc_hd__o22a_4
X_22340_ _23330_/Q VGND VGND VPWR VPWR _22340_/X sky130_fd_sc_hd__buf_2
XFILLER_109_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21692__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13948__A _13863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22271_ _22169_/X _22244_/A _23381_/Q _22226_/X VGND VGND VPWR VPWR _23381_/D sky130_fd_sc_hd__o22a_4
XFILLER_145_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24010_ _23558_/CLK _24010_/D VGND VGND VPWR VPWR _24010_/Q sky130_fd_sc_hd__dfxtp_4
X_21222_ _20841_/X _21219_/X _23965_/Q _21216_/X VGND VGND VPWR VPWR _23965_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21444__A2 _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21153_ _20509_/X _21148_/X _12632_/B _21152_/X VGND VGND VPWR VPWR _21153_/X sky130_fd_sc_hd__o22a_4
XFILLER_160_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24211__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20104_ _20124_/B _20093_/X _20098_/X _11640_/B VGND VGND VPWR VPWR _20104_/X sky130_fd_sc_hd__or4_4
XFILLER_104_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21084_ _21083_/X VGND VGND VPWR VPWR _21118_/A sky130_fd_sc_hd__buf_2
XFILLER_150_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13683__A _15447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20035_ _20034_/X VGND VGND VPWR VPWR _20035_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17155__A _12842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20955__A1 _20305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22996__A _18394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20955__B2 _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12299__A _12299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21986_ _21883_/X _21981_/X _14946_/B _21950_/A VGND VGND VPWR VPWR _23542_/D sky130_fd_sc_hd__o22a_4
XFILLER_73_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23725_ _23501_/CLK _21672_/X VGND VGND VPWR VPWR _16226_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21405__A _21405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20937_ _20937_/A VGND VGND VPWR VPWR _20938_/A sky130_fd_sc_hd__buf_2
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20183__A2 IRQ[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21380__B2 _21374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15403__A _13656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _13566_/A VGND VGND VPWR VPWR _13417_/A sky130_fd_sc_hd__buf_2
X_23656_ _23656_/CLK _23656_/D VGND VGND VPWR VPWR _23656_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20868_ _20871_/A _20865_/A VGND VGND VPWR VPWR _20869_/A sky130_fd_sc_hd__and2_4
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22607_ _22435_/X _22601_/X _12794_/B _22605_/X VGND VGND VPWR VPWR _23178_/D sky130_fd_sc_hd__o22a_4
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15122__B _15122_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23587_ _23587_/CLK _21918_/X VGND VGND VPWR VPWR _15866_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17336__B1 _21081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20799_ _24223_/Q _20773_/X _20798_/X VGND VGND VPWR VPWR _22461_/A sky130_fd_sc_hd__o21a_4
XANTENNA__14019__A _13877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13340_ _13453_/A _13315_/X _13322_/X _13331_/X _13339_/X VGND VGND VPWR VPWR _13340_/X
+ sky130_fd_sc_hd__a32o_4
X_22538_ _22537_/X VGND VGND VPWR VPWR _22539_/A sky130_fd_sc_hd__buf_2
XANTENNA__21683__A2 _21677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21140__A _21136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13271_ _13192_/X _13270_/X _13265_/Y VGND VGND VPWR VPWR _13271_/X sky130_fd_sc_hd__a21o_4
XANTENNA__13858__A _15447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12762__A _12762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22469_ _22433_/A VGND VGND VPWR VPWR _22469_/X sky130_fd_sc_hd__buf_2
XANTENNA__16234__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15010_ _13974_/A _23157_/Q VGND VGND VPWR VPWR _15010_/X sky130_fd_sc_hd__or2_4
X_12222_ _12269_/A VGND VGND VPWR VPWR _12721_/A sky130_fd_sc_hd__buf_2
X_24208_ _24184_/CLK _19608_/X HRESETn VGND VGND VPWR VPWR _17398_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21435__A2 _21434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22632__B2 _22626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18300__A2 _18278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12153_ _12129_/A _12151_/X _12152_/X VGND VGND VPWR VPWR _12153_/X sky130_fd_sc_hd__and3_4
X_24139_ _24137_/CLK _20091_/Y HRESETn VGND VGND VPWR VPWR _16967_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16961_ _24145_/Q VGND VGND VPWR VPWR _16983_/A sky130_fd_sc_hd__inv_2
X_12084_ _16725_/A _12084_/B _12083_/X VGND VGND VPWR VPWR _12085_/C sky130_fd_sc_hd__and3_4
XFILLER_89_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21199__B2 _21195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18700_ _16939_/X _18697_/Y _16940_/Y _18699_/X VGND VGND VPWR VPWR _18700_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13593__A _13593_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15912_ _13566_/A _15912_/B _15912_/C VGND VGND VPWR VPWR _15912_/X sky130_fd_sc_hd__and3_4
XANTENNA__17065__A _17100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19680_ _19680_/A VGND VGND VPWR VPWR _19683_/A sky130_fd_sc_hd__inv_2
X_16892_ _12846_/X _16891_/X _12846_/X _16891_/X VGND VGND VPWR VPWR _16895_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18631_ _18627_/X _18630_/X _17741_/A VGND VGND VPWR VPWR _18632_/A sky130_fd_sc_hd__or3_4
X_15843_ _12905_/A _15843_/B VGND VGND VPWR VPWR _15845_/B sky130_fd_sc_hd__or2_4
XANTENNA__22148__B1 _23455_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18562_ _18562_/A _18202_/Y VGND VGND VPWR VPWR _18562_/X sky130_fd_sc_hd__and2_4
XANTENNA__22699__B2 _22698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15774_ _15741_/X _15701_/B VGND VGND VPWR VPWR _15774_/X sky130_fd_sc_hd__or2_4
XANTENNA__12002__A _12105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12986_ _12846_/X _12986_/B VGND VGND VPWR VPWR _12986_/X sky130_fd_sc_hd__or2_4
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17513_ _17165_/Y _17515_/B VGND VGND VPWR VPWR _17513_/X sky130_fd_sc_hd__or2_4
X_14725_ _11913_/A _14723_/X _14725_/C VGND VGND VPWR VPWR _14726_/C sky130_fd_sc_hd__and3_4
X_11937_ _15978_/A VGND VGND VPWR VPWR _16129_/A sky130_fd_sc_hd__buf_2
X_18493_ _17396_/A _18491_/X _18008_/A VGND VGND VPWR VPWR _18493_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12937__A _12975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17444_ _17437_/A _17443_/X VGND VGND VPWR VPWR _17444_/Y sky130_fd_sc_hd__nor2_4
X_14656_ _14656_/A VGND VGND VPWR VPWR _14680_/A sky130_fd_sc_hd__buf_2
X_11868_ _11867_/X VGND VGND VPWR VPWR _11868_/X sky130_fd_sc_hd__buf_2
XFILLER_60_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13607_ _13607_/A VGND VGND VPWR VPWR _13823_/A sky130_fd_sc_hd__buf_2
XANTENNA__11560__B IRQ[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17375_ _17375_/A _17375_/B VGND VGND VPWR VPWR _18415_/B sky130_fd_sc_hd__or2_4
XANTENNA__21123__B2 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11799_ _11704_/X VGND VGND VPWR VPWR _12129_/A sky130_fd_sc_hd__buf_2
XFILLER_14_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14587_ _13601_/A _14587_/B VGND VGND VPWR VPWR _14587_/X sky130_fd_sc_hd__or2_4
XFILLER_41_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19114_ _11518_/A VGND VGND VPWR VPWR _19114_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24362__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16326_ _16313_/A _16324_/X _16325_/X VGND VGND VPWR VPWR _16326_/X sky130_fd_sc_hd__and3_4
XFILLER_174_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13538_ _12955_/A VGND VGND VPWR VPWR _13539_/A sky130_fd_sc_hd__buf_2
XFILLER_174_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22146__A _22461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13768__A _12623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19045_ _19038_/X _19044_/X _19038_/X _24357_/Q VGND VGND VPWR VPWR _19045_/X sky130_fd_sc_hd__a2bb2o_4
X_13469_ _13441_/A _13469_/B VGND VGND VPWR VPWR _13471_/B sky130_fd_sc_hd__or2_4
X_16257_ _16157_/A _16257_/B VGND VGND VPWR VPWR _16257_/X sky130_fd_sc_hd__or2_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24234__CLK _24271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15208_ _14635_/A _15208_/B _15207_/X VGND VGND VPWR VPWR _15209_/C sky130_fd_sc_hd__and3_4
XFILLER_173_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16188_ _16215_/A _23949_/Q VGND VGND VPWR VPWR _16190_/B sky130_fd_sc_hd__or2_4
XANTENNA__22623__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15139_ _14267_/A _15139_/B VGND VGND VPWR VPWR _15141_/B sky130_fd_sc_hd__or2_4
XFILLER_173_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19947_ _22908_/A VGND VGND VPWR VPWR _19953_/A sky130_fd_sc_hd__buf_2
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19878_ _19834_/A _19578_/Y _19601_/B _19877_/X VGND VGND VPWR VPWR _19878_/X sky130_fd_sc_hd__a211o_4
XFILLER_67_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18829_ _15380_/A _18824_/X _24440_/Q _18825_/X VGND VGND VPWR VPWR _18829_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14111__B _23999_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21840_ _21838_/X _21839_/X _23625_/Q _21834_/X VGND VGND VPWR VPWR _21840_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13008__A _12911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21771_ _21541_/X _21770_/X _23662_/Q _21767_/X VGND VGND VPWR VPWR _23662_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12847__A _12847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23510_ _23511_/CLK _23510_/D VGND VGND VPWR VPWR _14850_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20722_ _20364_/B _20671_/A VGND VGND VPWR VPWR _20722_/X sky130_fd_sc_hd__or2_4
X_24490_ _24277_/CLK _24490_/D HRESETn VGND VGND VPWR VPWR _20027_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23441_ _23409_/CLK _23441_/D VGND VGND VPWR VPWR _16799_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_149_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20653_ _18426_/X _20469_/X _20514_/X _20652_/Y VGND VGND VPWR VPWR _20653_/X sky130_fd_sc_hd__a211o_4
XFILLER_17_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_100_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR _23649_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21114__B2 _21108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23372_ _23852_/CLK _22290_/X VGND VGND VPWR VPWR _12204_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21665__A2 _21663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20584_ _20270_/X VGND VGND VPWR VPWR _20584_/X sky130_fd_sc_hd__buf_2
XFILLER_139_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13678__A _15439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22323_ _12142_/B VGND VGND VPWR VPWR _23347_/D sky130_fd_sc_hd__buf_2
X_22254_ _22139_/X _22251_/X _15432_/B _22248_/X VGND VGND VPWR VPWR _23394_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21895__A _21909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21417__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22614__B2 _22612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23601__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21205_ _21198_/A VGND VGND VPWR VPWR _21205_/X sky130_fd_sc_hd__buf_2
XFILLER_105_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22185_ _22105_/X _22180_/X _16432_/B _22184_/X VGND VGND VPWR VPWR _23440_/D sky130_fd_sc_hd__o22a_4
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19491__B1 HRDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21136_ _21136_/A VGND VGND VPWR VPWR _21152_/A sky130_fd_sc_hd__inv_2
XFILLER_28_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20304__A _20977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11926__A _16713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21067_ _20801_/X _21066_/X _24063_/Q _21063_/X VGND VGND VPWR VPWR _24063_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20389__C1 _20388_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14302__A _14302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23751__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21050__B1 _12647_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20018_ _19950_/X VGND VGND VPWR VPWR _20018_/X sky130_fd_sc_hd__buf_2
XFILLER_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11645__B _17060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12840_ _13415_/A _12832_/X _12840_/C VGND VGND VPWR VPWR _12840_/X sky130_fd_sc_hd__and3_4
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12771_ _13556_/A _12764_/X _12770_/X VGND VGND VPWR VPWR _12771_/X sky130_fd_sc_hd__or3_4
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ _21853_/X _21967_/X _15807_/B _21964_/X VGND VGND VPWR VPWR _23555_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12757__A _13067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11661__A _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21353__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _14510_/A _23323_/Q VGND VGND VPWR VPWR _14512_/B sky130_fd_sc_hd__or2_4
XANTENNA__15133__A _14169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11722_ _15606_/A VGND VGND VPWR VPWR _14658_/A sky130_fd_sc_hd__buf_2
X_15490_ _15502_/A _15490_/B VGND VGND VPWR VPWR _15491_/C sky130_fd_sc_hd__or2_4
X_23708_ _23675_/CLK _21696_/X VGND VGND VPWR VPWR _14399_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _13011_/A _14441_/B _14440_/X VGND VGND VPWR VPWR _14441_/X sky130_fd_sc_hd__and3_4
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11653_/A VGND VGND VPWR VPWR _11654_/A sky130_fd_sc_hd__buf_2
X_23639_ _23770_/CLK _23639_/D VGND VGND VPWR VPWR _15173_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21105__B2 _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24257__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14372_ _14372_/A _14368_/X _14372_/C VGND VGND VPWR VPWR _14373_/C sky130_fd_sc_hd__or3_4
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17160_ _17160_/A VGND VGND VPWR VPWR _17160_/X sky130_fd_sc_hd__buf_2
XFILLER_128_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11584_ _20124_/A _20125_/A _11583_/X VGND VGND VPWR VPWR _11585_/D sky130_fd_sc_hd__or3_4
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16111_ _16138_/A _16107_/X _16111_/C VGND VGND VPWR VPWR _16111_/X sky130_fd_sc_hd__or3_4
X_13323_ _12866_/A VGND VGND VPWR VPWR _13475_/A sky130_fd_sc_hd__buf_2
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13588__A _15029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12492__A _12492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17091_ _17091_/A _17090_/A _17077_/A VGND VGND VPWR VPWR _17091_/X sky130_fd_sc_hd__and3_4
XFILLER_122_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16042_ _16049_/A _23470_/Q VGND VGND VPWR VPWR _16042_/X sky130_fd_sc_hd__or2_4
X_13254_ _12338_/X _13254_/B _13254_/C VGND VGND VPWR VPWR _13258_/B sky130_fd_sc_hd__and3_4
XFILLER_6_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18809__B1 _20157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21408__A2 _21405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23281__CLK _23281_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16899__A _16899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12205_ _12512_/A VGND VGND VPWR VPWR _12687_/A sky130_fd_sc_hd__buf_2
XFILLER_170_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13185_ _12301_/A _13185_/B _13184_/X VGND VGND VPWR VPWR _13189_/B sky130_fd_sc_hd__and3_4
XFILLER_135_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19801_ _19683_/A _19800_/X _19613_/X _19811_/B VGND VGND VPWR VPWR _19801_/X sky130_fd_sc_hd__a2bb2o_4
X_12136_ _12167_/A _12136_/B VGND VGND VPWR VPWR _12136_/X sky130_fd_sc_hd__or2_4
XFILLER_124_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17993_ _17922_/X _17858_/X _17945_/X _17860_/X VGND VGND VPWR VPWR _17993_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11836__A _11836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19732_ _19439_/A VGND VGND VPWR VPWR _19732_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16944_ _24161_/Q VGND VGND VPWR VPWR _16945_/A sky130_fd_sc_hd__inv_2
XANTENNA__15308__A _15017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12067_ _16710_/A _12067_/B _12066_/X VGND VGND VPWR VPWR _12067_/X sky130_fd_sc_hd__or3_4
XANTENNA__14212__A _14635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19785__A1 _20598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19663_ _19690_/B VGND VGND VPWR VPWR _19663_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16875_ _15388_/X _14552_/Y _15389_/B VGND VGND VPWR VPWR _16875_/X sky130_fd_sc_hd__o21a_4
X_18614_ _18613_/X VGND VGND VPWR VPWR _18614_/Y sky130_fd_sc_hd__inv_2
X_15826_ _12884_/A _15826_/B VGND VGND VPWR VPWR _15826_/X sky130_fd_sc_hd__or2_4
X_19594_ _19528_/A _19479_/A _19524_/A VGND VGND VPWR VPWR _19681_/B sky130_fd_sc_hd__or3_4
XANTENNA__21045__A _21045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18545_ _18545_/A _17434_/A VGND VGND VPWR VPWR _18545_/X sky130_fd_sc_hd__and2_4
XFILLER_79_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15757_ _12778_/X _15755_/X _15756_/X VGND VGND VPWR VPWR _15757_/X sky130_fd_sc_hd__and3_4
XANTENNA__19363__A2_N _18496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12969_ _12945_/A _12965_/X _12968_/X VGND VGND VPWR VPWR _12977_/B sky130_fd_sc_hd__or3_4
XANTENNA__12667__A _12945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21344__B2 _21338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15043__A _13662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14708_ _13791_/A _14706_/X _14708_/C VGND VGND VPWR VPWR _14708_/X sky130_fd_sc_hd__and3_4
X_18476_ _18453_/X _18475_/X _24482_/Q _18453_/X VGND VGND VPWR VPWR _24482_/D sky130_fd_sc_hd__a2bb2o_4
X_15688_ _12721_/A _15688_/B VGND VGND VPWR VPWR _15689_/C sky130_fd_sc_hd__or2_4
XANTENNA__20552__C1 _20551_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12386__B _24076_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17427_ _17427_/A _17280_/B VGND VGND VPWR VPWR _17427_/X sky130_fd_sc_hd__or2_4
X_14639_ _14684_/A _14564_/B VGND VGND VPWR VPWR _14639_/X sky130_fd_sc_hd__or2_4
XFILLER_14_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21647__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22844__A1 _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17358_ _17342_/Y _17358_/B VGND VGND VPWR VPWR _17358_/Y sky130_fd_sc_hd__nor2_4
XFILLER_158_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16309_ _11858_/A _11631_/X _16278_/X _11608_/A _16308_/X VGND VGND VPWR VPWR _16309_/X
+ sky130_fd_sc_hd__a32o_4
X_17289_ _14701_/Y _17292_/B VGND VGND VPWR VPWR _17289_/X sky130_fd_sc_hd__or2_4
XFILLER_174_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19028_ _19024_/X _19027_/X _19024_/X _24360_/Q VGND VGND VPWR VPWR _24360_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22072__A2 _22067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11746__A _16080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15218__A _11673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23990_ _23991_/CLK _23990_/D VGND VGND VPWR VPWR _23990_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_25_0_HCLK clkbuf_6_12_0_HCLK/X VGND VGND VPWR VPWR _24306_/CLK sky130_fd_sc_hd__clkbuf_1
X_22941_ _22940_/X VGND VGND VPWR VPWR HADDR[6] sky130_fd_sc_hd__inv_2
Xclkbuf_7_88_0_HCLK clkbuf_7_89_0_HCLK/A VGND VGND VPWR VPWR _23391_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21583__B2 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22872_ _17273_/Y _22800_/Y _22815_/X VGND VGND VPWR VPWR _22872_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18248__B _17906_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21823_ _21821_/X _21815_/X _16424_/B _21822_/X VGND VGND VPWR VPWR _23632_/D sky130_fd_sc_hd__o22a_4
XFILLER_58_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12577__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16049__A _16049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21335__B2 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23154__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21754_ _21600_/X _21727_/A _23669_/Q _21717_/A VGND VGND VPWR VPWR _23669_/D sky130_fd_sc_hd__o22a_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21886__A2 _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20705_ _24418_/Q _20645_/X _20161_/A _20704_/X VGND VGND VPWR VPWR _20705_/X sky130_fd_sc_hd__o22a_4
XFILLER_145_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24473_ _24471_/CLK _18686_/X HRESETn VGND VGND VPWR VPWR _24473_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21685_ _21565_/X _21684_/X _23716_/Q _21681_/X VGND VGND VPWR VPWR _23716_/D sky130_fd_sc_hd__o22a_4
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23424_ _23744_/CLK _23424_/D VGND VGND VPWR VPWR _23424_/Q sky130_fd_sc_hd__dfxtp_4
X_20636_ _20895_/A VGND VGND VPWR VPWR _20636_/X sky130_fd_sc_hd__buf_2
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15400__B _23778_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23355_ _23772_/CLK _22314_/X VGND VGND VPWR VPWR _14487_/B sky130_fd_sc_hd__dfxtp_4
X_20567_ _20515_/X _20566_/X _19149_/A _20522_/X VGND VGND VPWR VPWR _20567_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22306_ _22141_/X _22301_/X _15525_/B _22305_/X VGND VGND VPWR VPWR _23361_/D sky130_fd_sc_hd__o22a_4
X_23286_ _23671_/CLK _23286_/D VGND VGND VPWR VPWR _14929_/B sky130_fd_sc_hd__dfxtp_4
X_20498_ _20490_/X _20497_/Y _24299_/Q _20323_/X VGND VGND VPWR VPWR _20498_/X sky130_fd_sc_hd__o22a_4
X_22237_ _22244_/A VGND VGND VPWR VPWR _22237_/X sky130_fd_sc_hd__buf_2
XANTENNA__22063__A2 _22060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22168_ _22167_/X _22159_/X _14875_/B _22106_/A VGND VGND VPWR VPWR _23446_/D sky130_fd_sc_hd__o22a_4
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21119_ _20801_/X _21118_/X _24031_/Q _21115_/X VGND VGND VPWR VPWR _24031_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15128__A _13788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11656__A _13923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19823__A _19823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22099_ _22123_/A VGND VGND VPWR VPWR _22099_/X sky130_fd_sc_hd__buf_2
X_14990_ _14171_/A _14990_/B _14990_/C VGND VGND VPWR VPWR _14991_/C sky130_fd_sc_hd__and3_4
XANTENNA__14032__A _13696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13941_ _13697_/A _13939_/X _13940_/X VGND VGND VPWR VPWR _13942_/C sky130_fd_sc_hd__and3_4
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21574__B2 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18439__A _18485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13871__A _13923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16660_ _16682_/A _16656_/X _16660_/C VGND VGND VPWR VPWR _16668_/B sky130_fd_sc_hd__or3_4
X_13872_ _13719_/A VGND VGND VPWR VPWR _14375_/A sky130_fd_sc_hd__buf_2
X_15611_ _15611_/A _24001_/Q VGND VGND VPWR VPWR _15612_/C sky130_fd_sc_hd__or2_4
X_12823_ _13400_/A _12815_/X _12822_/X VGND VGND VPWR VPWR _12823_/X sky130_fd_sc_hd__and3_4
XANTENNA__17062__B _17077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20129__A2 _20128_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16591_ _16556_/A _16589_/X _16591_/C VGND VGND VPWR VPWR _16592_/C sky130_fd_sc_hd__and3_4
XANTENNA__12487__A _12487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22523__B1 _23231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18330_ _16941_/X VGND VGND VPWR VPWR _18330_/X sky130_fd_sc_hd__buf_2
XANTENNA__24462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15542_ _12546_/A _15538_/X _15541_/X VGND VGND VPWR VPWR _15542_/X sky130_fd_sc_hd__or3_4
X_12754_ _12945_/A VGND VGND VPWR VPWR _13556_/A sky130_fd_sc_hd__buf_2
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11704_/X VGND VGND VPWR VPWR _11705_/X sky130_fd_sc_hd__buf_2
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18261_ _18261_/A VGND VGND VPWR VPWR _18261_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12685_ _13046_/A VGND VGND VPWR VPWR _13339_/A sky130_fd_sc_hd__buf_2
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ _13053_/A _15473_/B VGND VGND VPWR VPWR _15473_/X sky130_fd_sc_hd__or2_4
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _12680_/X _17197_/X _17153_/Y _17198_/X VGND VGND VPWR VPWR _17212_/X sky130_fd_sc_hd__o22a_4
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424_ _13687_/A VGND VGND VPWR VPWR _14431_/A sky130_fd_sc_hd__buf_2
X_11636_ _11636_/A VGND VGND VPWR VPWR _11636_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21629__A2 _21627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18192_ _18310_/A _17600_/D VGND VGND VPWR VPWR _18192_/X sky130_fd_sc_hd__or2_4
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17143_ _14413_/Y _17131_/X _16242_/X _17133_/X VGND VGND VPWR VPWR _17143_/X sky130_fd_sc_hd__o22a_4
XFILLER_156_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11567_ _11567_/A IRQ[10] VGND VGND VPWR VPWR _11567_/X sky130_fd_sc_hd__and2_4
X_14355_ _14367_/A _14355_/B VGND VGND VPWR VPWR _14355_/X sky130_fd_sc_hd__or2_4
XANTENNA__21031__C _21184_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14207__A _11654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13111__A _13103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23797__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13306_ _13306_/A _13302_/X _13306_/C VGND VGND VPWR VPWR _13306_/X sky130_fd_sc_hd__or3_4
XFILLER_6_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17074_ _17146_/A VGND VGND VPWR VPWR _17074_/X sky130_fd_sc_hd__buf_2
X_14286_ _13823_/A VGND VGND VPWR VPWR _15400_/A sky130_fd_sc_hd__buf_2
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16025_ _16066_/A _16025_/B _16024_/X VGND VGND VPWR VPWR _16026_/C sky130_fd_sc_hd__and3_4
X_13237_ _13220_/A _13237_/B VGND VGND VPWR VPWR _13237_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22054__A2 _22053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17518__A _13192_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12950__A _12950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16422__A _16009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13168_ _13164_/A _13237_/B VGND VGND VPWR VPWR _13170_/B sky130_fd_sc_hd__or2_4
XANTENNA__13765__B _13765_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12119_ _12127_/A _12119_/B VGND VGND VPWR VPWR _12119_/X sky130_fd_sc_hd__or2_4
XFILLER_170_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19733__A HRDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13099_ _13099_/A _13099_/B _13099_/C VGND VGND VPWR VPWR _13099_/X sky130_fd_sc_hd__and3_4
X_17976_ _17809_/A VGND VGND VPWR VPWR _17976_/X sky130_fd_sc_hd__buf_2
XFILLER_66_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19715_ _19563_/X _19691_/A _19647_/Y VGND VGND VPWR VPWR _19715_/X sky130_fd_sc_hd__a21o_4
X_16927_ _11593_/A VGND VGND VPWR VPWR _16927_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20598__B _20598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13781__A _15517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19646_ _19690_/B _19646_/B VGND VGND VPWR VPWR _19657_/B sky130_fd_sc_hd__nor2_4
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16858_ _16853_/X _16858_/B _16857_/X VGND VGND VPWR VPWR _16858_/X sky130_fd_sc_hd__and3_4
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15809_ _12874_/A _15805_/X _15809_/C VGND VGND VPWR VPWR _15809_/X sky130_fd_sc_hd__or3_4
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19577_ _20364_/B _19573_/X _19575_/X _19576_/X VGND VGND VPWR VPWR _19577_/X sky130_fd_sc_hd__a211o_4
XFILLER_20_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12397__A _11682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16789_ _16639_/A _23985_/Q VGND VGND VPWR VPWR _16790_/C sky130_fd_sc_hd__or2_4
X_18528_ _17762_/X _17724_/X _17723_/A VGND VGND VPWR VPWR _18528_/X sky130_fd_sc_hd__o21a_4
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21868__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20525__C1 _20524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24132__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21503__A _21489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18459_ _18406_/A _17446_/B VGND VGND VPWR VPWR _18459_/X sky130_fd_sc_hd__and2_4
XANTENNA__17941__B1 _17811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21470_ _22687_/A VGND VGND VPWR VPWR _21806_/A sky130_fd_sc_hd__buf_2
XFILLER_159_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12844__B _12842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20421_ _20226_/X VGND VGND VPWR VPWR _20438_/A sky130_fd_sc_hd__buf_2
XANTENNA__15220__B _15156_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22293__A2 _22287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18497__B2 _18496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13021__A _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23140_ _23203_/CLK _23140_/D VGND VGND VPWR VPWR _15759_/B sky130_fd_sc_hd__dfxtp_4
X_20352_ _20352_/A VGND VGND VPWR VPWR _20352_/X sky130_fd_sc_hd__buf_2
XFILLER_101_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23071_ _19953_/A _17655_/A _23048_/X _23070_/X VGND VGND VPWR VPWR _23071_/X sky130_fd_sc_hd__a211o_4
XFILLER_161_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12860__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20283_ _24436_/Q _18837_/B _24468_/Q _20282_/X VGND VGND VPWR VPWR _20283_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16332__A _11714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22022_ _21857_/X _22017_/X _15523_/B _22021_/X VGND VGND VPWR VPWR _23521_/D sky130_fd_sc_hd__o22a_4
XFILLER_115_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20789__A _20267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21005__B1 _14895_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23973_ _23493_/CLK _23973_/D VGND VGND VPWR VPWR _23973_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20359__A2 _20304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14787__A _15103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22924_ _23078_/A _18661_/A _22924_/C VGND VGND VPWR VPWR _22926_/B sky130_fd_sc_hd__or3_4
XFILLER_17_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20764__C1 _20763_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22855_ _13342_/Y _22847_/X _22853_/X _22854_/X VGND VGND VPWR VPWR _22856_/A sky130_fd_sc_hd__a211o_4
XFILLER_147_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21308__B2 _21300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21806_ _21806_/A _21420_/B _21320_/C _22487_/B VGND VGND VPWR VPWR _21806_/X sky130_fd_sc_hd__or4_4
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22786_ _22784_/Y _22786_/B VGND VGND VPWR VPWR _22788_/B sky130_fd_sc_hd__or2_4
XANTENNA__12100__A _12061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21859__A2 _21851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21737_ _21570_/X _21734_/X _15477_/B _21731_/X VGND VGND VPWR VPWR _21737_/X sky130_fd_sc_hd__o22a_4
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12470_ _12470_/A VGND VGND VPWR VPWR _12492_/A sky130_fd_sc_hd__buf_2
X_21668_ _21536_/X _21663_/X _16445_/B _21667_/X VGND VGND VPWR VPWR _21668_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24456_ _23347_/CLK _24456_/D HRESETn VGND VGND VPWR VPWR _24456_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23407_ _23983_/CLK _23407_/D VGND VGND VPWR VPWR _16289_/B sky130_fd_sc_hd__dfxtp_4
X_20619_ _20619_/A _20494_/B VGND VGND VPWR VPWR _20619_/X sky130_fd_sc_hd__or2_4
XFILLER_165_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24387_ _24419_/CLK _18924_/X HRESETn VGND VGND VPWR VPWR _24387_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_126_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21599_ _21598_/X _21590_/X _23766_/Q _21524_/X VGND VGND VPWR VPWR _23766_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14027__A _13719_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20295__A1 _20235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14140_ _14140_/A _23615_/Q VGND VGND VPWR VPWR _14140_/X sky130_fd_sc_hd__or2_4
X_23338_ _23723_/CLK _22332_/X VGND VGND VPWR VPWR _12803_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19838__A2_N _19837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22244__A _22244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14071_ _11660_/A _23712_/Q VGND VGND VPWR VPWR _14071_/X sky130_fd_sc_hd__or2_4
XANTENNA__13866__A _13866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23269_ _23750_/CLK _23269_/D VGND VGND VPWR VPWR _23269_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22036__A2 _22031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17338__A _17339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12770__A _13349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13022_ _12506_/A _24072_/Q VGND VGND VPWR VPWR _13022_/X sky130_fd_sc_hd__or2_4
XFILLER_3_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17830_ _17813_/X _17822_/Y _17824_/X _17829_/Y VGND VGND VPWR VPWR _17830_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20699__A _20339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17761_ _17730_/X _17731_/X _17760_/X VGND VGND VPWR VPWR _17762_/C sky130_fd_sc_hd__or3_4
XANTENNA__13485__B1 _11608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14973_ _14973_/A _23478_/Q VGND VGND VPWR VPWR _14973_/X sky130_fd_sc_hd__or2_4
XANTENNA__14697__A _15625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21547__B2 _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22744__B1 _23086_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19500_ _19624_/A _19528_/B VGND VGND VPWR VPWR _19537_/B sky130_fd_sc_hd__or2_4
XANTENNA__18169__A _17452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16712_ _16594_/A _23601_/Q VGND VGND VPWR VPWR _16713_/C sky130_fd_sc_hd__or2_4
X_13924_ _14390_/A _13841_/B VGND VGND VPWR VPWR _13924_/X sky130_fd_sc_hd__or2_4
X_17692_ _17688_/A _17520_/X _17688_/X VGND VGND VPWR VPWR _17697_/B sky130_fd_sc_hd__a21bo_4
Xclkbuf_7_71_0_HCLK clkbuf_6_35_0_HCLK/X VGND VGND VPWR VPWR _23671_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19431_ _19399_/X _18699_/X _19402_/X _24216_/Q VGND VGND VPWR VPWR _19431_/X sky130_fd_sc_hd__o22a_4
XFILLER_35_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16643_ _16788_/A VGND VGND VPWR VPWR _16676_/A sky130_fd_sc_hd__buf_2
XFILLER_90_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13855_ _15444_/A _13930_/B VGND VGND VPWR VPWR _13855_/X sky130_fd_sc_hd__or2_4
XANTENNA__13106__A _13090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12806_ _13556_/A _12806_/B _12805_/X VGND VGND VPWR VPWR _12807_/C sky130_fd_sc_hd__or3_4
X_19362_ _19372_/A VGND VGND VPWR VPWR _19362_/X sky130_fd_sc_hd__buf_2
XFILLER_50_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12010__A _11939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16574_ _16558_/A _23634_/Q VGND VGND VPWR VPWR _16576_/B sky130_fd_sc_hd__or2_4
X_13786_ _11928_/A VGND VGND VPWR VPWR _14991_/A sky130_fd_sc_hd__buf_2
X_18313_ _18378_/A _17523_/Y VGND VGND VPWR VPWR _18313_/X sky130_fd_sc_hd__and2_4
XANTENNA__21323__A _21338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15525_ _12239_/A _15525_/B VGND VGND VPWR VPWR _15525_/X sky130_fd_sc_hd__or2_4
X_12737_ _13304_/A _24106_/Q VGND VGND VPWR VPWR _12738_/C sky130_fd_sc_hd__or2_4
X_19293_ _19240_/B VGND VGND VPWR VPWR _19293_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12945__A _12945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16417__A _11882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18244_ _17900_/A VGND VGND VPWR VPWR _18244_/X sky130_fd_sc_hd__buf_2
XANTENNA__15321__A _15321_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15456_ _14543_/A _15454_/X _15456_/C VGND VGND VPWR VPWR _15456_/X sky130_fd_sc_hd__and3_4
X_12668_ _12942_/A _12668_/B VGND VGND VPWR VPWR _12668_/X sky130_fd_sc_hd__or2_4
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12664__B _12664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _15487_/A _23644_/Q VGND VGND VPWR VPWR _14407_/X sky130_fd_sc_hd__or2_4
XANTENNA__19728__A _19724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18175_ _17490_/C _18175_/B VGND VGND VPWR VPWR _18175_/X sky130_fd_sc_hd__or2_4
X_11619_ _11877_/A VGND VGND VPWR VPWR _12299_/A sky130_fd_sc_hd__buf_2
XFILLER_117_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15387_ _14703_/A _15387_/B VGND VGND VPWR VPWR _15387_/X sky130_fd_sc_hd__and2_4
X_12599_ _12651_/A _12599_/B VGND VGND VPWR VPWR _12599_/X sky130_fd_sc_hd__or2_4
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17126_ _17339_/A _17107_/X _17015_/X _17074_/X VGND VGND VPWR VPWR _17126_/X sky130_fd_sc_hd__o22a_4
X_14338_ _14377_/A VGND VGND VPWR VPWR _14517_/A sky130_fd_sc_hd__buf_2
XFILLER_143_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22154__A _22118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13776__A _12610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17057_ _17103_/A _17057_/B VGND VGND VPWR VPWR _17085_/A sky130_fd_sc_hd__or2_4
XANTENNA__22027__A2 _22024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14269_ _14269_/A VGND VGND VPWR VPWR _14270_/A sky130_fd_sc_hd__buf_2
XANTENNA__16152__A _16138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16008_ _16007_/X _23726_/Q VGND VGND VPWR VPWR _16011_/B sky130_fd_sc_hd__or2_4
XANTENNA__21993__A _22000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18100__B1 _18009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21786__B2 _21781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17959_ _17959_/A _17657_/Y VGND VGND VPWR VPWR _17959_/X sky130_fd_sc_hd__and2_4
XANTENNA__21538__B2 _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18079__A _18283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20970_ _20425_/A _20969_/X _19228_/A _20349_/A VGND VGND VPWR VPWR _20970_/X sky130_fd_sc_hd__o22a_4
XFILLER_38_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14400__A _12583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19629_ _19629_/A VGND VGND VPWR VPWR _19797_/A sky130_fd_sc_hd__buf_2
XFILLER_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13016__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22640_ _22655_/A VGND VGND VPWR VPWR _22648_/A sky130_fd_sc_hd__buf_2
XFILLER_81_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22571_ _22459_/X _22565_/X _23200_/Q _22569_/X VGND VGND VPWR VPWR _23200_/D sky130_fd_sc_hd__o22a_4
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12855__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16327__A _13414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24310_ _24287_/CLK _19222_/X HRESETn VGND VGND VPWR VPWR _24310_/Q sky130_fd_sc_hd__dfrtp_4
X_21522_ _21521_/X VGND VGND VPWR VPWR _21523_/A sky130_fd_sc_hd__buf_2
XFILLER_22_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17390__A1 _15915_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24318__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17390__B2 _17389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24241_ _24240_/CLK _24241_/D HRESETn VGND VGND VPWR VPWR _24241_/Q sky130_fd_sc_hd__dfrtp_4
X_21453_ _21287_/X _21448_/X _15560_/B _21452_/X VGND VGND VPWR VPWR _23841_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22266__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20404_ _20404_/A VGND VGND VPWR VPWR _20404_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24172_ _23383_/CLK _24172_/D HRESETn VGND VGND VPWR VPWR _24172_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21384_ _21391_/A VGND VGND VPWR VPWR _21384_/X sky130_fd_sc_hd__buf_2
XANTENNA__22064__A _22057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23123_ _23764_/CLK _23123_/D VGND VGND VPWR VPWR _23123_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22018__A2 _22017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13686__A _12294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20335_ _24243_/Q _20304_/X _20334_/X VGND VGND VPWR VPWR _20336_/A sky130_fd_sc_hd__o21a_4
XANTENNA__12590__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22999__A _22998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23054_ _22931_/A _23054_/B VGND VGND VPWR VPWR _23056_/B sky130_fd_sc_hd__nand2_4
X_20266_ _20266_/A _20352_/A VGND VGND VPWR VPWR _20266_/X sky130_fd_sc_hd__or2_4
XFILLER_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22005_ _21829_/X _22003_/X _16167_/B _22000_/X VGND VGND VPWR VPWR _22005_/X sky130_fd_sc_hd__o22a_4
XFILLER_1_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20197_ _18623_/Y _20155_/Y _20196_/X VGND VGND VPWR VPWR _20197_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20312__A _20233_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15406__A _15406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11934__A _12266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11970_ _11970_/A VGND VGND VPWR VPWR _13453_/A sky130_fd_sc_hd__buf_2
X_23956_ _23764_/CLK _23956_/D VGND VGND VPWR VPWR _23956_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14310__A _14310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_58_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__20201__A1 _19906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22907_ _22906_/X VGND VGND VPWR VPWR HADDR[1] sky130_fd_sc_hd__inv_2
X_23887_ _23119_/CLK _21383_/X VGND VGND VPWR VPWR _16304_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13640_ _13677_/A _13636_/X _13640_/C VGND VGND VPWR VPWR _13641_/C sky130_fd_sc_hd__and3_4
X_22838_ _15453_/Y _22836_/X _22817_/X _22837_/X VGND VGND VPWR VPWR _22839_/B sky130_fd_sc_hd__o22a_4
XFILLER_60_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _13342_/Y _13417_/X VGND VGND VPWR VPWR _13581_/A sky130_fd_sc_hd__or2_4
XANTENNA__16237__A _16187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12765__A _12634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20504__A2 _20488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22769_ _22769_/A _22754_/X _22757_/X _22769_/D VGND VGND VPWR VPWR _22769_/X sky130_fd_sc_hd__or4_4
XANTENNA__21701__A1 _21594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21701__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15141__A _13791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15310_ _15029_/A _15306_/X _15310_/C VGND VGND VPWR VPWR _15310_/X sky130_fd_sc_hd__or3_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12522_ _12493_/A _12522_/B _12522_/C VGND VGND VPWR VPWR _12523_/C sky130_fd_sc_hd__and3_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16290_ _11904_/X _16290_/B VGND VGND VPWR VPWR _16290_/X sky130_fd_sc_hd__or2_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15241_ _14199_/A _15169_/B VGND VGND VPWR VPWR _15243_/B sky130_fd_sc_hd__or2_4
XANTENNA__19658__B1 _11611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19548__A _19687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24439_ _24445_/CLK _24439_/D HRESETn VGND VGND VPWR VPWR _24439_/Q sky130_fd_sc_hd__dfrtp_4
X_12453_ _12453_/A VGND VGND VPWR VPWR _12454_/A sky130_fd_sc_hd__buf_2
XANTENNA__22257__A2 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12384_ _11739_/A _12384_/B _12384_/C VGND VGND VPWR VPWR _12384_/X sky130_fd_sc_hd__and3_4
X_15172_ _13617_/A _15172_/B VGND VGND VPWR VPWR _15172_/X sky130_fd_sc_hd__or2_4
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14123_ _13788_/A _14112_/X _14122_/X VGND VGND VPWR VPWR _14123_/X sky130_fd_sc_hd__or3_4
XANTENNA__13596__A _13596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22009__A2 _22003_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19980_ _19961_/X _19977_/X _19978_/Y _19979_/X VGND VGND VPWR VPWR _19980_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18881__A1 _14844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18931_ _17153_/A _18927_/X _24382_/Q _18928_/X VGND VGND VPWR VPWR _24382_/D sky130_fd_sc_hd__o22a_4
X_14054_ _13719_/A _14052_/X _14053_/X VGND VGND VPWR VPWR _14054_/X sky130_fd_sc_hd__and3_4
XANTENNA__21768__B2 _21767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14204__B _23935_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13005_ _12510_/A _23336_/Q VGND VGND VPWR VPWR _13007_/B sky130_fd_sc_hd__or2_4
X_18862_ _17172_/X _18856_/X _24422_/Q _18857_/X VGND VGND VPWR VPWR _24422_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12005__A _12106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17813_ _17812_/X VGND VGND VPWR VPWR _17813_/X sky130_fd_sc_hd__buf_2
XANTENNA__21318__A _21028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17515__B _17515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18793_ _17255_/X _18787_/X _24466_/Q _18790_/X VGND VGND VPWR VPWR _18793_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22717__B1 _15840_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17744_ _17744_/A _17743_/X VGND VGND VPWR VPWR _17744_/X sky130_fd_sc_hd__or2_4
X_14956_ _14925_/X _14954_/X _14955_/X VGND VGND VPWR VPWR _14956_/X sky130_fd_sc_hd__and3_4
XANTENNA__23985__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14220__A _12336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22193__B2 _22191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13907_ _13710_/A _13818_/B VGND VGND VPWR VPWR _13907_/X sky130_fd_sc_hd__or2_4
X_17675_ _17675_/A _17473_/Y VGND VGND VPWR VPWR _17675_/X sky130_fd_sc_hd__and2_4
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14887_ _14127_/A _14958_/B VGND VGND VPWR VPWR _14889_/B sky130_fd_sc_hd__or2_4
XFILLER_78_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19414_ _19406_/X VGND VGND VPWR VPWR _19414_/X sky130_fd_sc_hd__buf_2
XFILLER_78_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16626_ _16639_/A VGND VGND VPWR VPWR _16658_/A sky130_fd_sc_hd__buf_2
X_13838_ _12497_/A _13838_/B VGND VGND VPWR VPWR _13838_/X sky130_fd_sc_hd__or2_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22149__A _20818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19345_ _19343_/X _18142_/X _19343_/X _24269_/Q VGND VGND VPWR VPWR _24269_/D sky130_fd_sc_hd__a2bb2o_4
X_16557_ _12001_/A VGND VGND VPWR VPWR _16588_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_1_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR _24292_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12675__A _12977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13769_ _12610_/A _13769_/B VGND VGND VPWR VPWR _13769_/X sky130_fd_sc_hd__or2_4
XANTENNA__19897__B1 _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22496__A2 _22494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15051__A _12329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15508_ _13744_/A _15508_/B VGND VGND VPWR VPWR _15508_/X sky130_fd_sc_hd__or2_4
XFILLER_148_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19276_ _24299_/Q _19248_/B _19275_/Y VGND VGND VPWR VPWR _19276_/X sky130_fd_sc_hd__o21a_4
XFILLER_149_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16488_ _11784_/X _16478_/X _16487_/X VGND VGND VPWR VPWR _16489_/C sky130_fd_sc_hd__and3_4
XANTENNA__20892__A _20892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18227_ _17876_/X _17845_/Y _17833_/A _17864_/Y VGND VGND VPWR VPWR _18227_/X sky130_fd_sc_hd__o22a_4
XFILLER_148_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15439_ _15439_/A _15511_/B VGND VGND VPWR VPWR _15439_/X sky130_fd_sc_hd__or2_4
XANTENNA__15383__B1 _15185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18158_ _17986_/X _17983_/X _17988_/X _17987_/X VGND VGND VPWR VPWR _18158_/X sky130_fd_sc_hd__o22a_4
XFILLER_11_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17109_ _17108_/X VGND VGND VPWR VPWR _17109_/X sky130_fd_sc_hd__buf_2
XFILLER_89_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18089_ _17869_/X VGND VGND VPWR VPWR _18089_/X sky130_fd_sc_hd__buf_2
XANTENNA__18872__A1 _17161_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16913__A1_N _16905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15686__A1 _13339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21208__B1 _23975_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20120_ _11572_/X _11574_/X VGND VGND VPWR VPWR _20120_/X sky130_fd_sc_hd__or2_4
XANTENNA__21812__A2_N _21810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20051_ _24485_/Q VGND VGND VPWR VPWR _20051_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11754__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23810_ _23650_/CLK _23810_/D VGND VGND VPWR VPWR _15502_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15226__A _14225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19921__A _19920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12569__B _12665_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23741_ _23678_/CLK _21644_/X VGND VGND VPWR VPWR _23741_/Q sky130_fd_sc_hd__dfxtp_4
X_20953_ _18696_/X _20342_/X _20753_/X _20952_/Y VGND VGND VPWR VPWR _20953_/X sky130_fd_sc_hd__a211o_4
XFILLER_22_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21931__B2 _21927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17441__A _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _20930_/A _20883_/X VGND VGND VPWR VPWR _20884_/Y sky130_fd_sc_hd__nor2_4
X_23672_ _23098_/CLK _23672_/D VGND VGND VPWR VPWR _23672_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24140__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22623_ _22461_/X _22622_/X _23167_/Q _22619_/X VGND VGND VPWR VPWR _22623_/X sky130_fd_sc_hd__o22a_4
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23708__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22554_ _22430_/X _22551_/X _12344_/B _22548_/X VGND VGND VPWR VPWR _23212_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21505_ _21290_/X _21499_/X _14068_/B _21503_/X VGND VGND VPWR VPWR _21505_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22239__A2 _22237_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22485_ _22484_/X _22438_/A _23253_/Q _22421_/A VGND VGND VPWR VPWR _23253_/D sky130_fd_sc_hd__o22a_4
XFILLER_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24290__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21436_ _21259_/X _21434_/X _16140_/B _21431_/X VGND VGND VPWR VPWR _21436_/X sky130_fd_sc_hd__o22a_4
X_24224_ _24137_/CLK _19420_/X HRESETn VGND VGND VPWR VPWR _24224_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20307__A _18779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21998__B2 _21993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24155_ _24306_/CLK _24155_/D HRESETn VGND VGND VPWR VPWR _24155_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21367_ _21313_/X _21362_/X _14880_/B _21331_/A VGND VGND VPWR VPWR _23894_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14305__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23106_ _23523_/CLK _23106_/D VGND VGND VPWR VPWR _15501_/B sky130_fd_sc_hd__dfxtp_4
X_20318_ _20318_/A _20318_/B VGND VGND VPWR VPWR _20318_/Y sky130_fd_sc_hd__nand2_4
X_24086_ _23544_/CLK _24086_/D VGND VGND VPWR VPWR _14895_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__11648__B _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21298_ _21297_/X _21293_/X _13896_/B _21288_/X VGND VGND VPWR VPWR _23933_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22522__A _22489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23037_ _22912_/X VGND VGND VPWR VPWR _23051_/A sky130_fd_sc_hd__buf_2
X_20249_ _20249_/A VGND VGND VPWR VPWR _20308_/A sky130_fd_sc_hd__buf_2
XANTENNA__16520__A _11815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21138__A _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20042__A _19950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14810_ _14682_/A _14810_/B _14810_/C VGND VGND VPWR VPWR _14811_/C sky130_fd_sc_hd__and3_4
XFILLER_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15790_ _11902_/A _15790_/B VGND VGND VPWR VPWR _15790_/X sky130_fd_sc_hd__or2_4
XANTENNA__14040__A _11698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20977__A _20977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14741_ _13622_/A _14741_/B _14741_/C VGND VGND VPWR VPWR _14742_/C sky130_fd_sc_hd__and3_4
X_23939_ _23939_/CLK _21284_/X VGND VGND VPWR VPWR _15865_/B sky130_fd_sc_hd__dfxtp_4
X_11953_ _12102_/A _21705_/A VGND VGND VPWR VPWR _11957_/B sky130_fd_sc_hd__or2_4
XFILLER_45_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21922__B2 _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17460_ _12982_/X _17460_/B VGND VGND VPWR VPWR _17460_/X sky130_fd_sc_hd__and2_4
XFILLER_33_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14672_ _14840_/A _14667_/X _14672_/C VGND VGND VPWR VPWR _14682_/B sky130_fd_sc_hd__or3_4
X_11884_ _16155_/A VGND VGND VPWR VPWR _16116_/A sky130_fd_sc_hd__buf_2
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14694__B _14600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16411_ _16159_/A _16407_/X _16411_/C VGND VGND VPWR VPWR _16411_/X sky130_fd_sc_hd__or3_4
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13623_ _12497_/A _24030_/Q VGND VGND VPWR VPWR _13625_/B sky130_fd_sc_hd__or2_4
XFILLER_38_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17391_ _15913_/Y _17448_/B VGND VGND VPWR VPWR _17391_/X sky130_fd_sc_hd__or2_4
X_19130_ _19223_/A _24309_/Q VGND VGND VPWR VPWR _19131_/B sky130_fd_sc_hd__and2_4
X_16342_ _16342_/A _16267_/B VGND VGND VPWR VPWR _16343_/C sky130_fd_sc_hd__or2_4
XFILLER_9_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13554_ _13554_/A _13480_/B VGND VGND VPWR VPWR _13555_/C sky130_fd_sc_hd__or2_4
XANTENNA__21150__A2 _21148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12505_ _12540_/A VGND VGND VPWR VPWR _12506_/A sky130_fd_sc_hd__buf_2
X_19061_ _19046_/X _19059_/Y _19060_/Y _19049_/X VGND VGND VPWR VPWR _19061_/X sky130_fd_sc_hd__o22a_4
X_16273_ _16096_/A _16273_/B VGND VGND VPWR VPWR _16273_/X sky130_fd_sc_hd__or2_4
X_13485_ _11858_/A _11631_/X _13454_/X _11608_/A _13484_/X VGND VGND VPWR VPWR _13485_/X
+ sky130_fd_sc_hd__a32o_4
X_18012_ _17963_/X _17966_/X _17014_/X _18011_/X VGND VGND VPWR VPWR _18012_/X sky130_fd_sc_hd__o22a_4
X_15224_ _14201_/A _15222_/X _15224_/C VGND VGND VPWR VPWR _15225_/C sky130_fd_sc_hd__and3_4
X_12436_ _12852_/A VGND VGND VPWR VPWR _12847_/A sky130_fd_sc_hd__buf_2
XFILLER_172_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15155_ _14154_/A _15155_/B VGND VGND VPWR VPWR _15157_/B sky130_fd_sc_hd__or2_4
XANTENNA__18854__A1 _12419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12367_ _12367_/A VGND VGND VPWR VPWR _13251_/A sky130_fd_sc_hd__buf_2
XANTENNA__22650__A2 _22644_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14106_ _14003_/A _14106_/B _14105_/X VGND VGND VPWR VPWR _14107_/C sky130_fd_sc_hd__and3_4
X_12298_ _12298_/A _12293_/X _12297_/X VGND VGND VPWR VPWR _12308_/B sky130_fd_sc_hd__and3_4
X_19963_ _18037_/X _19963_/B VGND VGND VPWR VPWR _19966_/B sky130_fd_sc_hd__nor2_4
X_15086_ _15086_/A _23957_/Q VGND VGND VPWR VPWR _15087_/C sky130_fd_sc_hd__or2_4
XANTENNA__22432__A _22117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18914_ _18900_/A VGND VGND VPWR VPWR _18914_/X sky130_fd_sc_hd__buf_2
XFILLER_80_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14037_ _13719_/A _14035_/X _14037_/C VGND VGND VPWR VPWR _14037_/X sky130_fd_sc_hd__and3_4
XANTENNA__22402__A2 _22397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16430__A _15998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19894_ _19507_/A _19507_/B _19894_/C _19903_/B VGND VGND VPWR VPWR _19894_/X sky130_fd_sc_hd__and4_4
XANTENNA__22542__A2_N _22541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13773__B _24094_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18845_ _12180_/X _18840_/X _20318_/A _18843_/X VGND VGND VPWR VPWR _24435_/D sky130_fd_sc_hd__o22a_4
XFILLER_121_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24385__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18776_ _24131_/Q _17343_/X _17752_/X VGND VGND VPWR VPWR _18776_/Y sky130_fd_sc_hd__o21ai_4
X_15988_ _15957_/A _15988_/B VGND VGND VPWR VPWR _15990_/B sky130_fd_sc_hd__or2_4
XANTENNA__22166__A1 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22166__B2 _22106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17727_ _17727_/A _17399_/X VGND VGND VPWR VPWR _17727_/X sky130_fd_sc_hd__or2_4
XANTENNA__24163__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14939_ _14970_/A _14875_/B VGND VGND VPWR VPWR _14939_/X sky130_fd_sc_hd__or2_4
XFILLER_24_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_41_0_HCLK clkbuf_5_20_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17658_ _16948_/A _17548_/X VGND VGND VPWR VPWR _17663_/A sky130_fd_sc_hd__and2_4
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17593__A1 _17132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16609_ _16621_/A _16609_/B VGND VGND VPWR VPWR _16609_/X sky130_fd_sc_hd__or2_4
X_17589_ _17583_/B _17587_/X _17588_/Y VGND VGND VPWR VPWR _17589_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19328_ _19328_/A VGND VGND VPWR VPWR _19328_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14109__B _23679_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19259_ _24308_/Q _19258_/A _19257_/Y _19258_/Y VGND VGND VPWR VPWR _19259_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16605__A _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18092__A _18562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22270_ _22167_/X _22265_/X _14961_/B _22226_/X VGND VGND VPWR VPWR _23382_/D sky130_fd_sc_hd__o22a_4
XFILLER_145_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21221_ _20819_/X _21219_/X _23966_/Q _21216_/X VGND VGND VPWR VPWR _21221_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11749__A _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19916__A _23083_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18845__A1 _12180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21152_ _21152_/A VGND VGND VPWR VPWR _21152_/X sky130_fd_sc_hd__buf_2
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20103_ _19433_/X _20102_/X _19433_/X _24138_/Q VGND VGND VPWR VPWR _24138_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21083_ _21134_/A _21370_/B _21184_/C _22487_/B VGND VGND VPWR VPWR _21083_/X sky130_fd_sc_hd__or4_4
XANTENNA__14779__B _14779_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20034_ _20016_/X _17681_/A _20022_/X _20033_/X VGND VGND VPWR VPWR _20034_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21601__B1 _23765_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13683__B _13766_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_123_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR _23561_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20955__A2 _20946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22157__B2 _22154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21985_ _21881_/X _21981_/X _15143_/B _21950_/A VGND VGND VPWR VPWR _23543_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21904__B2 _21899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23724_ _24045_/CLK _23724_/D VGND VGND VPWR VPWR _23724_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _24217_/Q _20895_/X _20935_/X VGND VGND VPWR VPWR _20937_/A sky130_fd_sc_hd__o21a_4
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21380__A2 _21377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23655_ _23750_/CLK _23655_/D VGND VGND VPWR VPWR _23655_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15403__B _15466_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _20867_/A _20672_/A VGND VGND VPWR VPWR _20867_/X sky130_fd_sc_hd__or2_4
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13204__A _13230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22606_ _22432_/X _22601_/X _12520_/B _22605_/X VGND VGND VPWR VPWR _23179_/D sky130_fd_sc_hd__o22a_4
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23586_ _23587_/CLK _23586_/D VGND VGND VPWR VPWR _15471_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20798_ _20935_/A _20797_/X VGND VGND VPWR VPWR _20798_/X sky130_fd_sc_hd__or2_4
XANTENNA__17336__A1 _12570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20340__B1 _20235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22537_ _22090_/A _22687_/B _21319_/A _22537_/D VGND VGND VPWR VPWR _22537_/X sky130_fd_sc_hd__or4_4
XFILLER_127_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13270_ _13270_/A VGND VGND VPWR VPWR _13270_/X sky130_fd_sc_hd__buf_2
X_22468_ _20859_/A VGND VGND VPWR VPWR _22468_/X sky130_fd_sc_hd__buf_2
XFILLER_108_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12221_ _13676_/A VGND VGND VPWR VPWR _12269_/A sky130_fd_sc_hd__buf_2
X_24207_ _24184_/CLK _24207_/D HRESETn VGND VGND VPWR VPWR _17274_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24487__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11659__A _11659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21419_ _23860_/Q VGND VGND VPWR VPWR _21419_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22632__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22399_ _22161_/X _22397_/X _14717_/B _22394_/X VGND VGND VPWR VPWR _22399_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14035__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12152_ _11746_/X _24083_/Q VGND VGND VPWR VPWR _12152_/X sky130_fd_sc_hd__or2_4
X_24138_ _24137_/CLK _24138_/D HRESETn VGND VGND VPWR VPWR _24138_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_2_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16960_ _24146_/Q VGND VGND VPWR VPWR _17708_/A sky130_fd_sc_hd__inv_2
XANTENNA__17346__A _16866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12083_ _12059_/X _24083_/Q VGND VGND VPWR VPWR _12083_/X sky130_fd_sc_hd__or2_4
X_24069_ _23493_/CLK _21058_/X VGND VGND VPWR VPWR _24069_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21199__A2 _21198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15911_ _12676_/A _15911_/B _15911_/C VGND VGND VPWR VPWR _15912_/C sky130_fd_sc_hd__or3_4
XANTENNA__22396__B2 _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24186__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16891_ _12986_/B _16832_/X _12983_/X VGND VGND VPWR VPWR _16891_/X sky130_fd_sc_hd__o21a_4
X_18630_ _18628_/X _17749_/A _18630_/C VGND VGND VPWR VPWR _18630_/X sky130_fd_sc_hd__or3_4
X_15842_ _12862_/A _15842_/B _15842_/C VGND VGND VPWR VPWR _15842_/X sky130_fd_sc_hd__and3_4
XANTENNA__19561__A _19450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22148__B2 _22142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18561_ _17436_/B _18560_/B VGND VGND VPWR VPWR _18561_/X sky130_fd_sc_hd__or2_4
XFILLER_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15773_ _11689_/X _15769_/X _15773_/C VGND VGND VPWR VPWR _15781_/B sky130_fd_sc_hd__or3_4
XANTENNA__22699__A2 _22694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12985_ _12914_/X _12982_/X _12984_/Y VGND VGND VPWR VPWR _12986_/B sky130_fd_sc_hd__a21o_4
XFILLER_131_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17512_ _13049_/Y _17022_/X _17031_/A _17511_/X VGND VGND VPWR VPWR _17515_/B sky130_fd_sc_hd__o22a_4
XFILLER_45_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17081__A _17017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_28_0_HCLK clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14724_ _15444_/A _14724_/B VGND VGND VPWR VPWR _14725_/C sky130_fd_sc_hd__or2_4
X_11936_ _12904_/A VGND VGND VPWR VPWR _15978_/A sky130_fd_sc_hd__buf_2
X_18492_ _17396_/A _18491_/X VGND VGND VPWR VPWR _18492_/X sky130_fd_sc_hd__or2_4
XFILLER_18_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17443_ _17162_/Y _17421_/B _17436_/C _17442_/X VGND VGND VPWR VPWR _17443_/X sky130_fd_sc_hd__o22a_4
X_14655_ _14685_/A _14655_/B _14655_/C VGND VGND VPWR VPWR _14660_/B sky130_fd_sc_hd__and3_4
XFILLER_162_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11867_ _16160_/A VGND VGND VPWR VPWR _11867_/X sky130_fd_sc_hd__buf_2
XFILLER_159_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13114__A _13090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13606_ _13606_/A VGND VGND VPWR VPWR _13607_/A sky130_fd_sc_hd__buf_2
X_17374_ _17374_/A VGND VGND VPWR VPWR _17375_/B sky130_fd_sc_hd__inv_2
X_14586_ _12530_/A _23610_/Q VGND VGND VPWR VPWR _14586_/X sky130_fd_sc_hd__or2_4
X_11798_ _11694_/X VGND VGND VPWR VPWR _12169_/A sky130_fd_sc_hd__buf_2
XFILLER_13_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22320__B2 _22284_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19113_ _19109_/X _19112_/X _19109_/X _11519_/A VGND VGND VPWR VPWR _24345_/D sky130_fd_sc_hd__a2bb2o_4
X_16325_ _16318_/A _16260_/B VGND VGND VPWR VPWR _16325_/X sky130_fd_sc_hd__or2_4
XANTENNA__21331__A _21331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13537_ _13520_/A _13533_/X _13537_/C VGND VGND VPWR VPWR _13549_/B sky130_fd_sc_hd__or3_4
XFILLER_9_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19044_ _19016_/X _19042_/X _19043_/Y _19021_/X VGND VGND VPWR VPWR _19044_/X sky130_fd_sc_hd__o22a_4
X_16256_ _16156_/A _16256_/B VGND VGND VPWR VPWR _16256_/X sky130_fd_sc_hd__or2_4
X_13468_ _13468_/A _13464_/X _13468_/C VGND VGND VPWR VPWR _13468_/X sky130_fd_sc_hd__or3_4
XFILLER_139_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12672__B _12672_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15207_ _14669_/A _15150_/B VGND VGND VPWR VPWR _15207_/X sky130_fd_sc_hd__or2_4
X_12419_ _12418_/X VGND VGND VPWR VPWR _12419_/X sky130_fd_sc_hd__buf_2
XANTENNA__18827__A1 _17290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16187_ _16187_/A _16187_/B _16187_/C VGND VGND VPWR VPWR _16207_/B sky130_fd_sc_hd__and3_4
X_13399_ _13399_/A _13399_/B _13399_/C VGND VGND VPWR VPWR _13400_/C sky130_fd_sc_hd__or3_4
XFILLER_114_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18640__A _18545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20634__A1 _20533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20634__B2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15138_ _14277_/A _15131_/X _15137_/X VGND VGND VPWR VPWR _15138_/X sky130_fd_sc_hd__or3_4
XFILLER_153_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17256__A _17255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19946_ _24129_/Q VGND VGND VPWR VPWR _22908_/A sky130_fd_sc_hd__buf_2
X_15069_ _14073_/A _15069_/B _15069_/C VGND VGND VPWR VPWR _15069_/X sky130_fd_sc_hd__and3_4
XFILLER_68_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19877_ _19834_/A _19711_/A _19811_/A VGND VGND VPWR VPWR _19877_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18828_ _14844_/X _18824_/X _20923_/A _18825_/X VGND VGND VPWR VPWR _24441_/D sky130_fd_sc_hd__o22a_4
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21506__A _21506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17703__B _17483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18759_ _17101_/A _17626_/A _18674_/A _18758_/X VGND VGND VPWR VPWR _18759_/X sky130_fd_sc_hd__o22a_4
X_21770_ _21770_/A VGND VGND VPWR VPWR _21770_/X sky130_fd_sc_hd__buf_2
XANTENNA__18763__B1 _17037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20721_ HRDATA[12] _20697_/A VGND VGND VPWR VPWR _20721_/X sky130_fd_sc_hd__or2_4
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13024__A _12881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23440_ _24080_/CLK _23440_/D VGND VGND VPWR VPWR _16432_/B sky130_fd_sc_hd__dfxtp_4
X_20652_ _20652_/A _20651_/X VGND VGND VPWR VPWR _20652_/Y sky130_fd_sc_hd__nor2_4
XFILLER_11_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21114__A2 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22311__B2 _22305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23371_ _23723_/CLK _22292_/X VGND VGND VPWR VPWR _23371_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_149_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13959__A _15029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20583_ _20583_/A VGND VGND VPWR VPWR _20583_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12863__A _12863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24059__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_48_0_HCLK clkbuf_7_49_0_HCLK/A VGND VGND VPWR VPWR _23537_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22322_ _11804_/B VGND VGND VPWR VPWR _23348_/D sky130_fd_sc_hd__buf_2
XFILLER_165_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22253_ _22137_/X _22251_/X _15829_/B _22248_/X VGND VGND VPWR VPWR _22253_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22075__B1 _23487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22614__A2 _22608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21204_ _20531_/X _21198_/X _23978_/Q _21202_/X VGND VGND VPWR VPWR _21204_/X sky130_fd_sc_hd__o22a_4
X_22184_ _22184_/A VGND VGND VPWR VPWR _22184_/X sky130_fd_sc_hd__buf_2
XFILLER_133_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21135_ _21134_/X VGND VGND VPWR VPWR _21136_/A sky130_fd_sc_hd__buf_2
XANTENNA__22378__B2 _22373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21066_ _21033_/A VGND VGND VPWR VPWR _21066_/X sky130_fd_sc_hd__buf_2
XFILLER_59_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22800__A _16922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20017_ _20017_/A VGND VGND VPWR VPWR _20017_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19381__A _19377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21050__B2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11942__A _16713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15414__A _13655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12770_ _13349_/A _12768_/X _12769_/X VGND VGND VPWR VPWR _12770_/X sky130_fd_sc_hd__and3_4
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21968_ _21850_/X _21967_/X _15675_/B _21964_/X VGND VGND VPWR VPWR _23556_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21353__A2 _21348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22550__B2 _22548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _23675_/CLK _23707_/D VGND VGND VPWR VPWR _14534_/B sky130_fd_sc_hd__dfxtp_4
X_11721_ _13868_/A VGND VGND VPWR VPWR _15606_/A sky130_fd_sc_hd__buf_2
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ _20864_/A _20917_/X _20918_/X HRDATA[12] _20869_/A VGND VGND VPWR VPWR _20919_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ _21899_/A VGND VGND VPWR VPWR _21899_/X sky130_fd_sc_hd__buf_2
XFILLER_70_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _13010_/A _14440_/B VGND VGND VPWR VPWR _14440_/X sky130_fd_sc_hd__or2_4
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23638_ _23770_/CLK _23638_/D VGND VGND VPWR VPWR _23638_/Q sky130_fd_sc_hd__dfxtp_4
X_11652_ _13865_/A VGND VGND VPWR VPWR _15616_/A sky130_fd_sc_hd__buf_2
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21105__A2 _21104_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22302__B2 _22298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13869__A _13877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14371_ _13752_/A _14369_/X _14371_/C VGND VGND VPWR VPWR _14372_/C sky130_fd_sc_hd__and3_4
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12773__A _12944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23569_ _23761_/CLK _23569_/D VGND VGND VPWR VPWR _23569_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11583_ _24466_/Q IRQ[29] _20188_/A VGND VGND VPWR VPWR _11583_/X sky130_fd_sc_hd__a21o_4
XFILLER_70_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16110_ _16110_/A _16110_/B _16110_/C VGND VGND VPWR VPWR _16111_/C sky130_fd_sc_hd__and3_4
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _12516_/A _13318_/X _13322_/C VGND VGND VPWR VPWR _13322_/X sky130_fd_sc_hd__or3_4
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17090_ _17090_/A _17090_/B VGND VGND VPWR VPWR _17090_/X sky130_fd_sc_hd__and2_4
XFILLER_6_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16041_ _16048_/A _16041_/B VGND VGND VPWR VPWR _16041_/X sky130_fd_sc_hd__or2_4
X_13253_ _13253_/A _24103_/Q VGND VGND VPWR VPWR _13254_/C sky130_fd_sc_hd__or2_4
XFILLER_108_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18809__A1 _17172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12204_ _12693_/A _12204_/B VGND VGND VPWR VPWR _12204_/X sky130_fd_sc_hd__or2_4
XFILLER_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16899__B _16898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_5_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__23078__A _23078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13184_ _13184_/A _23815_/Q VGND VGND VPWR VPWR _13184_/X sky130_fd_sc_hd__or2_4
XFILLER_135_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19800_ _19681_/B _19798_/X _19809_/A VGND VGND VPWR VPWR _19800_/X sky130_fd_sc_hd__o21a_4
XFILLER_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12135_ _12166_/A _12135_/B VGND VGND VPWR VPWR _12135_/X sky130_fd_sc_hd__or2_4
XFILLER_150_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23576__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17992_ _17977_/X _17984_/Y _17985_/X _17991_/Y VGND VGND VPWR VPWR _17992_/X sky130_fd_sc_hd__o22a_4
XFILLER_145_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20214__B _21028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19731_ _19441_/X _19730_/X _17813_/X _19700_/X VGND VGND VPWR VPWR _24202_/D sky130_fd_sc_hd__o22a_4
X_16943_ _16943_/A VGND VGND VPWR VPWR _16943_/X sky130_fd_sc_hd__buf_2
XFILLER_133_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12066_ _16732_/A _12063_/X _12065_/X VGND VGND VPWR VPWR _12066_/X sky130_fd_sc_hd__and3_4
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21041__B2 _21035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19662_ _19659_/Y _19662_/B VGND VGND VPWR VPWR _19662_/X sky130_fd_sc_hd__and2_4
X_16874_ _16873_/X VGND VGND VPWR VPWR _16874_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12013__A _11951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15825_ _12866_/A _15821_/X _15824_/X VGND VGND VPWR VPWR _15825_/X sky130_fd_sc_hd__or3_4
X_18613_ _17890_/X _18605_/Y _18606_/X _18009_/X _18612_/X VGND VGND VPWR VPWR _18613_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21326__A _21322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19593_ _19589_/A VGND VGND VPWR VPWR _19681_/A sky130_fd_sc_hd__inv_2
XANTENNA__12948__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11852__A _11603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15756_ _15743_/X _15756_/B VGND VGND VPWR VPWR _15756_/X sky130_fd_sc_hd__or2_4
X_18544_ _18518_/X _17429_/X _17798_/A VGND VGND VPWR VPWR _18544_/X sky130_fd_sc_hd__a21o_4
X_12968_ _12944_/A _12966_/X _12967_/X VGND VGND VPWR VPWR _12968_/X sky130_fd_sc_hd__and3_4
XANTENNA__21344__A2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14707_ _13799_/A _23513_/Q VGND VGND VPWR VPWR _14708_/C sky130_fd_sc_hd__or2_4
XANTENNA__11571__B IRQ[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11919_ _16123_/A VGND VGND VPWR VPWR _16148_/A sky130_fd_sc_hd__buf_2
X_18475_ _18356_/X _18473_/X _18396_/X _18474_/X VGND VGND VPWR VPWR _18475_/X sky130_fd_sc_hd__o22a_4
X_15687_ _12696_/A _23908_/Q VGND VGND VPWR VPWR _15687_/X sky130_fd_sc_hd__or2_4
XANTENNA__20552__B1 _20538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12899_ _12872_/A _24105_/Q VGND VGND VPWR VPWR _12900_/C sky130_fd_sc_hd__or2_4
XFILLER_166_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17426_ _24210_/Q VGND VGND VPWR VPWR _17427_/A sky130_fd_sc_hd__inv_2
X_14638_ _14653_/A _14563_/B VGND VGND VPWR VPWR _14640_/B sky130_fd_sc_hd__or2_4
XFILLER_92_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13779__A _12576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17357_ _17357_/A _17357_/B VGND VGND VPWR VPWR _17358_/B sky130_fd_sc_hd__and2_4
X_14569_ _14448_/A _14567_/X _14569_/C VGND VGND VPWR VPWR _14573_/B sky130_fd_sc_hd__and3_4
XFILLER_158_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16308_ _16130_/A _16285_/X _16292_/X _16299_/X _16307_/X VGND VGND VPWR VPWR _16308_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_14_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24338__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21996__A _22010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17288_ _17287_/X VGND VGND VPWR VPWR _17292_/B sky130_fd_sc_hd__inv_2
X_19027_ _19016_/X _19025_/Y _19026_/Y _19021_/X VGND VGND VPWR VPWR _19027_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15994__A _15971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16239_ _13417_/A _16239_/B _16238_/X VGND VGND VPWR VPWR _16239_/X sky130_fd_sc_hd__and3_4
XFILLER_174_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20607__A1 _18350_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14403__A _14510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20124__B _20124_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19225__A1 _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19929_ _19921_/X _24176_/Q _19925_/X _20364_/B VGND VGND VPWR VPWR _24176_/D sky130_fd_sc_hd__o22a_4
XFILLER_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13019__A _12487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22940_ _22908_/X _17738_/X _22909_/X _22939_/X VGND VGND VPWR VPWR _22940_/X sky130_fd_sc_hd__a211o_4
XFILLER_96_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21583__A2 _21578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21236__A _21134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13961__B _23776_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22871_ _22870_/X VGND VGND VPWR VPWR HWDATA[22] sky130_fd_sc_hd__inv_2
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12858__A _12858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11762__A _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21822_ _21809_/X VGND VGND VPWR VPWR _21822_/X sky130_fd_sc_hd__buf_2
XFILLER_110_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21335__A2 _21334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22532__B2 _22526_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_11_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21753_ _21598_/X _21748_/X _14864_/B _21717_/A VGND VGND VPWR VPWR _23670_/D sky130_fd_sc_hd__o22a_4
XFILLER_19_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18545__A _18545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20704_ _20450_/B VGND VGND VPWR VPWR _20704_/X sky130_fd_sc_hd__buf_2
XANTENNA__15888__B _15826_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24472_ _24472_/CLK _18707_/Y HRESETn VGND VGND VPWR VPWR _24472_/Q sky130_fd_sc_hd__dfrtp_4
X_21684_ _21677_/A VGND VGND VPWR VPWR _21684_/X sky130_fd_sc_hd__buf_2
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22067__A _22060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21099__B2 _21094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13689__A _13689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23423_ _23294_/CLK _22209_/X VGND VGND VPWR VPWR _23423_/Q sky130_fd_sc_hd__dfxtp_4
X_20635_ _20533_/A VGND VGND VPWR VPWR _20635_/X sky130_fd_sc_hd__buf_2
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12593__A _12971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20566_ _20516_/X _20565_/X _24360_/Q _20475_/X VGND VGND VPWR VPWR _20566_/X sky130_fd_sc_hd__o22a_4
X_23354_ _24057_/CLK _22316_/X VGND VGND VPWR VPWR _23354_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22305_ _22291_/A VGND VGND VPWR VPWR _22305_/X sky130_fd_sc_hd__buf_2
XFILLER_165_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19376__A _19324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20497_ _20497_/A VGND VGND VPWR VPWR _20497_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18280__A _18406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23285_ _23392_/CLK _23285_/D VGND VGND VPWR VPWR _23285_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_164_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22599__B2 _22598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22236_ _22108_/X _22230_/X _16289_/B _22234_/X VGND VGND VPWR VPWR _23407_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15409__A _12191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22167_ _22482_/A VGND VGND VPWR VPWR _22167_/X sky130_fd_sc_hd__buf_2
XFILLER_132_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14313__A _14448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21118_ _21118_/A VGND VGND VPWR VPWR _21118_/X sky130_fd_sc_hd__buf_2
XFILLER_59_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19823__B _19823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22098_ _22147_/A VGND VGND VPWR VPWR _22123_/A sky130_fd_sc_hd__buf_2
XFILLER_75_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21049_ _21049_/A VGND VGND VPWR VPWR _21049_/X sky130_fd_sc_hd__buf_2
X_13940_ _13706_/A _23645_/Q VGND VGND VPWR VPWR _13940_/X sky130_fd_sc_hd__or2_4
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21574__A2 _21566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22771__A1 SYSTICKCLKDIV[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13871_ _13923_/A _13867_/X _13870_/X VGND VGND VPWR VPWR _13871_/X sky130_fd_sc_hd__and3_4
XFILLER_35_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16450__A1 _16130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15610_ _15610_/A _23681_/Q VGND VGND VPWR VPWR _15612_/B sky130_fd_sc_hd__or2_4
X_12822_ _13556_/A _12818_/X _12821_/X VGND VGND VPWR VPWR _12822_/X sky130_fd_sc_hd__or3_4
XANTENNA__15144__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24224__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16590_ _16554_/X _23666_/Q VGND VGND VPWR VPWR _16591_/C sky130_fd_sc_hd__or2_4
XFILLER_74_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22523__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15541_ _14431_/A _15541_/B _15541_/C VGND VGND VPWR VPWR _15541_/X sky130_fd_sc_hd__and3_4
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _12752_/X VGND VGND VPWR VPWR _12753_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14983__A _14983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _16047_/A VGND VGND VPWR VPWR _11704_/X sky130_fd_sc_hd__buf_2
X_18260_ _18314_/A _18257_/Y _18258_/Y _18260_/D VGND VGND VPWR VPWR _18261_/A sky130_fd_sc_hd__or4_4
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _12587_/A _15470_/X _15471_/X VGND VGND VPWR VPWR _15472_/X sky130_fd_sc_hd__and3_4
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12423_/X _12683_/X VGND VGND VPWR VPWR _12684_/X sky130_fd_sc_hd__or2_4
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17950__A1 _17875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17539_/A _17192_/X _14262_/X _17193_/X VGND VGND VPWR VPWR _17211_/X sky130_fd_sc_hd__o22a_4
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14418_/X _14420_/X _14423_/C VGND VGND VPWR VPWR _14423_/X sky130_fd_sc_hd__and3_4
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18191_ _23030_/B _18190_/X _23030_/B _18190_/X VGND VGND VPWR VPWR _19400_/A sky130_fd_sc_hd__a2bb2o_4
X_11635_ _11635_/A _11634_/X VGND VGND VPWR VPWR _11636_/A sky130_fd_sc_hd__or2_4
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11578__A1 _24464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17142_ _17114_/X _17138_/X _17124_/X _17141_/X VGND VGND VPWR VPWR _17142_/X sky130_fd_sc_hd__o22a_4
XFILLER_129_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14354_ _14366_/A _24028_/Q VGND VGND VPWR VPWR _14356_/B sky130_fd_sc_hd__or2_4
XFILLER_156_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _24446_/Q IRQ[9] _11565_/X VGND VGND VPWR VPWR _11566_/X sky130_fd_sc_hd__a21o_4
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22705__A _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13305_ _13290_/A _13305_/B _13305_/C VGND VGND VPWR VPWR _13306_/C sky130_fd_sc_hd__and3_4
Xclkbuf_7_31_0_HCLK clkbuf_7_31_0_HCLK/A VGND VGND VPWR VPWR _23409_/CLK sky130_fd_sc_hd__clkbuf_1
X_17073_ _17198_/A VGND VGND VPWR VPWR _17146_/A sky130_fd_sc_hd__buf_2
X_14285_ _14307_/A _14366_/B VGND VGND VPWR VPWR _14288_/B sky130_fd_sc_hd__or2_4
XANTENNA__12008__A _12106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16703__A _16592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_94_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR _23515_/CLK sky130_fd_sc_hd__clkbuf_1
X_16024_ _16062_/A _23758_/Q VGND VGND VPWR VPWR _16024_/X sky130_fd_sc_hd__or2_4
X_13236_ _13258_/A _13232_/X _13236_/C VGND VGND VPWR VPWR _13236_/X sky130_fd_sc_hd__or3_4
XFILLER_108_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20225__A _20396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21262__B2 _21252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11847__A _16635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13167_ _13306_/A _13163_/X _13167_/C VGND VGND VPWR VPWR _13167_/X sky130_fd_sc_hd__or3_4
XFILLER_124_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14223__A _11674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12118_ _16079_/A VGND VGND VPWR VPWR _12127_/A sky130_fd_sc_hd__buf_2
XFILLER_111_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13098_ _13085_/A _24072_/Q VGND VGND VPWR VPWR _13099_/C sky130_fd_sc_hd__or2_4
XANTENNA__22440__A _22440_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17975_ _17974_/X VGND VGND VPWR VPWR _17975_/X sky130_fd_sc_hd__buf_2
Xclkbuf_3_0_0_HCLK clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19714_ _19683_/B _19712_/X _19899_/A VGND VGND VPWR VPWR _19714_/X sky130_fd_sc_hd__a21o_4
X_16926_ _11645_/X _16926_/B _16926_/C VGND VGND VPWR VPWR _16931_/A sky130_fd_sc_hd__or3_4
X_12049_ _16595_/A VGND VGND VPWR VPWR _16725_/A sky130_fd_sc_hd__buf_2
XFILLER_66_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19645_ _19622_/X _19642_/Y _19644_/Y _19890_/B VGND VGND VPWR VPWR _19646_/B sky130_fd_sc_hd__o22a_4
X_16857_ _16855_/Y _16857_/B VGND VGND VPWR VPWR _16857_/X sky130_fd_sc_hd__or2_4
XANTENNA__12678__A _12677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11582__A _24465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15808_ _12536_/A _15808_/B _15808_/C VGND VGND VPWR VPWR _15809_/C sky130_fd_sc_hd__and3_4
XFILLER_81_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16788_ _16788_/A _23921_/Q VGND VGND VPWR VPWR _16790_/B sky130_fd_sc_hd__or2_4
X_19576_ _19889_/A VGND VGND VPWR VPWR _19576_/X sky130_fd_sc_hd__buf_2
XFILLER_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20895__A _20895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22514__B2 _22512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15739_ _11701_/A _15737_/X _15738_/X VGND VGND VPWR VPWR _15739_/X sky130_fd_sc_hd__and3_4
X_18527_ _18064_/X VGND VGND VPWR VPWR _18527_/X sky130_fd_sc_hd__buf_2
XANTENNA__14893__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18458_ _18405_/A _18415_/B VGND VGND VPWR VPWR _18458_/X sky130_fd_sc_hd__or2_4
XFILLER_166_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17409_ _17153_/Y _17410_/A VGND VGND VPWR VPWR _17412_/A sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_3_5_0_HCLK_A clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15501__B _15501_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18389_ _18389_/A _18388_/Y VGND VGND VPWR VPWR _18389_/X sky130_fd_sc_hd__and2_4
XANTENNA__13302__A _13276_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20420_ _20895_/A VGND VGND VPWR VPWR _20420_/X sky130_fd_sc_hd__buf_2
XANTENNA__24172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22615__A _22608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20351_ _20344_/X _20350_/X _24370_/Q _20269_/X VGND VGND VPWR VPWR _20351_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16613__A _11762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23070_ _23080_/A _23070_/B _23069_/X VGND VGND VPWR VPWR _23070_/X sky130_fd_sc_hd__and3_4
X_20282_ _20282_/A VGND VGND VPWR VPWR _20282_/X sky130_fd_sc_hd__buf_2
X_22021_ _22007_/A VGND VGND VPWR VPWR _22021_/X sky130_fd_sc_hd__buf_2
XANTENNA__11757__A _13392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21253__B2 _21252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21005__A1 _20894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21005__B2 _20396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23972_ _23908_/CLK _23972_/D VGND VGND VPWR VPWR _15688_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24247__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22923_ _18628_/X _18718_/X _18627_/X VGND VGND VPWR VPWR _22924_/C sky130_fd_sc_hd__o21a_4
XANTENNA__12588__A _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22854_ _15117_/Y _22848_/X _22849_/X VGND VGND VPWR VPWR _22854_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21308__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15899__A _13543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21805_ _21805_/A VGND VGND VPWR VPWR _21805_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22785_ _22784_/Y _22786_/B VGND VGND VPWR VPWR _22787_/A sky130_fd_sc_hd__nand2_4
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21736_ _21568_/X _21734_/X _15803_/B _21731_/X VGND VGND VPWR VPWR _21736_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24455_ _23347_/CLK _18808_/X HRESETn VGND VGND VPWR VPWR _11573_/A sky130_fd_sc_hd__dfrtp_4
X_21667_ _21667_/A VGND VGND VPWR VPWR _21667_/X sky130_fd_sc_hd__buf_2
XANTENNA__14308__A _12485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23406_ _23438_/CLK _23406_/D VGND VGND VPWR VPWR _23406_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20618_ _24453_/Q VGND VGND VPWR VPWR _20619_/A sky130_fd_sc_hd__inv_2
X_24386_ _24388_/CLK _24386_/D HRESETn VGND VGND VPWR VPWR _24386_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21598_ _21313_/A VGND VGND VPWR VPWR _21598_/X sky130_fd_sc_hd__buf_2
XFILLER_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20295__A2 _20252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23337_ _23337_/CLK _22333_/X VGND VGND VPWR VPWR _23337_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_18_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20549_ _20264_/X VGND VGND VPWR VPWR _20549_/X sky130_fd_sc_hd__buf_2
XANTENNA__16523__A _16452_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14070_ _11735_/A VGND VGND VPWR VPWR _14073_/A sky130_fd_sc_hd__buf_2
X_23268_ _23203_/CLK _23268_/D VGND VGND VPWR VPWR _15657_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13021_ _12499_/A _23624_/Q VGND VGND VPWR VPWR _13021_/X sky130_fd_sc_hd__or2_4
XANTENNA__11667__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22219_ _22165_/X _22215_/X _15166_/B _22184_/A VGND VGND VPWR VPWR _22219_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15139__A _14267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23199_ _23229_/CLK _23199_/D VGND VGND VPWR VPWR _23199_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_156_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14978__A _14771_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13882__A _13882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17760_ _17736_/A _17760_/B _17760_/C VGND VGND VPWR VPWR _17760_/X sky130_fd_sc_hd__and3_4
X_14972_ _14769_/A _14968_/X _14971_/X VGND VGND VPWR VPWR _14972_/X sky130_fd_sc_hd__or3_4
XANTENNA__13485__A1 _11858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21547__A2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13485__B2 _13484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13923_ _13923_/A _13923_/B _13923_/C VGND VGND VPWR VPWR _13927_/B sky130_fd_sc_hd__and3_4
X_16711_ _16711_/A _23953_/Q VGND VGND VPWR VPWR _16711_/X sky130_fd_sc_hd__or2_4
X_17691_ _17691_/A _17690_/Y VGND VGND VPWR VPWR _17697_/A sky130_fd_sc_hd__or2_4
X_16642_ _16682_/A _16642_/B _16641_/X VGND VGND VPWR VPWR _16642_/X sky130_fd_sc_hd__or3_4
X_19430_ _19428_/X _18682_/X _19428_/X _24217_/Q VGND VGND VPWR VPWR _24217_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13854_ _13628_/A _13929_/B VGND VGND VPWR VPWR _13856_/B sky130_fd_sc_hd__or2_4
XFILLER_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12805_ _13349_/A _12803_/X _12804_/X VGND VGND VPWR VPWR _12805_/X sky130_fd_sc_hd__and3_4
XANTENNA__23091__A _16901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16573_ _16588_/A _16573_/B _16572_/X VGND VGND VPWR VPWR _16577_/B sky130_fd_sc_hd__and3_4
X_19361_ _19358_/X _18474_/X _19358_/X _20713_/A VGND VGND VPWR VPWR _24258_/D sky130_fd_sc_hd__a2bb2o_4
X_13785_ _13782_/X _13785_/B VGND VGND VPWR VPWR _15391_/A sky130_fd_sc_hd__or2_4
XFILLER_76_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15524_ _12300_/A _15522_/X _15524_/C VGND VGND VPWR VPWR _15524_/X sky130_fd_sc_hd__and3_4
X_18312_ _18377_/A _17524_/X VGND VGND VPWR VPWR _18312_/Y sky130_fd_sc_hd__nor2_4
X_12736_ _12747_/A VGND VGND VPWR VPWR _13304_/A sky130_fd_sc_hd__buf_2
X_19292_ _19240_/A _19240_/B _19291_/Y VGND VGND VPWR VPWR _24291_/D sky130_fd_sc_hd__o21a_4
XFILLER_30_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18243_ _18215_/X _18239_/X _18240_/X _18242_/X VGND VGND VPWR VPWR _18243_/X sky130_fd_sc_hd__o22a_4
X_15455_ _15487_/A _15455_/B VGND VGND VPWR VPWR _15456_/C sky130_fd_sc_hd__or2_4
X_12667_ _12945_/A _12667_/B _12666_/X VGND VGND VPWR VPWR _12667_/X sky130_fd_sc_hd__or3_4
XFILLER_129_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13122__A _13100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14406_ _15486_/A _14406_/B VGND VGND VPWR VPWR _14406_/X sky130_fd_sc_hd__or2_4
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18174_ _18095_/X _17485_/X _18167_/X _18168_/X _18173_/Y VGND VGND VPWR VPWR _18175_/B
+ sky130_fd_sc_hd__a32o_4
X_11618_ _11618_/A VGND VGND VPWR VPWR _11877_/A sky130_fd_sc_hd__buf_2
X_15386_ _15121_/X _15385_/X _15384_/A _15382_/X VGND VGND VPWR VPWR _15386_/X sky130_fd_sc_hd__o22a_4
X_12598_ _12925_/A VGND VGND VPWR VPWR _12651_/A sky130_fd_sc_hd__buf_2
XFILLER_129_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22435__A _20530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17125_ _17124_/X VGND VGND VPWR VPWR _17817_/A sky130_fd_sc_hd__buf_2
XFILLER_156_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14337_ _14516_/A _14337_/B VGND VGND VPWR VPWR _14340_/B sky130_fd_sc_hd__or2_4
XANTENNA__21483__B2 _21482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22680__B1 _14590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17529__A _17515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11549_ _11549_/A _11549_/B VGND VGND VPWR VPWR _11549_/X sky130_fd_sc_hd__or2_4
XANTENNA__12961__A _12659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17056_ _17015_/X _17054_/B VGND VGND VPWR VPWR _17057_/B sky130_fd_sc_hd__and2_4
X_14268_ _14278_/A _14337_/B VGND VGND VPWR VPWR _14271_/B sky130_fd_sc_hd__or2_4
X_16007_ _13441_/A VGND VGND VPWR VPWR _16007_/X sky130_fd_sc_hd__buf_2
XFILLER_143_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13219_ _13258_/A _13214_/X _13218_/X VGND VGND VPWR VPWR _13219_/X sky130_fd_sc_hd__or3_4
XANTENNA__15049__A _14771_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14199_ _14199_/A _24031_/Q VGND VGND VPWR VPWR _14199_/X sky130_fd_sc_hd__or2_4
XFILLER_170_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21786__A2 _21784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13792__A _13792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17958_ _16943_/X _17910_/X _17014_/X _17957_/X VGND VGND VPWR VPWR _17958_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21538__A2 _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22735__B2 _22698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16909_ _16532_/Y _16908_/X _16824_/X _16906_/B VGND VGND VPWR VPWR _16910_/A sky130_fd_sc_hd__a211o_4
X_17889_ _17095_/X VGND VGND VPWR VPWR _18409_/A sky130_fd_sc_hd__buf_2
XFILLER_39_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19628_ _19690_/B _19628_/B VGND VGND VPWR VPWR _19634_/C sky130_fd_sc_hd__nor2_4
XFILLER_0_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12201__A _11881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19559_ _19510_/X _19558_/X VGND VGND VPWR VPWR _19559_/Y sky130_fd_sc_hd__nand2_4
XFILLER_146_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15512__A _12626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22570_ _22456_/X _22565_/X _23201_/Q _22569_/X VGND VGND VPWR VPWR _23201_/D sky130_fd_sc_hd__o22a_4
XFILLER_90_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21521_ _21134_/A _21370_/B _21320_/C _21184_/D VGND VGND VPWR VPWR _21521_/X sky130_fd_sc_hd__or4_4
XFILLER_142_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19919__A _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17390__A2 _17020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14128__A _14110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13032__A _12510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24240_ _24240_/CLK _19393_/X HRESETn VGND VGND VPWR VPWR _24240_/Q sky130_fd_sc_hd__dfrtp_4
X_21452_ _21438_/A VGND VGND VPWR VPWR _21452_/X sky130_fd_sc_hd__buf_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20403_ _18891_/X _20400_/Y _20402_/X _18983_/Y _20275_/X VGND VGND VPWR VPWR _20404_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21383_ _21254_/X _21377_/X _16304_/B _21381_/X VGND VGND VPWR VPWR _21383_/X sky130_fd_sc_hd__o22a_4
X_24171_ _23383_/CLK _24171_/D HRESETn VGND VGND VPWR VPWR _24171_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17439__A _17153_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22671__B1 _23136_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12871__A _12871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23122_ _23922_/CLK _22696_/X VGND VGND VPWR VPWR _23122_/Q sky130_fd_sc_hd__dfxtp_4
X_20334_ _20334_/A _20334_/B VGND VGND VPWR VPWR _20334_/X sky130_fd_sc_hd__or2_4
XANTENNA__12590__B _23371_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20265_ _20264_/X VGND VGND VPWR VPWR _20352_/A sky130_fd_sc_hd__buf_2
X_23053_ _23053_/A VGND VGND VPWR VPWR HADDR[25] sky130_fd_sc_hd__inv_2
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22004_ _21826_/X _22003_/X _15940_/B _22000_/X VGND VGND VPWR VPWR _22004_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20196_ _20196_/A _20195_/X VGND VGND VPWR VPWR _20196_/X sky130_fd_sc_hd__or2_4
XFILLER_163_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20985__B1 _20598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23637__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23955_ _23764_/CLK _21246_/X VGND VGND VPWR VPWR _23955_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_9_0_HCLK clkbuf_5_8_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22906_ _22742_/A _19319_/X _22738_/A _19910_/X VGND VGND VPWR VPWR _22906_/X sky130_fd_sc_hd__or4_4
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23886_ _23438_/CLK _21385_/X VGND VGND VPWR VPWR _16010_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21424__A _21431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22837_ _20700_/A _17284_/Y VGND VGND VPWR VPWR _22837_/X sky130_fd_sc_hd__or2_4
XFILLER_32_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16518__A _16370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11950__A _16116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15422__A _12477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19408__A1_N _19396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _13570_/A VGND VGND VPWR VPWR _13570_/Y sky130_fd_sc_hd__inv_2
X_22768_ _22759_/X _22761_/X _22768_/C _22768_/D VGND VGND VPWR VPWR _22769_/D sky130_fd_sc_hd__or4_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _12506_/A _23467_/Q VGND VGND VPWR VPWR _12522_/C sky130_fd_sc_hd__or2_4
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21719_ _21539_/X _21713_/X _16338_/B _21717_/X VGND VGND VPWR VPWR _21719_/X sky130_fd_sc_hd__o22a_4
XFILLER_13_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22699_ _21821_/A _22694_/X _16442_/B _22698_/X VGND VGND VPWR VPWR _23120_/D sky130_fd_sc_hd__o22a_4
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20982__B HRDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15240_ _14615_/A _15236_/X _15240_/C VGND VGND VPWR VPWR _15240_/X sky130_fd_sc_hd__or3_4
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12452_ _15017_/A VGND VGND VPWR VPWR _12453_/A sky130_fd_sc_hd__buf_2
X_24438_ _24419_/CLK _24438_/D HRESETn VGND VGND VPWR VPWR _24438_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22255__A _22226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15171_ _14297_/A _15169_/X _15170_/X VGND VGND VPWR VPWR _15175_/B sky130_fd_sc_hd__and3_4
XANTENNA__21465__B2 _21459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13877__A _13877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12383_ _12829_/A _23980_/Q VGND VGND VPWR VPWR _12384_/C sky130_fd_sc_hd__or2_4
X_24369_ _24397_/CLK _24369_/D HRESETn VGND VGND VPWR VPWR _24369_/Q sky130_fd_sc_hd__dfstp_4
X_14122_ _14149_/A _14117_/X _14121_/X VGND VGND VPWR VPWR _14122_/X sky130_fd_sc_hd__and3_4
XFILLER_125_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21217__B2 _21216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18930_ _14261_/A _18927_/X _19078_/A _18928_/X VGND VGND VPWR VPWR _18930_/X sky130_fd_sc_hd__o22a_4
X_14053_ _13705_/A _23968_/Q VGND VGND VPWR VPWR _14053_/X sky130_fd_sc_hd__or2_4
XFILLER_4_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13004_ _12493_/A _13004_/B _13004_/C VGND VGND VPWR VPWR _13008_/B sky130_fd_sc_hd__and3_4
XANTENNA__21768__A2 _21763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18861_ _13262_/X _18856_/X _20579_/A _18857_/X VGND VGND VPWR VPWR _24423_/D sky130_fd_sc_hd__o22a_4
X_17812_ _17878_/A VGND VGND VPWR VPWR _17812_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18792_ _12180_/X _18787_/X _24467_/Q _18790_/X VGND VGND VPWR VPWR _24467_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22717__B2 _22712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17743_ _17743_/A _17298_/X VGND VGND VPWR VPWR _17743_/X sky130_fd_sc_hd__or2_4
X_14955_ _14967_/A _14884_/B VGND VGND VPWR VPWR _14955_/X sky130_fd_sc_hd__or2_4
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22193__A2 _22187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13906_ _14385_/A _13904_/X _13906_/C VGND VGND VPWR VPWR _13910_/B sky130_fd_sc_hd__and3_4
X_17674_ _17667_/A _17576_/Y _17668_/Y VGND VGND VPWR VPWR _18013_/B sky130_fd_sc_hd__a21o_4
X_14886_ _14133_/A _14882_/X _14885_/X VGND VGND VPWR VPWR _14886_/X sky130_fd_sc_hd__or3_4
XANTENNA__12021__A _12020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21334__A _21341_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19413_ _19411_/X _18372_/X _19411_/X _24229_/Q VGND VGND VPWR VPWR _19413_/X sky130_fd_sc_hd__a2bb2o_4
X_16625_ _11772_/X VGND VGND VPWR VPWR _16639_/A sky130_fd_sc_hd__buf_2
X_13837_ _15405_/A _13837_/B _13837_/C VGND VGND VPWR VPWR _13837_/X sky130_fd_sc_hd__or3_4
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12956__A _12949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11860__A _14012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19344_ _19340_/X _18104_/X _19343_/X _20436_/A VGND VGND VPWR VPWR _24270_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16556_ _16556_/A _16556_/B _16556_/C VGND VGND VPWR VPWR _16561_/B sky130_fd_sc_hd__and3_4
XANTENNA__21153__B1 _12632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13768_ _12623_/A _13768_/B VGND VGND VPWR VPWR _13768_/X sky130_fd_sc_hd__or2_4
XFILLER_149_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15507_ _12630_/A _15503_/X _15506_/X VGND VGND VPWR VPWR _15507_/X sky130_fd_sc_hd__or3_4
X_12719_ _12279_/A VGND VGND VPWR VPWR _12722_/A sky130_fd_sc_hd__buf_2
XANTENNA__15051__B _23509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16487_ _16362_/X _16483_/X _16487_/C VGND VGND VPWR VPWR _16487_/X sky130_fd_sc_hd__or3_4
X_19275_ _19248_/X VGND VGND VPWR VPWR _19275_/Y sky130_fd_sc_hd__inv_2
X_13699_ _13699_/A VGND VGND VPWR VPWR _13700_/A sky130_fd_sc_hd__buf_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15438_ _13677_/A _15438_/B _15438_/C VGND VGND VPWR VPWR _15442_/B sky130_fd_sc_hd__and3_4
X_18226_ _18225_/X VGND VGND VPWR VPWR _18226_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15383__A1 _15382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24345__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13787__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15369_ _15369_/A _15365_/X _15369_/C VGND VGND VPWR VPWR _15369_/X sky130_fd_sc_hd__or3_4
X_18157_ _17976_/X _18128_/X _17883_/X VGND VGND VPWR VPWR _18157_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21456__B2 _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16163__A _13413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24092__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17108_ _17107_/X VGND VGND VPWR VPWR _17108_/X sky130_fd_sc_hd__buf_2
X_18088_ _18088_/A VGND VGND VPWR VPWR _18637_/B sky130_fd_sc_hd__inv_2
XFILLER_171_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21208__B2 _21202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17039_ _17039_/A VGND VGND VPWR VPWR _17039_/X sky130_fd_sc_hd__buf_2
XFILLER_131_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20050_ _20050_/A VGND VGND VPWR VPWR _20050_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20967__B1 _20262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20413__A _20334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14411__A _11813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15226__B _15162_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14130__B _23167_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19585__B1 HRDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23740_ _23772_/CLK _23740_/D VGND VGND VPWR VPWR _14345_/B sky130_fd_sc_hd__dfxtp_4
X_20952_ _21017_/A _20951_/X VGND VGND VPWR VPWR _20952_/Y sky130_fd_sc_hd__nor2_4
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21931__A2 _21930_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21244__A _21238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ _23671_/CLK _23671_/D VGND VGND VPWR VPWR _15139_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12866__A _12866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20883_ _20781_/X _20882_/X _19136_/A _20791_/X VGND VGND VPWR VPWR _20883_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22622_ _22622_/A VGND VGND VPWR VPWR _22622_/X sky130_fd_sc_hd__buf_2
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20498__A2 _20497_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22553_ _22428_/X _22551_/X _16177_/B _22548_/X VGND VGND VPWR VPWR _22553_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22892__B1 _17353_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21504_ _21287_/X _21499_/X _15574_/B _21503_/X VGND VGND VPWR VPWR _23809_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15896__B _15840_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22484_ _22169_/A VGND VGND VPWR VPWR _22484_/X sky130_fd_sc_hd__buf_2
XFILLER_10_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13697__A _13697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24223_ _24248_/CLK _24223_/D HRESETn VGND VGND VPWR VPWR _24223_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21447__B2 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21435_ _21256_/X _21434_/X _15989_/B _21431_/X VGND VGND VPWR VPWR _23854_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17169__A _15517_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16073__A _16049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21998__A2 _21996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24154_ _24302_/CLK _24154_/D HRESETn VGND VGND VPWR VPWR _17702_/A sky130_fd_sc_hd__dfrtp_4
X_21366_ _21311_/X _21362_/X _15155_/B _21331_/A VGND VGND VPWR VPWR _23895_/D sky130_fd_sc_hd__o22a_4
X_23105_ _23744_/CLK _23105_/D VGND VGND VPWR VPWR _15634_/B sky130_fd_sc_hd__dfxtp_4
X_20317_ _20316_/X VGND VGND VPWR VPWR _20318_/B sky130_fd_sc_hd__buf_2
X_24085_ _23617_/CLK _21025_/X VGND VGND VPWR VPWR _24085_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12106__A _12106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21297_ _20841_/A VGND VGND VPWR VPWR _21297_/X sky130_fd_sc_hd__buf_2
XFILLER_162_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23036_ _22908_/A VGND VGND VPWR VPWR _23036_/X sky130_fd_sc_hd__buf_2
X_20248_ _20244_/X _20248_/B VGND VGND VPWR VPWR _20249_/A sky130_fd_sc_hd__or2_4
XFILLER_88_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20323__A _20270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15417__A _14329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20179_ _24456_/Q IRQ[19] _20178_/X VGND VGND VPWR VPWR _20179_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__14321__A _12191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11664__B _15377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_HCLK_A clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14740_ _12503_/A _24057_/Q VGND VGND VPWR VPWR _14741_/C sky130_fd_sc_hd__or2_4
X_23938_ _23587_/CLK _23938_/D VGND VGND VPWR VPWR _15470_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11952_ _11975_/A VGND VGND VPWR VPWR _12102_/A sky130_fd_sc_hd__buf_2
XFILLER_44_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21922__A2 _21916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14671_ _14685_/A _14668_/X _14671_/C VGND VGND VPWR VPWR _14672_/C sky130_fd_sc_hd__and3_4
X_11883_ _11882_/X VGND VGND VPWR VPWR _16155_/A sky130_fd_sc_hd__buf_2
X_23869_ _23101_/CLK _21408_/X VGND VGND VPWR VPWR _13933_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12776__A _12773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16410_ _16094_/A _16408_/X _16409_/X VGND VGND VPWR VPWR _16411_/C sky130_fd_sc_hd__and3_4
XANTENNA__11680__A _11680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15152__A _15022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13622_ _13622_/A VGND VGND VPWR VPWR _15404_/A sky130_fd_sc_hd__buf_2
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17390_ _15915_/Y _17020_/X _17028_/X _17389_/X VGND VGND VPWR VPWR _17448_/B sky130_fd_sc_hd__o22a_4
XFILLER_38_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16341_ _16333_/A _16266_/B VGND VGND VPWR VPWR _16341_/X sky130_fd_sc_hd__or2_4
X_13553_ _13515_/X _23717_/Q VGND VGND VPWR VPWR _13555_/B sky130_fd_sc_hd__or2_4
XANTENNA__21686__B2 _21681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14991__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12504_ _12504_/A VGND VGND VPWR VPWR _12540_/A sky130_fd_sc_hd__buf_2
X_19060_ _24386_/Q VGND VGND VPWR VPWR _19060_/Y sky130_fd_sc_hd__inv_2
X_16272_ _11917_/X _16270_/X _16272_/C VGND VGND VPWR VPWR _16272_/X sky130_fd_sc_hd__and3_4
X_13484_ _11971_/X _13461_/X _13468_/X _13475_/X _13483_/X VGND VGND VPWR VPWR _13484_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_160_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15223_ _15198_/X _15223_/B VGND VGND VPWR VPWR _15224_/C sky130_fd_sc_hd__or2_4
X_18011_ _17967_/X _17973_/Y _18000_/X _18007_/X _18010_/Y VGND VGND VPWR VPWR _18011_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_145_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12435_ _12435_/A VGND VGND VPWR VPWR _12852_/A sky130_fd_sc_hd__buf_2
XFILLER_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15154_ _13586_/A _15128_/X _15138_/X _15145_/X _15153_/X VGND VGND VPWR VPWR _15154_/X
+ sky130_fd_sc_hd__a32o_4
X_12366_ _15887_/A _12359_/X _12365_/X VGND VGND VPWR VPWR _12366_/X sky130_fd_sc_hd__or3_4
XFILLER_5_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14105_ _11898_/A _23295_/Q VGND VGND VPWR VPWR _14105_/X sky130_fd_sc_hd__or2_4
X_19962_ _18150_/A _19962_/B VGND VGND VPWR VPWR _19962_/X sky130_fd_sc_hd__or2_4
X_15085_ _12322_/A _23893_/Q VGND VGND VPWR VPWR _15085_/X sky130_fd_sc_hd__or2_4
X_12297_ _13145_/A _24108_/Q VGND VGND VPWR VPWR _12297_/X sky130_fd_sc_hd__or2_4
XANTENNA__12016__A _12001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18913_ _18897_/A VGND VGND VPWR VPWR _18913_/X sky130_fd_sc_hd__buf_2
XFILLER_84_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14036_ _14056_/A _23584_/Q VGND VGND VPWR VPWR _14037_/C sky130_fd_sc_hd__or2_4
X_19893_ _19749_/X _19752_/D _19763_/Y VGND VGND VPWR VPWR _19903_/B sky130_fd_sc_hd__o21ai_4
XFILLER_136_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11855__A _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18844_ _11851_/X _18840_/X _24436_/Q _18843_/X VGND VGND VPWR VPWR _18844_/X sky130_fd_sc_hd__o22a_4
XFILLER_132_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18775_ _17013_/X _18774_/X _17751_/A _16943_/X VGND VGND VPWR VPWR _18775_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15987_ _16003_/A _15983_/X _15987_/C VGND VGND VPWR VPWR _15987_/X sky130_fd_sc_hd__or3_4
XANTENNA__22166__A2 _22159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17726_ _17726_/A _17407_/X VGND VGND VPWR VPWR _17730_/B sky130_fd_sc_hd__and2_4
XFILLER_76_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14938_ _12327_/A VGND VGND VPWR VPWR _14970_/A sky130_fd_sc_hd__buf_2
XFILLER_94_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17657_ _17780_/A _17263_/Y VGND VGND VPWR VPWR _17657_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12686__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14869_ _14114_/A _14867_/X _14868_/X VGND VGND VPWR VPWR _14869_/X sky130_fd_sc_hd__and3_4
XFILLER_1_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11590__A _17060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16608_ _16608_/A VGND VGND VPWR VPWR _16621_/A sky130_fd_sc_hd__buf_2
X_17588_ _16381_/X _17561_/B VGND VGND VPWR VPWR _17588_/Y sky130_fd_sc_hd__nand2_4
XFILLER_143_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19327_ _19327_/A VGND VGND VPWR VPWR _19327_/Y sky130_fd_sc_hd__inv_2
X_16539_ _12015_/A VGND VGND VPWR VPWR _16539_/X sky130_fd_sc_hd__buf_2
XFILLER_143_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18373__A _18032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20885__C1 _20884_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19258_ _19258_/A VGND VGND VPWR VPWR _19258_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20408__A _20313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18209_ _17490_/D _18207_/X _18060_/X VGND VGND VPWR VPWR _18209_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__22096__A2_N _22094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21429__B2 _21424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19189_ _19148_/B VGND VGND VPWR VPWR _19189_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20127__B _20126_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21220_ _20801_/X _21219_/X _23967_/Q _21216_/X VGND VGND VPWR VPWR _23967_/D sky130_fd_sc_hd__o22a_4
XFILLER_144_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21151_ _20486_/X _21148_/X _24012_/Q _21145_/X VGND VGND VPWR VPWR _21151_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20102_ _20150_/A _20100_/X _20101_/Y _19959_/A VGND VGND VPWR VPWR _20102_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21239__A _21264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21082_ _22637_/D VGND VGND VPWR VPWR _22487_/B sky130_fd_sc_hd__buf_2
XANTENNA__13964__B _23296_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20033_ _18275_/X _20031_/X _20032_/Y _20018_/X VGND VGND VPWR VPWR _20033_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11765__A _11762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19932__A _22745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15237__A _14677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14141__A _11898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21601__B2 _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20955__A3 _20953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17281__A1 _14483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22157__A2 _22147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13980__A _11930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21984_ _21879_/X _21981_/X _15343_/B _21978_/X VGND VGND VPWR VPWR _23544_/D sky130_fd_sc_hd__o22a_4
XFILLER_66_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21904__A2 _21902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23723_ _23723_/CLK _23723_/D VGND VGND VPWR VPWR _12664_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20935_ _20935_/A _20934_/X VGND VGND VPWR VPWR _20935_/X sky130_fd_sc_hd__or2_4
XANTENNA__12596__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16068__A _16222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _23397_/CLK _21782_/X VGND VGND VPWR VPWR _23654_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21117__B1 _24032_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _20940_/A _20866_/B VGND VGND VPWR VPWR _20866_/X sky130_fd_sc_hd__or2_4
XFILLER_148_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22605_ _22605_/A VGND VGND VPWR VPWR _22605_/X sky130_fd_sc_hd__buf_2
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21668__B2 _21667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23585_ _23617_/CLK _23585_/D VGND VGND VPWR VPWR _15602_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20797_ _24255_/Q _20661_/X _20796_/X VGND VGND VPWR VPWR _20797_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18283__A _18283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15700__A _13338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22536_ _11763_/B VGND VGND VPWR VPWR _22536_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22617__B1 _15868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22467_ _22466_/X _22462_/X _13796_/B _22457_/X VGND VGND VPWR VPWR _23261_/D sky130_fd_sc_hd__o22a_4
X_12220_ _12294_/A VGND VGND VPWR VPWR _13676_/A sky130_fd_sc_hd__buf_2
X_24206_ _24184_/CLK _19658_/X HRESETn VGND VGND VPWR VPWR _11611_/B sky130_fd_sc_hd__dfrtp_4
X_21418_ _21315_/X _21391_/A _15104_/B _21381_/A VGND VGND VPWR VPWR _23861_/D sky130_fd_sc_hd__o22a_4
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22398_ _22158_/X _22397_/X _14564_/B _22394_/X VGND VGND VPWR VPWR _22398_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24391__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21840__A1 _21838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24137_ _24137_/CLK _20107_/Y HRESETn VGND VGND VPWR VPWR _24137_/Q sky130_fd_sc_hd__dfrtp_4
X_12151_ _12151_/A _23635_/Q VGND VGND VPWR VPWR _12151_/X sky130_fd_sc_hd__or2_4
XANTENNA__21840__B2 _21834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21349_ _21280_/X _21348_/X _23908_/Q _21345_/X VGND VGND VPWR VPWR _21349_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23205__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24068_ _23908_/CLK _21060_/X VGND VGND VPWR VPWR _15756_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17346__B _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12082_ _12051_/A _23635_/Q VGND VGND VPWR VPWR _12084_/B sky130_fd_sc_hd__or2_4
XFILLER_104_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11675__A _11675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22396__A2 _22390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15910_ _13564_/A _15910_/B _15910_/C VGND VGND VPWR VPWR _15911_/C sky130_fd_sc_hd__and3_4
X_23019_ _23048_/A VGND VGND VPWR VPWR _23019_/X sky130_fd_sc_hd__buf_2
XANTENNA__15147__A _14170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14051__A _11812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16890_ _16246_/A _16889_/X _16246_/A _16889_/X VGND VGND VPWR VPWR _16890_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15841_ _12487_/A _15841_/B VGND VGND VPWR VPWR _15842_/C sky130_fd_sc_hd__or2_4
XFILLER_134_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14986__A _14170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22148__A2 _22147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17362__A _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13890__A _13877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18560_ _17436_/B _18560_/B VGND VGND VPWR VPWR _18560_/Y sky130_fd_sc_hd__nand2_4
X_15772_ _11739_/A _15772_/B _15772_/C VGND VGND VPWR VPWR _15773_/C sky130_fd_sc_hd__and3_4
X_12984_ _12983_/X VGND VGND VPWR VPWR _12984_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17511_ _17493_/A _17511_/B VGND VGND VPWR VPWR _17511_/X sky130_fd_sc_hd__or2_4
X_11935_ _11935_/A VGND VGND VPWR VPWR _12904_/A sky130_fd_sc_hd__buf_2
X_14723_ _12190_/A _14723_/B VGND VGND VPWR VPWR _14723_/X sky130_fd_sc_hd__or2_4
XFILLER_91_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18491_ _17250_/X _18419_/X _17250_/X _18415_/C VGND VGND VPWR VPWR _18491_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17442_ _17435_/Y _17440_/X _17441_/X VGND VGND VPWR VPWR _17442_/X sky130_fd_sc_hd__o21a_4
X_14654_ _14684_/A _14568_/B VGND VGND VPWR VPWR _14655_/C sky130_fd_sc_hd__or2_4
X_11866_ _11865_/X VGND VGND VPWR VPWR _16160_/A sky130_fd_sc_hd__buf_2
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22708__A _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _12477_/A _13605_/B VGND VGND VPWR VPWR _13610_/B sky130_fd_sc_hd__or2_4
XPHY_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21612__A _21608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17373_ _17169_/X _17446_/B VGND VGND VPWR VPWR _17374_/A sky130_fd_sc_hd__or2_4
X_14585_ _14280_/A _14583_/X _14584_/X VGND VGND VPWR VPWR _14585_/X sky130_fd_sc_hd__and3_4
X_11797_ _12138_/A _11790_/X _11796_/X VGND VGND VPWR VPWR _11797_/X sky130_fd_sc_hd__or3_4
XANTENNA__22320__A2 _22315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19112_ _18987_/A _19110_/Y _19111_/Y _19106_/X VGND VGND VPWR VPWR _19112_/X sky130_fd_sc_hd__o22a_4
X_13536_ _13503_/X _13536_/B _13536_/C VGND VGND VPWR VPWR _13537_/C sky130_fd_sc_hd__and3_4
X_16324_ _16316_/A _16259_/B VGND VGND VPWR VPWR _16324_/X sky130_fd_sc_hd__or2_4
XFILLER_9_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20228__A _20216_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16255_ _16159_/A _16255_/B _16254_/X VGND VGND VPWR VPWR _16255_/X sky130_fd_sc_hd__or3_4
X_19043_ _24389_/Q VGND VGND VPWR VPWR _19043_/Y sky130_fd_sc_hd__inv_2
X_13467_ _13467_/A _13465_/X _13467_/C VGND VGND VPWR VPWR _13468_/C sky130_fd_sc_hd__and3_4
XFILLER_12_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13130__A _12696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15206_ _14677_/A _15149_/B VGND VGND VPWR VPWR _15208_/B sky130_fd_sc_hd__or2_4
XFILLER_51_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12418_ _13566_/A _12380_/X _12417_/X VGND VGND VPWR VPWR _12418_/X sky130_fd_sc_hd__and3_4
X_16186_ _16214_/A _16179_/X _16186_/C VGND VGND VPWR VPWR _16187_/C sky130_fd_sc_hd__or3_4
XANTENNA__22084__B2 _22078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13398_ _13398_/A _13396_/X _13398_/C VGND VGND VPWR VPWR _13399_/C sky130_fd_sc_hd__and3_4
XFILLER_114_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15137_ _15269_/A _15137_/B _15137_/C VGND VGND VPWR VPWR _15137_/X sky130_fd_sc_hd__and3_4
X_12349_ _11712_/X _24044_/Q VGND VGND VPWR VPWR _12349_/X sky130_fd_sc_hd__or2_4
XFILLER_47_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21059__A _21045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19945_ _19920_/X _24164_/Q _22745_/A _22737_/A VGND VGND VPWR VPWR _19945_/X sky130_fd_sc_hd__o22a_4
X_15068_ _15086_/A _23573_/Q VGND VGND VPWR VPWR _15069_/C sky130_fd_sc_hd__or2_4
XANTENNA__24130__CLK _24342_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15057__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14019_ _13877_/A _23520_/Q VGND VGND VPWR VPWR _14019_/X sky130_fd_sc_hd__or2_4
XFILLER_136_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19876_ _19665_/A _19875_/X VGND VGND VPWR VPWR _19876_/X sky130_fd_sc_hd__and2_4
XANTENNA__21595__B1 _23768_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18827_ _17290_/X _18824_/X _24442_/Q _18825_/X VGND VGND VPWR VPWR _18827_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14896__A _14114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17272__A _14412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24280__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18758_ _18744_/A _17346_/B VGND VGND VPWR VPWR _18758_/X sky130_fd_sc_hd__and2_4
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17709_ _16983_/A _17389_/X VGND VGND VPWR VPWR _17710_/B sky130_fd_sc_hd__or2_4
XANTENNA__23848__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21898__B2 _21892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18689_ _18689_/A _18687_/Y VGND VGND VPWR VPWR _18689_/Y sky130_fd_sc_hd__nand2_4
XFILLER_63_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18763__A1 _12021_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20720_ _20635_/X _20719_/X _15509_/B _20614_/X VGND VGND VPWR VPWR _24098_/D sky130_fd_sc_hd__o22a_4
XFILLER_169_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20651_ _20515_/X _20650_/X _24324_/Q _20522_/X VGND VGND VPWR VPWR _20651_/X sky130_fd_sc_hd__o22a_4
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16616__A _11836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22311__A2 _22308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23370_ _23404_/CLK _22293_/X VGND VGND VPWR VPWR _12768_/B sky130_fd_sc_hd__dfxtp_4
X_20582_ _20447_/X _20579_/Y _20581_/X _19032_/Y _20495_/X VGND VGND VPWR VPWR _20583_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22321_ _22169_/X _22294_/A _23349_/Q _22284_/A VGND VGND VPWR VPWR _23349_/D sky130_fd_sc_hd__o22a_4
XFILLER_118_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14136__A _15281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22252_ _22134_/X _22251_/X _15762_/B _22248_/X VGND VGND VPWR VPWR _23396_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24401__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22075__B2 _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21203_ _20509_/X _21198_/X _23979_/Q _21202_/X VGND VGND VPWR VPWR _21203_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22183_ _22103_/X _22180_/X _16799_/B _22177_/X VGND VGND VPWR VPWR _23441_/D sky130_fd_sc_hd__o22a_4
XFILLER_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21134_ _21134_/A _21134_/B _21134_/C _21134_/D VGND VGND VPWR VPWR _21134_/X sky130_fd_sc_hd__or4_4
XFILLER_132_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22378__A2 _22376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23378__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21065_ _20770_/X _21059_/X _24064_/Q _21063_/X VGND VGND VPWR VPWR _24064_/D sky130_fd_sc_hd__o22a_4
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22800__B _18774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21050__A2 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20016_ _18670_/A VGND VGND VPWR VPWR _20016_/X sky130_fd_sc_hd__buf_2
XFILLER_101_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17182__A _12027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15414__B _15471_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21967_ _21960_/A VGND VGND VPWR VPWR _21967_/X sky130_fd_sc_hd__buf_2
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13215__A _12372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22550__A2 _22544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11720_ _11720_/A VGND VGND VPWR VPWR _13868_/A sky130_fd_sc_hd__buf_2
X_23706_ _23101_/CLK _23706_/D VGND VGND VPWR VPWR _14686_/B sky130_fd_sc_hd__dfxtp_4
X_20918_ _20867_/A _20364_/B VGND VGND VPWR VPWR _20918_/X sky130_fd_sc_hd__or2_4
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ _21819_/X _21895_/X _23601_/Q _21892_/X VGND VGND VPWR VPWR _23601_/D sky130_fd_sc_hd__o22a_4
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _15321_/A VGND VGND VPWR VPWR _13865_/A sky130_fd_sc_hd__buf_2
X_23637_ _23392_/CLK _21804_/X VGND VGND VPWR VPWR _23637_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20849_ _20703_/X _20848_/X _19094_/A _20647_/X VGND VGND VPWR VPWR _20849_/X sky130_fd_sc_hd__o22a_4
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22302__A2 _22301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15430__A _14319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14370_ _12583_/A _23548_/Q VGND VGND VPWR VPWR _14371_/C sky130_fd_sc_hd__or2_4
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23568_ _23533_/CLK _23568_/D VGND VGND VPWR VPWR _16409_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_126_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ _24465_/Q IRQ[28] VGND VGND VPWR VPWR _20188_/A sky130_fd_sc_hd__and2_4
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _13321_/A _13319_/X _13320_/X VGND VGND VPWR VPWR _13322_/C sky130_fd_sc_hd__and3_4
XFILLER_167_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22519_ _22505_/A VGND VGND VPWR VPWR _22519_/X sky130_fd_sc_hd__buf_2
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23499_ _24074_/CLK _22058_/X VGND VGND VPWR VPWR _12668_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14046__A _12581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16040_ _16056_/A _16038_/X _16039_/X VGND VGND VPWR VPWR _16040_/X sky130_fd_sc_hd__and3_4
XANTENNA__22066__A1 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13252_ _13252_/A _23495_/Q VGND VGND VPWR VPWR _13254_/B sky130_fd_sc_hd__or2_4
XANTENNA__22066__B2 _22064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24153__CLK _24302_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ _13042_/A VGND VGND VPWR VPWR _12693_/A sky130_fd_sc_hd__buf_2
XANTENNA__20616__A2 _22737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17357__A _17357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13885__A _13885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13183_ _13183_/A _23111_/Q VGND VGND VPWR VPWR _13185_/B sky130_fd_sc_hd__or2_4
XFILLER_163_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12134_ _12122_/A _12134_/B _12134_/C VGND VGND VPWR VPWR _12138_/B sky130_fd_sc_hd__and3_4
XFILLER_150_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17991_ _17991_/A VGND VGND VPWR VPWR _17991_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19730_ _19556_/X _19723_/X _19726_/Y _19729_/X VGND VGND VPWR VPWR _19730_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20214__C _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16942_ _16941_/X VGND VGND VPWR VPWR _16943_/A sky130_fd_sc_hd__buf_2
XANTENNA__19572__A HRDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12065_ _12064_/X _23571_/Q VGND VGND VPWR VPWR _12065_/X sky130_fd_sc_hd__or2_4
XFILLER_150_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21041__A2 _21038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19661_ _19661_/A _19665_/B VGND VGND VPWR VPWR _19662_/B sky130_fd_sc_hd__or2_4
XFILLER_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16873_ _16865_/X _16867_/X _16873_/C _16873_/D VGND VGND VPWR VPWR _16873_/X sky130_fd_sc_hd__or4_4
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18612_ _18565_/A _17307_/X _18608_/X _18611_/Y VGND VGND VPWR VPWR _18612_/X sky130_fd_sc_hd__a211o_4
X_15824_ _12440_/A _15824_/B _15823_/X VGND VGND VPWR VPWR _15824_/X sky130_fd_sc_hd__and3_4
X_19592_ _19750_/A VGND VGND VPWR VPWR _19724_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_54_0_HCLK clkbuf_6_27_0_HCLK/X VGND VGND VPWR VPWR _23404_/CLK sky130_fd_sc_hd__clkbuf_1
X_18543_ _18467_/X _18230_/Y _17869_/X _18542_/X VGND VGND VPWR VPWR _18543_/X sky130_fd_sc_hd__a211o_4
XFILLER_79_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12967_ _12943_/A _23881_/Q VGND VGND VPWR VPWR _12967_/X sky130_fd_sc_hd__or2_4
X_15755_ _15741_/X _15755_/B VGND VGND VPWR VPWR _15755_/X sky130_fd_sc_hd__or2_4
XFILLER_166_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13125__A _12979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11918_ _11917_/X VGND VGND VPWR VPWR _16123_/A sky130_fd_sc_hd__buf_2
X_14706_ _14295_/A _14774_/B VGND VGND VPWR VPWR _14706_/X sky130_fd_sc_hd__or2_4
XFILLER_73_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20552__A1 _18272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18474_ _17715_/X _17765_/X _17715_/X _17765_/X VGND VGND VPWR VPWR _18474_/X sky130_fd_sc_hd__a2bb2o_4
X_12898_ _12871_/A _23497_/Q VGND VGND VPWR VPWR _12900_/B sky130_fd_sc_hd__or2_4
X_15686_ _13339_/A _15663_/X _15670_/X _15677_/X _15685_/X VGND VGND VPWR VPWR _15686_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22438__A _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17425_ _14263_/A VGND VGND VPWR VPWR _17425_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11849_ _11686_/X _11849_/B _11848_/X VGND VGND VPWR VPWR _11850_/C sky130_fd_sc_hd__and3_4
X_14637_ _14677_/A VGND VGND VPWR VPWR _14653_/A sky130_fd_sc_hd__buf_2
XFILLER_92_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17356_ _17044_/B VGND VGND VPWR VPWR _17378_/A sky130_fd_sc_hd__inv_2
X_14568_ _13601_/A _14568_/B VGND VGND VPWR VPWR _14569_/C sky130_fd_sc_hd__or2_4
XFILLER_159_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16307_ _11865_/X _16306_/X VGND VGND VPWR VPWR _16307_/X sky130_fd_sc_hd__and2_4
X_13519_ _13562_/A _13516_/X _13518_/X VGND VGND VPWR VPWR _13520_/C sky130_fd_sc_hd__and3_4
X_14499_ _14506_/A _14499_/B VGND VGND VPWR VPWR _14499_/X sky130_fd_sc_hd__or2_4
X_17287_ _17284_/Y _17019_/X _17026_/X _17286_/X VGND VGND VPWR VPWR _17287_/X sky130_fd_sc_hd__o22a_4
XFILLER_174_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18651__A _18483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19026_ _24392_/Q VGND VGND VPWR VPWR _19026_/Y sky130_fd_sc_hd__inv_2
X_16238_ _11815_/X _16238_/B _16238_/C VGND VGND VPWR VPWR _16238_/X sky130_fd_sc_hd__or3_4
XFILLER_127_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13795__A _14574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17267__A _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16169_ _13398_/A VGND VGND VPWR VPWR _16220_/A sky130_fd_sc_hd__buf_2
XANTENNA__21804__B2 _21767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17484__A1 _17480_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24307__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17484__B2 _17483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19928_ _19921_/X _24177_/Q _19925_/X _20339_/B VGND VGND VPWR VPWR _24177_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12204__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19859_ _19859_/A _19859_/B VGND VGND VPWR VPWR _19859_/X sky130_fd_sc_hd__or2_4
XANTENNA__20421__A _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15515__A _11682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22870_ _17480_/Y _22846_/X _22799_/X _22869_/X VGND VGND VPWR VPWR _22870_/X sky130_fd_sc_hd__a211o_4
XFILLER_3_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21821_ _21821_/A VGND VGND VPWR VPWR _21821_/X sky130_fd_sc_hd__buf_2
XANTENNA__15234__B _15176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13035__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21752_ _21596_/X _21748_/X _15139_/B _21717_/A VGND VGND VPWR VPWR _23671_/D sky130_fd_sc_hd__o22a_4
XFILLER_52_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21252__A _21239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20703_ _20275_/X VGND VGND VPWR VPWR _20703_/X sky130_fd_sc_hd__buf_2
X_24471_ _24471_/CLK _24471_/D HRESETn VGND VGND VPWR VPWR _20154_/A sky130_fd_sc_hd__dfrtp_4
X_21683_ _21563_/X _21677_/X _23717_/Q _21681_/X VGND VGND VPWR VPWR _21683_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12874__A _12874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16346__A _13383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15250__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23422_ _23101_/CLK _23422_/D VGND VGND VPWR VPWR _13761_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21099__A2 _21097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20634_ _20533_/X _20633_/X _13470_/B _20614_/X VGND VGND VPWR VPWR _20634_/X sky130_fd_sc_hd__o22a_4
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22296__B2 _22291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12593__B _23755_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24176__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23353_ _23290_/CLK _22317_/X VGND VGND VPWR VPWR _14779_/B sky130_fd_sc_hd__dfxtp_4
X_20565_ _20425_/X _20564_/X _24296_/Q _20519_/X VGND VGND VPWR VPWR _20565_/X sky130_fd_sc_hd__o22a_4
XFILLER_149_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22304_ _22139_/X _22301_/X _15458_/B _22298_/X VGND VGND VPWR VPWR _23362_/D sky130_fd_sc_hd__o22a_4
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22048__B2 _22043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23284_ _23475_/CLK _22411_/X VGND VGND VPWR VPWR _11718_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20496_ _20447_/X _20491_/Y _20494_/X _19007_/Y _20495_/X VGND VGND VPWR VPWR _20497_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_69_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22599__A2 _22594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22235_ _22105_/X _22230_/X _16431_/B _22234_/X VGND VGND VPWR VPWR _23408_/D sky130_fd_sc_hd__o22a_4
XFILLER_106_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22166_ _22165_/X _22159_/X _15150_/B _22106_/A VGND VGND VPWR VPWR _23447_/D sky130_fd_sc_hd__o22a_4
XFILLER_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22811__A _14483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21117_ _20770_/X _21111_/X _24032_/Q _21115_/X VGND VGND VPWR VPWR _24032_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19392__A _19377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21559__B1 _23783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22097_ _20336_/A VGND VGND VPWR VPWR _22097_/X sky130_fd_sc_hd__buf_2
X_21048_ _20486_/X _21045_/X _24076_/Q _21042_/X VGND VGND VPWR VPWR _21048_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21427__A _21441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22220__B2 _22184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15425__A _15406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13870_ _13885_/A _13800_/B VGND VGND VPWR VPWR _13870_/X sky130_fd_sc_hd__or2_4
XFILLER_41_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12821_ _13349_/A _12821_/B _12820_/X VGND VGND VPWR VPWR _12821_/X sky130_fd_sc_hd__and3_4
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18727__A1 _18022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22999_ _22998_/X VGND VGND VPWR VPWR HADDR[16] sky130_fd_sc_hd__inv_2
XFILLER_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12752_ _11856_/A _11630_/A _12717_/X _12264_/X _12751_/X VGND VGND VPWR VPWR _12752_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_131_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15540_ _11900_/A _15540_/B VGND VGND VPWR VPWR _15541_/C sky130_fd_sc_hd__or2_4
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22258__A _22258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11703_ _11702_/X VGND VGND VPWR VPWR _16047_/A sky130_fd_sc_hd__buf_2
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21162__A _21155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15471_ _12592_/A _15471_/B VGND VGND VPWR VPWR _15471_/X sky130_fd_sc_hd__or2_4
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12574_/X _12680_/X _12682_/Y VGND VGND VPWR VPWR _12683_/X sky130_fd_sc_hd__a21o_4
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12784__A _12783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14430_/A _14485_/B VGND VGND VPWR VPWR _14423_/C sky130_fd_sc_hd__or2_4
XANTENNA__15160__A _13791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17210_ _17128_/A _17206_/X _12093_/X _17209_/X VGND VGND VPWR VPWR _17210_/X sky130_fd_sc_hd__o22a_4
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _20095_/D _11633_/X VGND VGND VPWR VPWR _11634_/X sky130_fd_sc_hd__or2_4
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18190_ _18190_/A _18217_/C _18148_/A _18148_/B VGND VGND VPWR VPWR _18190_/X sky130_fd_sc_hd__and4_4
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11578__A2 IRQ[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17141_ _14549_/Y _17115_/X _17140_/Y _17116_/X VGND VGND VPWR VPWR _17141_/X sky130_fd_sc_hd__o22a_4
X_14353_ _14390_/A VGND VGND VPWR VPWR _14366_/A sky130_fd_sc_hd__buf_2
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _24445_/Q IRQ[8] VGND VGND VPWR VPWR _11565_/X sky130_fd_sc_hd__and2_4
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17163__B1 _12982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13304_ _13304_/A _23462_/Q VGND VGND VPWR VPWR _13305_/C sky130_fd_sc_hd__or2_4
XANTENNA__23543__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17072_ _17197_/A VGND VGND VPWR VPWR _17198_/A sky130_fd_sc_hd__inv_2
XFILLER_171_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14284_ _14310_/A _14284_/B _14284_/C VGND VGND VPWR VPWR _14284_/X sky130_fd_sc_hd__or3_4
XFILLER_109_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20506__A _20334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16023_ _16033_/A VGND VGND VPWR VPWR _16062_/A sky130_fd_sc_hd__buf_2
X_13235_ _13235_/A _13233_/X _13234_/X VGND VGND VPWR VPWR _13236_/C sky130_fd_sc_hd__and3_4
XFILLER_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17087__A _17087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13166_ _13290_/A _13166_/B _13166_/C VGND VGND VPWR VPWR _13167_/C sky130_fd_sc_hd__and3_4
XANTENNA__21262__A2 _21257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12117_ _11705_/X _12114_/X _12116_/X VGND VGND VPWR VPWR _12123_/B sky130_fd_sc_hd__and3_4
X_13097_ _13097_/A _23624_/Q VGND VGND VPWR VPWR _13099_/B sky130_fd_sc_hd__or2_4
X_17974_ _18413_/A VGND VGND VPWR VPWR _17974_/X sky130_fd_sc_hd__buf_2
XANTENNA__12024__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19713_ _19508_/A VGND VGND VPWR VPWR _19899_/A sky130_fd_sc_hd__buf_2
X_16925_ _16899_/Y _16925_/B _16924_/X VGND VGND VPWR VPWR _16926_/C sky130_fd_sc_hd__and3_4
X_12048_ _16695_/A _12045_/X _12048_/C VGND VGND VPWR VPWR _12054_/B sky130_fd_sc_hd__and3_4
XANTENNA__22211__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12959__A _12971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11863__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24049__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19644_ _19811_/A VGND VGND VPWR VPWR _19644_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15335__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16856_ _15919_/D _16845_/X _15914_/X VGND VGND VPWR VPWR _16857_/B sky130_fd_sc_hd__o21a_4
XFILLER_168_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15807_ _12868_/A _15807_/B VGND VGND VPWR VPWR _15808_/C sky130_fd_sc_hd__or2_4
XANTENNA__11582__B IRQ[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19575_ _19703_/A HRDATA[12] VGND VGND VPWR VPWR _19575_/X sky130_fd_sc_hd__and2_4
XANTENNA__15054__B _23349_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16787_ _16053_/A _16787_/B _16787_/C VGND VGND VPWR VPWR _16819_/B sky130_fd_sc_hd__or3_4
XFILLER_81_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13999_ _12250_/A _13999_/B _13998_/X VGND VGND VPWR VPWR _13999_/X sky130_fd_sc_hd__and3_4
XANTENNA__22514__A2 _22508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18526_ _18477_/X _18503_/Y _18504_/X _18525_/X VGND VGND VPWR VPWR _18526_/X sky130_fd_sc_hd__o22a_4
X_15738_ _15778_/A _15682_/B VGND VGND VPWR VPWR _15738_/X sky130_fd_sc_hd__or2_4
XANTENNA__20525__A1 _18238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18457_ _18456_/X VGND VGND VPWR VPWR _18457_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12694__A _12687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15669_ _12704_/A _15667_/X _15669_/C VGND VGND VPWR VPWR _15669_/X sky130_fd_sc_hd__and3_4
XANTENNA__16166__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15070__A _14773_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17408_ _13692_/Y _17354_/X _17027_/X _17407_/X VGND VGND VPWR VPWR _17410_/A sky130_fd_sc_hd__o22a_4
XFILLER_21_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18388_ _18131_/X _18387_/X _18053_/X VGND VGND VPWR VPWR _18388_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__22278__B2 _22277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17339_ _17339_/A _17339_/B VGND VGND VPWR VPWR _17341_/A sky130_fd_sc_hd__or2_4
XFILLER_146_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17154__B1 _12680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20350_ _20273_/X _20346_/X _24306_/Q _20349_/X VGND VGND VPWR VPWR _20350_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17709__B _17389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19009_ _19009_/A VGND VGND VPWR VPWR _19024_/A sky130_fd_sc_hd__buf_2
X_20281_ _20450_/B VGND VGND VPWR VPWR _20282_/A sky130_fd_sc_hd__buf_2
XFILLER_143_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14414__A _14334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13191__A1 _13307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22020_ _21855_/X _22017_/X _15455_/B _22014_/X VGND VGND VPWR VPWR _22020_/X sky130_fd_sc_hd__o22a_4
XFILLER_115_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17457__A1 _17453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21253__A2 _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24141__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17457__B2 _17456_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23971_ _23939_/CLK _21214_/X VGND VGND VPWR VPWR _15820_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22202__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12869__A _12869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11773__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22922_ _22922_/A VGND VGND VPWR VPWR _23078_/A sky130_fd_sc_hd__buf_2
XFILLER_151_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20764__A1 _18525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23416__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22853_ _22799_/X VGND VGND VPWR VPWR _22853_/X sky130_fd_sc_hd__buf_2
XFILLER_72_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17460__A _12982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21804_ _21600_/X _21770_/A _23637_/Q _21767_/A VGND VGND VPWR VPWR _21804_/X sky130_fd_sc_hd__o22a_4
X_22784_ _22784_/A VGND VGND VPWR VPWR _22784_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22078__A _22057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21735_ _21565_/X _21734_/X _23684_/Q _21731_/X VGND VGND VPWR VPWR _23684_/D sky130_fd_sc_hd__o22a_4
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16076__A _16048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22269__A1 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24454_ _23347_/CLK _24454_/D HRESETn VGND VGND VPWR VPWR _20157_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_101_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21666_ _21534_/X _21663_/X _23729_/Q _21660_/X VGND VGND VPWR VPWR _21666_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22269__B2 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22806__A _15117_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23405_ _23501_/CLK _22239_/X VGND VGND VPWR VPWR _16142_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21710__A _21717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20617_ _24421_/Q _20617_/B VGND VGND VPWR VPWR _20617_/Y sky130_fd_sc_hd__nand2_4
X_24385_ _24419_/CLK _24385_/D HRESETn VGND VGND VPWR VPWR _19066_/A sky130_fd_sc_hd__dfstp_4
X_21597_ _21596_/X _21590_/X _15130_/B _21524_/X VGND VGND VPWR VPWR _21597_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12109__A _11868_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23336_ _23592_/CLK _22334_/X VGND VGND VPWR VPWR _23336_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20548_ _20540_/X _20546_/X _11535_/A _20547_/X VGND VGND VPWR VPWR _20548_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16523__B _16523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11948__A _11939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23267_ _23203_/CLK _23267_/D VGND VGND VPWR VPWR _15789_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14324__A _11933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20479_ _18178_/X _20469_/X _20341_/X _20478_/Y VGND VGND VPWR VPWR _20479_/X sky130_fd_sc_hd__a211o_4
X_13020_ _12877_/A _13018_/X _13019_/X VGND VGND VPWR VPWR _13024_/B sky130_fd_sc_hd__and3_4
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22218_ _22163_/X _22215_/X _23416_/Q _22212_/X VGND VGND VPWR VPWR _23416_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15139__B _15139_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22441__B2 _22433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23198_ _23679_/CLK _22574_/X VGND VGND VPWR VPWR _13721_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14043__B _24000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22541__A _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22149_ _20818_/A VGND VGND VPWR VPWR _22149_/X sky130_fd_sc_hd__buf_2
XFILLER_160_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14971_ _14786_/A _14971_/B _14970_/X VGND VGND VPWR VPWR _14971_/X sky130_fd_sc_hd__and3_4
XFILLER_94_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13485__A2 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12779__A _12778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20204__B1 _20200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11683__A _13123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16710_ _16710_/A _16710_/B _16710_/C VGND VGND VPWR VPWR _16710_/X sky130_fd_sc_hd__or3_4
X_13922_ _14377_/A _13839_/B VGND VGND VPWR VPWR _13923_/C sky130_fd_sc_hd__or2_4
X_17690_ _17698_/A VGND VGND VPWR VPWR _17690_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16641_ _16659_/A _16638_/X _16641_/C VGND VGND VPWR VPWR _16641_/X sky130_fd_sc_hd__and3_4
XANTENNA__24341__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13853_ _13853_/A VGND VGND VPWR VPWR _15450_/A sky130_fd_sc_hd__buf_2
XANTENNA__14994__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17370__A _17170_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12804_ _12834_/A _12804_/B VGND VGND VPWR VPWR _12804_/X sky130_fd_sc_hd__or2_4
X_19360_ _19358_/X _18450_/X _19358_/X _24259_/Q VGND VGND VPWR VPWR _24259_/D sky130_fd_sc_hd__a2bb2o_4
X_16572_ _16539_/X _23986_/Q VGND VGND VPWR VPWR _16572_/X sky130_fd_sc_hd__or2_4
X_13784_ _13784_/A VGND VGND VPWR VPWR _13785_/B sky130_fd_sc_hd__inv_2
X_18311_ _18376_/A _17522_/B VGND VGND VPWR VPWR _18311_/Y sky130_fd_sc_hd__nor2_4
X_15523_ _12258_/A _15523_/B VGND VGND VPWR VPWR _15524_/C sky130_fd_sc_hd__or2_4
X_12735_ _12735_/A _12833_/B VGND VGND VPWR VPWR _12735_/X sky130_fd_sc_hd__or2_4
X_19291_ _19240_/X VGND VGND VPWR VPWR _19291_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21180__B2 _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18242_ _17683_/A _18241_/X _17683_/A _18241_/X VGND VGND VPWR VPWR _18242_/X sky130_fd_sc_hd__a2bb2o_4
X_12666_ _12944_/A _12664_/X _12665_/X VGND VGND VPWR VPWR _12666_/X sky130_fd_sc_hd__and3_4
X_15454_ _14369_/A _15454_/B VGND VGND VPWR VPWR _15454_/X sky130_fd_sc_hd__or2_4
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21620__A _21620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14405_ _14512_/A _14405_/B _14404_/X VGND VGND VPWR VPWR _14409_/B sky130_fd_sc_hd__and3_4
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _12466_/A VGND VGND VPWR VPWR _11618_/A sky130_fd_sc_hd__buf_2
X_18173_ _17490_/D _18172_/X _17541_/Y VGND VGND VPWR VPWR _18173_/Y sky130_fd_sc_hd__o21ai_4
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12597_/A VGND VGND VPWR VPWR _12954_/A sky130_fd_sc_hd__buf_2
X_15385_ _15185_/X _15252_/X _15382_/X _15384_/Y VGND VGND VPWR VPWR _15385_/X sky130_fd_sc_hd__a211o_4
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ _17164_/A VGND VGND VPWR VPWR _17124_/X sky130_fd_sc_hd__buf_2
XANTENNA__21483__A2 _21478_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11548_ _24444_/Q IRQ[7] _11547_/X VGND VGND VPWR VPWR _11549_/B sky130_fd_sc_hd__a21o_4
X_14336_ _13884_/A VGND VGND VPWR VPWR _14516_/A sky130_fd_sc_hd__buf_2
XFILLER_156_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22680__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20236__A _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11858__A _11858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17055_ _17055_/A VGND VGND VPWR VPWR _17103_/A sky130_fd_sc_hd__inv_2
X_14267_ _14267_/A VGND VGND VPWR VPWR _14278_/A sky130_fd_sc_hd__buf_2
XFILLER_109_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16006_ _16006_/A _16006_/B _16006_/C VGND VGND VPWR VPWR _16012_/B sky130_fd_sc_hd__and3_4
X_13218_ _13235_/A _13216_/X _13217_/X VGND VGND VPWR VPWR _13218_/X sky130_fd_sc_hd__and3_4
XANTENNA__11577__B IRQ[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14198_ _11654_/A VGND VGND VPWR VPWR _14201_/A sky130_fd_sc_hd__buf_2
XFILLER_124_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13149_ _13333_/A _23559_/Q VGND VGND VPWR VPWR _13150_/C sky130_fd_sc_hd__or2_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17957_ _17911_/X _17917_/Y _17952_/X _17955_/Y _17956_/X VGND VGND VPWR VPWR _17957_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_111_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18939__A1 _15380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22735__A2 _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15065__A _15091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16908_ _13580_/Y _16907_/X _16528_/X VGND VGND VPWR VPWR _16908_/X sky130_fd_sc_hd__a21o_4
X_17888_ _17260_/A _17887_/X VGND VGND VPWR VPWR _17888_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24368__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19627_ _19898_/B _19622_/X _19533_/B _19890_/B VGND VGND VPWR VPWR _19628_/B sky130_fd_sc_hd__o22a_4
XFILLER_38_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16839_ _16830_/X _13585_/X _13573_/B VGND VGND VPWR VPWR _16839_/X sky130_fd_sc_hd__o21a_4
XFILLER_26_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23589__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19558_ _19558_/A _19557_/Y VGND VGND VPWR VPWR _19558_/X sky130_fd_sc_hd__or2_4
XFILLER_59_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22499__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_24_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18509_ _18418_/Y _17436_/A _17438_/X VGND VGND VPWR VPWR _18509_/X sky130_fd_sc_hd__o21a_4
XFILLER_90_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19489_ _19539_/A VGND VGND VPWR VPWR _19545_/A sky130_fd_sc_hd__inv_2
XANTENNA__21171__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21520_ _23796_/Q VGND VGND VPWR VPWR _21520_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14128__B _23583_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21530__A _21542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21451_ _21285_/X _21448_/X _15494_/B _21445_/X VGND VGND VPWR VPWR _23842_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20402_ _20402_/A _20450_/B VGND VGND VPWR VPWR _20402_/X sky130_fd_sc_hd__or2_4
XANTENNA__24322__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24170_ _24184_/CLK _24170_/D HRESETn VGND VGND VPWR VPWR _24170_/Q sky130_fd_sc_hd__dfrtp_4
X_21382_ _21251_/X _21377_/X _16446_/B _21381_/X VGND VGND VPWR VPWR _21382_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22671__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23121_ _23889_/CLK _22697_/X VGND VGND VPWR VPWR _23121_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11768__A _16048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20333_ _24275_/Q _20305_/X _20332_/X VGND VGND VPWR VPWR _20334_/B sky130_fd_sc_hd__o21a_4
XANTENNA__24214__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23052_ _23036_/X _18070_/A _23048_/X _23051_/X VGND VGND VPWR VPWR _23053_/A sky130_fd_sc_hd__a211o_4
X_20264_ _11634_/X _18889_/B VGND VGND VPWR VPWR _20264_/X sky130_fd_sc_hd__or2_4
XANTENNA__22361__A _22357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22003_ _22010_/A VGND VGND VPWR VPWR _22003_/X sky130_fd_sc_hd__buf_2
XFILLER_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20195_ _11636_/A _20195_/B VGND VGND VPWR VPWR _20195_/X sky130_fd_sc_hd__and2_4
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_106_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR _24102_/CLK sky130_fd_sc_hd__clkbuf_1
X_23954_ _23728_/CLK _23954_/D VGND VGND VPWR VPWR _23954_/Q sky130_fd_sc_hd__dfxtp_4
X_22905_ _22904_/X VGND VGND VPWR VPWR HADDR[0] sky130_fd_sc_hd__inv_2
XFILLER_29_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23885_ _24077_/CLK _21386_/X VGND VGND VPWR VPWR _23885_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15703__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22836_ _22801_/X VGND VGND VPWR VPWR _22836_/X sky130_fd_sc_hd__buf_2
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15422__B _23906_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22767_ SYSTICKCLKDIV[5] _22766_/A _22765_/Y _22766_/Y VGND VGND VPWR VPWR _22768_/D
+ sky130_fd_sc_hd__o22a_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14319__A _14319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _12499_/A _12520_/B VGND VGND VPWR VPWR _12522_/B sky130_fd_sc_hd__or2_4
X_21718_ _21536_/X _21713_/X _16403_/B _21717_/X VGND VGND VPWR VPWR _21718_/X sky130_fd_sc_hd__o22a_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22698_ _22698_/A VGND VGND VPWR VPWR _22698_/X sky130_fd_sc_hd__buf_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14038__B _23168_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12450_/X VGND VGND VPWR VPWR _15017_/A sky130_fd_sc_hd__buf_2
XFILLER_36_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24437_ _24422_/CLK _24437_/D HRESETn VGND VGND VPWR VPWR _24437_/Q sky130_fd_sc_hd__dfrtp_4
X_21649_ _21589_/X _21648_/X _14627_/B _21645_/X VGND VGND VPWR VPWR _23738_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16534__A _11960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15170_ _13799_/A _15170_/B VGND VGND VPWR VPWR _15170_/X sky130_fd_sc_hd__or2_4
X_12382_ _12827_/A _12268_/B VGND VGND VPWR VPWR _12384_/B sky130_fd_sc_hd__or2_4
X_24368_ _24368_/CLK _24368_/D HRESETn VGND VGND VPWR VPWR _24368_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21465__A2 _21462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14121_ _14148_/A _23551_/Q VGND VGND VPWR VPWR _14121_/X sky130_fd_sc_hd__or2_4
XANTENNA__11678__A _13383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23319_ _23416_/CLK _23319_/D VGND VGND VPWR VPWR _15213_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19845__A _17296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24299_ _24357_/CLK _19276_/X HRESETn VGND VGND VPWR VPWR _24299_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_67_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14054__A _13719_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21217__A2 _21212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14052_ _13700_/A _14052_/B VGND VGND VPWR VPWR _14052_/X sky130_fd_sc_hd__or2_4
XFILLER_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14989__A _15017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13003_ _12506_/A _24008_/Q VGND VGND VPWR VPWR _13004_/C sky130_fd_sc_hd__or2_4
XFILLER_106_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13893__A _14348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18860_ _13266_/X _18856_/X _24424_/Q _18857_/X VGND VGND VPWR VPWR _18860_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23086__B _23086_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20976__A1 _20305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20976__B2 _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17811_ _17810_/X VGND VGND VPWR VPWR _17811_/X sky130_fd_sc_hd__buf_2
X_18791_ _11851_/X _18787_/X _24468_/Q _18790_/X VGND VGND VPWR VPWR _24468_/D sky130_fd_sc_hd__o22a_4
XFILLER_130_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22717__A2 _22715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17742_ _17741_/A _17286_/X VGND VGND VPWR VPWR _17744_/A sky130_fd_sc_hd__and2_4
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14954_ _14973_/A _23606_/Q VGND VGND VPWR VPWR _14954_/X sky130_fd_sc_hd__or2_4
XANTENNA__12302__A _11887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13905_ _14507_/A _23997_/Q VGND VGND VPWR VPWR _13906_/C sky130_fd_sc_hd__or2_4
X_17673_ _17666_/X _17672_/Y VGND VGND VPWR VPWR _17673_/X sky130_fd_sc_hd__or2_4
X_14885_ _12425_/A _14883_/X _14884_/X VGND VGND VPWR VPWR _14885_/X sky130_fd_sc_hd__and3_4
XFILLER_78_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19412_ _19411_/X _18332_/X _19411_/X _24230_/Q VGND VGND VPWR VPWR _19412_/X sky130_fd_sc_hd__a2bb2o_4
X_16624_ _16654_/A _24050_/Q VGND VGND VPWR VPWR _16624_/X sky130_fd_sc_hd__or2_4
X_13836_ _15404_/A _13834_/X _13835_/X VGND VGND VPWR VPWR _13837_/C sky130_fd_sc_hd__and3_4
XFILLER_35_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19343_ _19340_/A VGND VGND VPWR VPWR _19343_/X sky130_fd_sc_hd__buf_2
XFILLER_62_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16555_ _16554_/X _24018_/Q VGND VGND VPWR VPWR _16556_/C sky130_fd_sc_hd__or2_4
X_13767_ _13743_/A _13767_/B _13766_/X VGND VGND VPWR VPWR _13767_/X sky130_fd_sc_hd__and3_4
XFILLER_16_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21153__B2 _21152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15506_ _13058_/A _15506_/B _15505_/X VGND VGND VPWR VPWR _15506_/X sky130_fd_sc_hd__and3_4
X_12718_ _13016_/A VGND VGND VPWR VPWR _13307_/A sky130_fd_sc_hd__buf_2
X_19274_ _24300_/Q _19248_/X _19273_/Y VGND VGND VPWR VPWR _24300_/D sky130_fd_sc_hd__o21a_4
X_16486_ _16210_/A _16486_/B _16485_/X VGND VGND VPWR VPWR _16487_/C sky130_fd_sc_hd__and3_4
X_13698_ _15325_/A VGND VGND VPWR VPWR _13699_/A sky130_fd_sc_hd__buf_2
X_18225_ _18283_/A _18225_/B _18225_/C _18224_/X VGND VGND VPWR VPWR _18225_/X sky130_fd_sc_hd__or4_4
X_15437_ _13639_/A _15509_/B VGND VGND VPWR VPWR _15438_/C sky130_fd_sc_hd__or2_4
XANTENNA__12972__A _12972_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12649_ _12954_/A _12645_/X _12649_/C VGND VGND VPWR VPWR _12649_/X sky130_fd_sc_hd__or3_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16444__A _11882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24237__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18156_ _18156_/A VGND VGND VPWR VPWR _18156_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21456__A2 _21455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22653__B2 _22648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15368_ _11735_/A _15368_/B _15367_/X VGND VGND VPWR VPWR _15369_/C sky130_fd_sc_hd__and3_4
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11588__A _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17107_ _17144_/A VGND VGND VPWR VPWR _17107_/X sky130_fd_sc_hd__buf_2
X_14319_ _14319_/A _24092_/Q VGND VGND VPWR VPWR _14320_/C sky130_fd_sc_hd__or2_4
XFILLER_116_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18087_ _17809_/A _18084_/X _17848_/A _18086_/X VGND VGND VPWR VPWR _18088_/A sky130_fd_sc_hd__o22a_4
X_15299_ _12444_/A _15299_/B _15299_/C VGND VGND VPWR VPWR _15303_/B sky130_fd_sc_hd__and3_4
XANTENNA__21208__A2 _21205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17038_ _17038_/A _17038_/B _17017_/A _16936_/A VGND VGND VPWR VPWR _17039_/A sky130_fd_sc_hd__or4_4
XANTENNA__14899__A _14170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18989_ _24398_/Q VGND VGND VPWR VPWR _18989_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12212__A _11880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21525__A _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20951_ _20754_/X _20950_/X _24312_/Q _20761_/X VGND VGND VPWR VPWR _20951_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17722__B _17427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21392__B2 _21388_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16619__A _16675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15523__A _12258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23670_ _23671_/CLK _23670_/D VGND VGND VPWR VPWR _14864_/B sky130_fd_sc_hd__dfxtp_4
X_20882_ _20782_/X _20881_/X _11521_/A _20789_/X VGND VGND VPWR VPWR _20882_/X sky130_fd_sc_hd__o22a_4
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22621_ _22459_/X _22615_/X _23168_/Q _22619_/X VGND VGND VPWR VPWR _23168_/D sky130_fd_sc_hd__o22a_4
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15242__B _15170_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21144__B2 _21138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18834__A _11609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13043__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22552_ _22425_/X _22551_/X _23214_/Q _22548_/X VGND VGND VPWR VPWR _23214_/D sky130_fd_sc_hd__o22a_4
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18553__B _18148_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21503_ _21489_/A VGND VGND VPWR VPWR _21503_/X sky130_fd_sc_hd__buf_2
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22483_ _22482_/X _22474_/X _14912_/B _22421_/A VGND VGND VPWR VPWR _23254_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12882__A _12882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24222_ _24248_/CLK _19423_/X HRESETn VGND VGND VPWR VPWR _24222_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21447__A2 _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21434_ _21441_/A VGND VGND VPWR VPWR _21434_/X sky130_fd_sc_hd__buf_2
XFILLER_148_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24153_ _24302_/CLK _20026_/Y HRESETn VGND VGND VPWR VPWR _17676_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_174_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21365_ _21309_/X _21362_/X _23896_/Q _21359_/X VGND VGND VPWR VPWR _21365_/X sky130_fd_sc_hd__o22a_4
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23104_ _23649_/CLK _23104_/D VGND VGND VPWR VPWR _23104_/Q sky130_fd_sc_hd__dfxtp_4
X_20316_ _20279_/B VGND VGND VPWR VPWR _20316_/X sky130_fd_sc_hd__buf_2
X_24084_ _23668_/CLK _24084_/D VGND VGND VPWR VPWR _24084_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_122_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21296_ _21295_/X _21293_/X _13732_/B _21288_/X VGND VGND VPWR VPWR _23934_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23035_ _23035_/A VGND VGND VPWR VPWR HADDR[22] sky130_fd_sc_hd__inv_2
X_20247_ _16918_/X _16922_/C _20247_/C _20247_/D VGND VGND VPWR VPWR _20248_/B sky130_fd_sc_hd__and4_4
XFILLER_66_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15417__B _15474_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20178_ _20178_/A _20177_/X VGND VGND VPWR VPWR _20178_/X sky130_fd_sc_hd__or2_4
XFILLER_103_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13218__A _13235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17913__A _18406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21907__B1 _12619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18728__B _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11951_ _11951_/A VGND VGND VPWR VPWR _11951_/X sky130_fd_sc_hd__buf_2
X_23937_ _23744_/CLK _23937_/D VGND VGND VPWR VPWR _15601_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21383__B2 _21381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22580__B1 _14560_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11961__A _12105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24351__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15433__A _12198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11882_ _13318_/A VGND VGND VPWR VPWR _11882_/X sky130_fd_sc_hd__buf_2
XFILLER_33_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14670_ _14679_/A _14587_/B VGND VGND VPWR VPWR _14671_/C sky130_fd_sc_hd__or2_4
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23868_ _23518_/CLK _21410_/X VGND VGND VPWR VPWR _14400_/B sky130_fd_sc_hd__dfxtp_4
X_13621_ _11877_/A VGND VGND VPWR VPWR _13622_/A sky130_fd_sc_hd__buf_2
X_22819_ _20700_/A VGND VGND VPWR VPWR _22819_/X sky130_fd_sc_hd__buf_2
XANTENNA__14049__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23799_ _23862_/CLK _23799_/D VGND VGND VPWR VPWR _15177_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18744__A _18744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16340_ _16313_/A _16338_/X _16339_/X VGND VGND VPWR VPWR _16340_/X sky130_fd_sc_hd__and3_4
XANTENNA__24244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13552_ _13503_/X _13552_/B _13552_/C VGND VGND VPWR VPWR _13556_/B sky130_fd_sc_hd__and3_4
XANTENNA__21686__A2 _21684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12503_ _12503_/A VGND VGND VPWR VPWR _12504_/A sky130_fd_sc_hd__buf_2
XANTENNA__13888__A _13888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13483_ _13483_/A _13483_/B VGND VGND VPWR VPWR _13483_/X sky130_fd_sc_hd__and2_4
X_16271_ _16099_/X _16271_/B VGND VGND VPWR VPWR _16272_/C sky130_fd_sc_hd__or2_4
XFILLER_41_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12792__A _13230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18010_ _17583_/A _18007_/B _18009_/X VGND VGND VPWR VPWR _18010_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15222_ _15196_/X _15222_/B VGND VGND VPWR VPWR _15222_/X sky130_fd_sc_hd__or2_4
X_12434_ _12434_/A VGND VGND VPWR VPWR _12435_/A sky130_fd_sc_hd__buf_2
XFILLER_139_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22635__B2 _22598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20217__C _17017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12365_ _12387_/A _12365_/B _12364_/X VGND VGND VPWR VPWR _12365_/X sky130_fd_sc_hd__and3_4
X_15153_ _15281_/A _15152_/X VGND VGND VPWR VPWR _15153_/X sky130_fd_sc_hd__and2_4
XFILLER_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14104_ _14137_/A _24031_/Q VGND VGND VPWR VPWR _14106_/B sky130_fd_sc_hd__or2_4
X_19961_ _19960_/X VGND VGND VPWR VPWR _19961_/X sky130_fd_sc_hd__buf_2
X_15084_ _11674_/A _15066_/X _15084_/C VGND VGND VPWR VPWR _15084_/X sky130_fd_sc_hd__or3_4
X_12296_ _13184_/A VGND VGND VPWR VPWR _13145_/A sky130_fd_sc_hd__buf_2
XANTENNA__22399__B1 _14717_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18912_ _12678_/X _18906_/X _19007_/A _18907_/X VGND VGND VPWR VPWR _24395_/D sky130_fd_sc_hd__o22a_4
X_14035_ _13700_/A _14035_/B VGND VGND VPWR VPWR _14035_/X sky130_fd_sc_hd__or2_4
XFILLER_136_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15608__A _13923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19892_ _19471_/X _19888_/X _19891_/Y _20216_/D _19512_/X VGND VGND VPWR VPWR _24185_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14512__A _14512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18843_ _18843_/A VGND VGND VPWR VPWR _18843_/X sky130_fd_sc_hd__buf_2
XFILLER_45_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14231__B _24063_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13128__A _12690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18774_ _18774_/A VGND VGND VPWR VPWR _18774_/X sky130_fd_sc_hd__buf_2
X_15986_ _15961_/A _15986_/B _15986_/C VGND VGND VPWR VPWR _15987_/C sky130_fd_sc_hd__and3_4
XFILLER_76_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21345__A _21338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17725_ _17726_/A _17407_/X VGND VGND VPWR VPWR _17729_/A sky130_fd_sc_hd__or2_4
X_14937_ _14976_/A _23158_/Q VGND VGND VPWR VPWR _14940_/B sky130_fd_sc_hd__or2_4
XFILLER_82_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12967__A _12943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22571__B1 _23200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11871__A _12186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15343__A _13704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17656_ _16997_/A VGND VGND VPWR VPWR _17780_/A sky130_fd_sc_hd__buf_2
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14868_ _14110_/A _14946_/B VGND VGND VPWR VPWR _14868_/X sky130_fd_sc_hd__or2_4
XFILLER_63_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16607_ _11705_/X VGND VGND VPWR VPWR _16646_/A sky130_fd_sc_hd__buf_2
X_13819_ _12198_/A _13819_/B VGND VGND VPWR VPWR _13819_/X sky130_fd_sc_hd__or2_4
XFILLER_50_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15062__B _24021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17587_ _18099_/A _17585_/Y _17586_/X VGND VGND VPWR VPWR _17587_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21126__B2 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14799_ _14679_/A _14731_/B VGND VGND VPWR VPWR _14800_/C sky130_fd_sc_hd__or2_4
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19326_ _16945_/X _17052_/Y _17654_/X _17784_/X VGND VGND VPWR VPWR _19327_/A sky130_fd_sc_hd__o22a_4
XFILLER_143_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16538_ _16534_/X _16615_/B VGND VGND VPWR VPWR _16541_/B sky130_fd_sc_hd__or2_4
XFILLER_50_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22176__A _22176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19257_ _24308_/Q VGND VGND VPWR VPWR _19257_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13798__A _13953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16469_ _16507_/A _16467_/X _16468_/X VGND VGND VPWR VPWR _16470_/C sky130_fd_sc_hd__and3_4
X_18208_ _17490_/D _18207_/X VGND VGND VPWR VPWR _18208_/X sky130_fd_sc_hd__or2_4
XFILLER_148_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21429__A2 _21427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19188_ _19148_/A _19148_/B _19187_/Y VGND VGND VPWR VPWR _24327_/D sky130_fd_sc_hd__o21a_4
XFILLER_157_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18139_ _18138_/A _18137_/X _17648_/X VGND VGND VPWR VPWR _18139_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17502__B1 _17028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21150_ _20464_/X _21148_/X _24013_/Q _21145_/X VGND VGND VPWR VPWR _21150_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20101_ _24476_/Q VGND VGND VPWR VPWR _20101_/Y sky130_fd_sc_hd__inv_2
X_21081_ _21081_/A _22039_/B _21234_/B VGND VGND VPWR VPWR _22637_/D sky130_fd_sc_hd__or3_4
XANTENNA__15518__A _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14422__A _14430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20032_ _24489_/Q VGND VGND VPWR VPWR _20032_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21601__A2 _21542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14141__B _24063_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13038__A _11935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21983_ _21877_/X _21981_/X _14724_/B _21978_/X VGND VGND VPWR VPWR _23545_/D sky130_fd_sc_hd__o22a_4
XFILLER_96_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12877__A _12877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21365__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23157__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11781__A _11781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23722_ _23723_/CLK _23722_/D VGND VGND VPWR VPWR _23722_/Q sky130_fd_sc_hd__dfxtp_4
X_20934_ _24249_/Q _20231_/A _20933_/X VGND VGND VPWR VPWR _20934_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24402__CLK _23281_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23653_ _23557_/CLK _21783_/X VGND VGND VPWR VPWR _23653_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _20865_/A VGND VGND VPWR VPWR _20940_/A sky130_fd_sc_hd__buf_2
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21117__B2 _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22604_ _22430_/X _22601_/X _12361_/B _22598_/X VGND VGND VPWR VPWR _23180_/D sky130_fd_sc_hd__o22a_4
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21668__A2 _21663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23584_ _23649_/CLK _23584_/D VGND VGND VPWR VPWR _23584_/Q sky130_fd_sc_hd__dfxtp_4
X_20796_ _20662_/X _20778_/X _20779_/X _20795_/Y VGND VGND VPWR VPWR _20796_/X sky130_fd_sc_hd__a211o_4
XFILLER_169_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22535_ _22484_/X _22508_/A _15033_/B _22498_/A VGND VGND VPWR VPWR _23221_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16084__A _11815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22466_ _20840_/A VGND VGND VPWR VPWR _22466_/X sky130_fd_sc_hd__buf_2
XFILLER_148_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22617__B2 _22612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22814__A _22884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20628__B1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24205_ _23126_/CLK _19674_/Y HRESETn VGND VGND VPWR VPWR _11611_/C sky130_fd_sc_hd__dfrtp_4
X_21417_ _21313_/X _21412_/X _23862_/Q _21381_/A VGND VGND VPWR VPWR _23862_/D sky130_fd_sc_hd__o22a_4
XFILLER_163_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12117__A _11705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22397_ _22357_/A VGND VGND VPWR VPWR _22397_/X sky130_fd_sc_hd__buf_2
X_12150_ _11762_/X _12148_/X _12150_/C VGND VGND VPWR VPWR _12150_/X sky130_fd_sc_hd__and3_4
X_24136_ _24137_/CLK _24136_/D HRESETn VGND VGND VPWR VPWR _24136_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21348_ _21341_/A VGND VGND VPWR VPWR _21348_/X sky130_fd_sc_hd__buf_2
XANTENNA__21840__A2 _21839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20334__A _20334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24067_ _23939_/CLK _21061_/X VGND VGND VPWR VPWR _15823_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15428__A _15405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12081_ _16695_/A _12081_/B _12081_/C VGND VGND VPWR VPWR _12085_/B sky130_fd_sc_hd__and3_4
X_21279_ _21278_/X _21269_/X _13512_/B _21276_/X VGND VGND VPWR VPWR _23941_/D sky130_fd_sc_hd__o22a_4
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14332__A _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23018_ _23018_/A VGND VGND VPWR VPWR HADDR[19] sky130_fd_sc_hd__inv_2
XFILLER_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18739__A _18738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15840_ _12878_/A _15840_/B VGND VGND VPWR VPWR _15842_/B sky130_fd_sc_hd__or2_4
XFILLER_77_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14986__B _23509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15771_ _15778_/A _15712_/B VGND VGND VPWR VPWR _15772_/C sky130_fd_sc_hd__or2_4
XANTENNA__24496__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17362__B _17445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12787__A _13563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23083__C _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12983_ _12914_/X _12983_/B VGND VGND VPWR VPWR _12983_/X sky130_fd_sc_hd__or2_4
XANTENNA__21356__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11691__A _13399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17510_ _11815_/X _17378_/X _17379_/X VGND VGND VPWR VPWR _17511_/B sky130_fd_sc_hd__o21a_4
X_14722_ _13622_/A _14722_/B _14722_/C VGND VGND VPWR VPWR _14722_/X sky130_fd_sc_hd__and3_4
X_11934_ _12266_/A VGND VGND VPWR VPWR _11935_/A sky130_fd_sc_hd__buf_2
X_18490_ _17805_/X _18285_/Y _18265_/X _18489_/Y VGND VGND VPWR VPWR _18490_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17441_ _14262_/X _17441_/B VGND VGND VPWR VPWR _17441_/X sky130_fd_sc_hd__or2_4
X_14653_ _14653_/A _14567_/B VGND VGND VPWR VPWR _14655_/B sky130_fd_sc_hd__or2_4
X_11865_ _13483_/A VGND VGND VPWR VPWR _11865_/X sky130_fd_sc_hd__buf_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13604_ _15415_/A VGND VGND VPWR VPWR _13657_/A sky130_fd_sc_hd__buf_2
XPHY_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17372_ _17372_/A VGND VGND VPWR VPWR _17446_/B sky130_fd_sc_hd__inv_2
X_11796_ _16635_/A _11793_/X _11796_/C VGND VGND VPWR VPWR _11796_/X sky130_fd_sc_hd__and3_4
X_14584_ _12454_/A _14584_/B VGND VGND VPWR VPWR _14584_/X sky130_fd_sc_hd__or2_4
XFILLER_159_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19111_ _24377_/Q VGND VGND VPWR VPWR _19111_/Y sky130_fd_sc_hd__inv_2
X_16323_ _16314_/X _16323_/B _16323_/C VGND VGND VPWR VPWR _16323_/X sky130_fd_sc_hd__and3_4
X_13535_ _13535_/A _24069_/Q VGND VGND VPWR VPWR _13536_/C sky130_fd_sc_hd__or2_4
XFILLER_159_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14507__A _14507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13411__A _13378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19042_ _19040_/Y _19041_/Y _11532_/B VGND VGND VPWR VPWR _19042_/X sky130_fd_sc_hd__o21a_4
XFILLER_51_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16254_ _16123_/A _16251_/X _16253_/X VGND VGND VPWR VPWR _16254_/X sky130_fd_sc_hd__and3_4
XFILLER_173_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13466_ _13443_/A _13546_/B VGND VGND VPWR VPWR _13467_/C sky130_fd_sc_hd__or2_4
XFILLER_158_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15205_ _14631_/A _15205_/B _15204_/X VGND VGND VPWR VPWR _15205_/X sky130_fd_sc_hd__and3_4
XANTENNA__13130__B _13199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12417_ _12676_/A _12396_/X _12417_/C VGND VGND VPWR VPWR _12417_/X sky130_fd_sc_hd__or3_4
X_16185_ _16185_/A _16185_/B _16184_/X VGND VGND VPWR VPWR _16186_/C sky130_fd_sc_hd__and3_4
XFILLER_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19485__B1 HRDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22084__A2 _22081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13397_ _13397_/A _23430_/Q VGND VGND VPWR VPWR _13398_/C sky130_fd_sc_hd__or2_4
XANTENNA__12027__A _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_14_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR _23347_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15136_ _15294_/A _15136_/B VGND VGND VPWR VPWR _15137_/C sky130_fd_sc_hd__or2_4
X_12348_ _13235_/A VGND VGND VPWR VPWR _12387_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_77_0_HCLK clkbuf_7_77_0_HCLK/A VGND VGND VPWR VPWR _23770_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_5_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11866__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15338__A _11752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12279_ _12279_/A VGND VGND VPWR VPWR _13276_/A sky130_fd_sc_hd__buf_2
X_19944_ _19938_/X _24165_/Q _19939_/X _20598_/B VGND VGND VPWR VPWR _24165_/D sky130_fd_sc_hd__o22a_4
X_15067_ _15075_/A _23925_/Q VGND VGND VPWR VPWR _15069_/B sky130_fd_sc_hd__or2_4
XANTENNA__14242__A _14615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14018_ _13888_/A _23264_/Q VGND VGND VPWR VPWR _14018_/X sky130_fd_sc_hd__or2_4
X_19875_ _19894_/C _19873_/X _19874_/X _19879_/D _19811_/A VGND VGND VPWR VPWR _19875_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21595__A1 _21594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21595__B2 _21585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22739__A2_N _22736_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17553__A _17120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18826_ _14548_/X _18824_/X _24443_/Q _18825_/X VGND VGND VPWR VPWR _24443_/D sky130_fd_sc_hd__o22a_4
X_18757_ _17980_/X _18753_/Y _17869_/A _18756_/Y VGND VGND VPWR VPWR _18757_/X sky130_fd_sc_hd__a211o_4
X_15969_ _15969_/A _23566_/Q VGND VGND VPWR VPWR _15970_/C sky130_fd_sc_hd__or2_4
XANTENNA__16169__A _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21347__B2 _21345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12697__A _12721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17708_ _17708_/A _17381_/X VGND VGND VPWR VPWR _17710_/A sky130_fd_sc_hd__and2_4
XANTENNA__15073__A _15112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21898__A2 _21895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18688_ _18689_/A _18687_/Y VGND VGND VPWR VPWR _18688_/X sky130_fd_sc_hd__or2_4
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17639_ _17639_/A _17605_/X _17638_/Y VGND VGND VPWR VPWR _17640_/D sky130_fd_sc_hd__or3_4
XFILLER_91_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20650_ _20516_/X _20649_/X _11530_/A _20475_/X VGND VGND VPWR VPWR _20650_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20419__A _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19309_ _19231_/X VGND VGND VPWR VPWR _19309_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20581_ _20581_/A _20494_/B VGND VGND VPWR VPWR _20581_/X sky130_fd_sc_hd__or2_4
XFILLER_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22320_ _22167_/X _22315_/X _14852_/B _22284_/A VGND VGND VPWR VPWR _22320_/X sky130_fd_sc_hd__o22a_4
XFILLER_149_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22251_ _22244_/A VGND VGND VPWR VPWR _22251_/X sky130_fd_sc_hd__buf_2
XANTENNA__22075__A2 _22074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21202_ _21202_/A VGND VGND VPWR VPWR _21202_/X sky130_fd_sc_hd__buf_2
XFILLER_105_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22182_ _22101_/X _22180_/X _16665_/B _22177_/X VGND VGND VPWR VPWR _22182_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21133_ _21133_/A VGND VGND VPWR VPWR _21134_/C sky130_fd_sc_hd__buf_2
XFILLER_160_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14152__A _13955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21064_ _20745_/X _21059_/X _24065_/Q _21063_/X VGND VGND VPWR VPWR _24065_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21586__A1 _21584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21586__B2 _21585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20015_ _20014_/X VGND VGND VPWR VPWR _24155_/D sky130_fd_sc_hd__inv_2
XFILLER_28_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13991__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17463__A _16702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18451__B2 _18450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20794__C1 _20793_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16079__A _16079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22535__B1 _15033_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21966_ _21848_/X _21960_/X _23557_/Q _21964_/X VGND VGND VPWR VPWR _21966_/X sky130_fd_sc_hd__o22a_4
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20010__A1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22809__A _14767_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21713__A _21727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23705_ _23101_/CLK _23705_/D VGND VGND VPWR VPWR _14760_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20917_ _20865_/A _20917_/B VGND VGND VPWR VPWR _20917_/X sky130_fd_sc_hd__or2_4
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _21817_/X _21895_/X _23602_/Q _21892_/X VGND VGND VPWR VPWR _23602_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16807__A _16611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15711__A _11887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11650_ _11750_/A VGND VGND VPWR VPWR _15321_/A sky130_fd_sc_hd__buf_2
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23636_ _23668_/CLK _23636_/D VGND VGND VPWR VPWR _21805_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22838__A1 _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20848_ _24412_/Q _20645_/X _24444_/Q _20704_/X VGND VGND VPWR VPWR _20848_/X sky130_fd_sc_hd__o22a_4
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20329__A _20313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _24467_/Q IRQ[30] VGND VGND VPWR VPWR _20125_/A sky130_fd_sc_hd__and2_4
XFILLER_156_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23567_ _23918_/CLK _23567_/D VGND VGND VPWR VPWR _16267_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ _20253_/Y VGND VGND VPWR VPWR _20779_/X sky130_fd_sc_hd__buf_2
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14327__A _12469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _13320_/A _23430_/Q VGND VGND VPWR VPWR _13320_/X sky130_fd_sc_hd__or2_4
XFILLER_35_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22518_ _22454_/X _22515_/X _15511_/B _22512_/X VGND VGND VPWR VPWR _22518_/X sky130_fd_sc_hd__o22a_4
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23498_ _23531_/CLK _22059_/X VGND VGND VPWR VPWR _12833_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_10_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22544__A _22558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22066__A2 _22060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13251_ _13251_/A _13247_/X _13251_/C VGND VGND VPWR VPWR _13259_/B sky130_fd_sc_hd__or3_4
XFILLER_129_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22449_ _20658_/A VGND VGND VPWR VPWR _22449_/X sky130_fd_sc_hd__buf_2
XANTENNA__16542__A _12108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12202_ _11915_/A VGND VGND VPWR VPWR _12691_/A sky130_fd_sc_hd__buf_2
X_13182_ _12866_/A _13182_/B _13181_/X VGND VGND VPWR VPWR _13182_/X sky130_fd_sc_hd__or3_4
XANTENNA__20064__A _18670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11686__A _16187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12133_ _12164_/A _23603_/Q VGND VGND VPWR VPWR _12134_/C sky130_fd_sc_hd__or2_4
X_24119_ _23991_/CLK _24119_/D HRESETn VGND VGND VPWR VPWR _22773_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17990_ _17986_/X _17987_/X _17988_/X _17989_/X VGND VGND VPWR VPWR _17991_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24448__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16941_ _16940_/Y VGND VGND VPWR VPWR _16941_/X sky130_fd_sc_hd__buf_2
X_12064_ _12103_/A VGND VGND VPWR VPWR _12064_/X sky130_fd_sc_hd__buf_2
XFILLER_123_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14997__A _13953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19660_ _19660_/A VGND VGND VPWR VPWR _19665_/B sky130_fd_sc_hd__inv_2
XANTENNA__17373__A _17169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16872_ _15388_/X _14552_/Y _16871_/Y _14552_/A VGND VGND VPWR VPWR _16873_/D sky130_fd_sc_hd__o22a_4
XFILLER_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18611_ _18610_/X VGND VGND VPWR VPWR _18611_/Y sky130_fd_sc_hd__inv_2
X_15823_ _12860_/A _15823_/B VGND VGND VPWR VPWR _15823_/X sky130_fd_sc_hd__or2_4
X_19591_ _19446_/A _19590_/X HRDATA[4] _19461_/X VGND VGND VPWR VPWR _19750_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21329__B2 _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13406__A _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18542_ _18095_/A _18229_/Y VGND VGND VPWR VPWR _18542_/X sky130_fd_sc_hd__and2_4
X_15754_ _13090_/A _15754_/B _15754_/C VGND VGND VPWR VPWR _15758_/B sky130_fd_sc_hd__and3_4
X_12966_ _12942_/A _23721_/Q VGND VGND VPWR VPWR _12966_/X sky130_fd_sc_hd__or2_4
XFILLER_161_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20001__A1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22719__A _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14705_ _14705_/A _14704_/X VGND VGND VPWR VPWR _14705_/X sky130_fd_sc_hd__or2_4
X_11917_ _12515_/A VGND VGND VPWR VPWR _11917_/X sky130_fd_sc_hd__buf_2
X_18473_ _18330_/X _18457_/Y _18373_/X _18472_/X VGND VGND VPWR VPWR _18473_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19942__B2 _20561_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15685_ _11970_/A _15684_/X VGND VGND VPWR VPWR _15685_/X sky130_fd_sc_hd__and2_4
X_12897_ _12874_/A _12893_/X _12897_/C VGND VGND VPWR VPWR _12897_/X sky130_fd_sc_hd__or3_4
XANTENNA__16717__A _16568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17424_ _17635_/A VGND VGND VPWR VPWR _17436_/C sky130_fd_sc_hd__inv_2
XFILLER_127_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14636_ _11708_/A VGND VGND VPWR VPWR _14677_/A sky130_fd_sc_hd__buf_2
X_11848_ _16768_/A _11848_/B _11847_/X VGND VGND VPWR VPWR _11848_/X sky130_fd_sc_hd__or3_4
XPHY_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17418_/A VGND VGND VPWR VPWR _17360_/A sky130_fd_sc_hd__inv_2
X_14567_ _12530_/A _14567_/B VGND VGND VPWR VPWR _14567_/X sky130_fd_sc_hd__or2_4
X_11779_ _15362_/A VGND VGND VPWR VPWR _11780_/A sky130_fd_sc_hd__buf_2
XANTENNA__14237__A _14616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21501__B2 _21496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16306_ _15934_/X _16302_/X _16305_/X VGND VGND VPWR VPWR _16306_/X sky130_fd_sc_hd__or3_4
XFILLER_147_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13141__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13518_ _13554_/A _13518_/B VGND VGND VPWR VPWR _13518_/X sky130_fd_sc_hd__or2_4
X_17286_ _17285_/Y _17280_/B VGND VGND VPWR VPWR _17286_/X sky130_fd_sc_hd__or2_4
X_14498_ _11681_/A _14490_/X _14497_/X VGND VGND VPWR VPWR _14498_/X sky130_fd_sc_hd__and3_4
XANTENNA__22454__A _20718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17181__A1 _12077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19025_ _24360_/Q _11533_/X _19018_/Y VGND VGND VPWR VPWR _19025_/Y sky130_fd_sc_hd__a21oi_4
X_16237_ _16187_/A _16237_/B _16237_/C VGND VGND VPWR VPWR _16238_/C sky130_fd_sc_hd__and3_4
XFILLER_173_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13449_ _12867_/A _13449_/B VGND VGND VPWR VPWR _13451_/B sky130_fd_sc_hd__or2_4
XANTENNA__19458__B1 HRDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12980__A _12979_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21265__B1 _12618_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16168_ _16163_/X _16165_/X _16168_/C VGND VGND VPWR VPWR _16168_/X sky130_fd_sc_hd__and3_4
XANTENNA__21804__A2 _21770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15119_ _14911_/X _14984_/A _15117_/Y _15118_/X VGND VGND VPWR VPWR _15119_/X sky130_fd_sc_hd__o22a_4
X_16099_ _12561_/A VGND VGND VPWR VPWR _16099_/X sky130_fd_sc_hd__buf_2
X_19927_ _19921_/X _24178_/Q _19925_/X _20672_/A VGND VGND VPWR VPWR _19927_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17283__A _14549_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_7_0_HCLK clkbuf_7_6_0_HCLK/A VGND VGND VPWR VPWR _24277_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_69_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19858_ _19649_/A _19856_/X _19725_/A _19857_/X VGND VGND VPWR VPWR _19859_/B sky130_fd_sc_hd__o22a_4
XANTENNA__14700__A _11668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18809_ _17172_/X _18803_/X _20157_/A _18804_/X VGND VGND VPWR VPWR _24454_/D sky130_fd_sc_hd__o22a_4
XFILLER_23_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22517__B1 _15836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19789_ _19767_/A _19786_/X _19781_/A _19788_/X VGND VGND VPWR VPWR _19789_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21236__C _21184_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21820_ _21819_/X _21815_/X _23633_/Q _21810_/X VGND VGND VPWR VPWR _23633_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12220__A _12294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22629__A _22622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19933__B2 _20776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21751_ _21594_/X _21748_/X _23672_/Q _21745_/X VGND VGND VPWR VPWR _23672_/D sky130_fd_sc_hd__o22a_4
XFILLER_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21740__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15531__A _12236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20702_ _20260_/A VGND VGND VPWR VPWR _20702_/X sky130_fd_sc_hd__buf_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21682_ _21560_/X _21677_/X _23718_/Q _21681_/X VGND VGND VPWR VPWR _21682_/X sky130_fd_sc_hd__o22a_4
XFILLER_145_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24470_ _24137_/CLK _18743_/X HRESETn VGND VGND VPWR VPWR _24470_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20633_ _21848_/A VGND VGND VPWR VPWR _20633_/X sky130_fd_sc_hd__buf_2
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23421_ _23582_/CLK _22211_/X VGND VGND VPWR VPWR _13842_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22296__A2 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21242__A2_N _21240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19938__A _19920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23352_ _23290_/CLK _23352_/D VGND VGND VPWR VPWR _23352_/Q sky130_fd_sc_hd__dfxtp_4
X_20564_ _20470_/X _20563_/X _24392_/Q _20429_/X VGND VGND VPWR VPWR _20564_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22303_ _22137_/X _22301_/X _15853_/B _22298_/X VGND VGND VPWR VPWR _23363_/D sky130_fd_sc_hd__o22a_4
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22048__A2 _22046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17458__A _12982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23283_ _23379_/CLK _22415_/X VGND VGND VPWR VPWR _12114_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12890__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16362__A _13399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20495_ _20495_/A VGND VGND VPWR VPWR _20495_/X sky130_fd_sc_hd__buf_2
XFILLER_121_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23345__CLK _23409_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22234_ _22226_/X VGND VGND VPWR VPWR _22234_/X sky130_fd_sc_hd__buf_2
XFILLER_30_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22165_ _22480_/A VGND VGND VPWR VPWR _22165_/X sky130_fd_sc_hd__buf_2
XFILLER_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_60_0_HCLK clkbuf_6_30_0_HCLK/X VGND VGND VPWR VPWR _23467_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21008__B1 HRDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21116_ _20745_/X _21111_/X _24033_/Q _21115_/X VGND VGND VPWR VPWR _24033_/D sky130_fd_sc_hd__o22a_4
XFILLER_59_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21708__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22096_ _22088_/Y _22094_/X _22095_/X _22094_/X VGND VGND VPWR VPWR _22096_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20612__A _20612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21559__B2 _21549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22756__B1 SYSTICKCLKDIV[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21047_ _20464_/X _21045_/X _24077_/Q _21042_/X VGND VGND VPWR VPWR _21047_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15706__A _12741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22220__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14610__A _13589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13226__A _12338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12820_ _12834_/A _12731_/B VGND VGND VPWR VPWR _12820_/X sky130_fd_sc_hd__or2_4
XFILLER_90_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22998_ _22977_/X _17906_/A _22989_/X _22997_/X VGND VGND VPWR VPWR _22998_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22539__A _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18727__A2 _17005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12751_ _13307_/A _12726_/X _12733_/X _12742_/X _12750_/X VGND VGND VPWR VPWR _12751_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ _21819_/X _21946_/X _23569_/Q _21943_/X VGND VGND VPWR VPWR _23569_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16537__A _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11702_ _13367_/A VGND VGND VPWR VPWR _11702_/X sky130_fd_sc_hd__buf_2
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15441__A _12300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15477_/A _15470_/B VGND VGND VPWR VPWR _15470_/X sky130_fd_sc_hd__or2_4
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/A VGND VGND VPWR VPWR _12682_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14421_/A VGND VGND VPWR VPWR _14430_/A sky130_fd_sc_hd__buf_2
XANTENNA__24120__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ _23587_/CLK _21854_/X VGND VGND VPWR VPWR _15822_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19848__A _19848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11633_ _11632_/X VGND VGND VPWR VPWR _11633_/X sky130_fd_sc_hd__buf_2
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14057__A _11698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17140_ _17139_/X VGND VGND VPWR VPWR _17140_/Y sky130_fd_sc_hd__inv_2
X_14352_ _13697_/A VGND VGND VPWR VPWR _14383_/A sky130_fd_sc_hd__buf_2
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ _11561_/X _11563_/X VGND VGND VPWR VPWR _11564_/X sky130_fd_sc_hd__or2_4
XANTENNA__17163__A1 _17162_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _13303_/A _23174_/Q VGND VGND VPWR VPWR _13305_/B sky130_fd_sc_hd__or2_4
XFILLER_7_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13896__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17368__A _17360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17071_ _17070_/X VGND VGND VPWR VPWR _17197_/A sky130_fd_sc_hd__buf_2
X_14283_ _14448_/A _14283_/B _14282_/X VGND VGND VPWR VPWR _14284_/C sky130_fd_sc_hd__and3_4
XANTENNA__16272__A _11917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24270__CLK _24271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16022_ _16061_/A _23374_/Q VGND VGND VPWR VPWR _16025_/B sky130_fd_sc_hd__or2_4
XFILLER_13_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18190__C _18148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13234_ _13253_/A _24071_/Q VGND VGND VPWR VPWR _13234_/X sky130_fd_sc_hd__or2_4
XANTENNA__17087__B _17188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22995__B1 _22949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13165_ _13301_/A _24071_/Q VGND VGND VPWR VPWR _13166_/C sky130_fd_sc_hd__or2_4
XFILLER_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12305__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12116_ _16775_/A _23539_/Q VGND VGND VPWR VPWR _12116_/X sky130_fd_sc_hd__or2_4
XFILLER_97_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13096_ _13096_/A _13096_/B _13096_/C VGND VGND VPWR VPWR _13100_/B sky130_fd_sc_hd__and3_4
X_17973_ _17973_/A VGND VGND VPWR VPWR _17973_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22747__B1 _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12024__B _12020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19712_ _19849_/B _19712_/B _19899_/B VGND VGND VPWR VPWR _19712_/X sky130_fd_sc_hd__and3_4
X_16924_ _16915_/A _17060_/B _17091_/A _16898_/X VGND VGND VPWR VPWR _16924_/X sky130_fd_sc_hd__or4_4
XANTENNA__15616__A _15616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12047_ _16724_/A _23795_/Q VGND VGND VPWR VPWR _12048_/C sky130_fd_sc_hd__or2_4
XANTENNA__24440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22211__A2 _22208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19643_ _19643_/A VGND VGND VPWR VPWR _19811_/A sky130_fd_sc_hd__buf_2
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15335__B _23160_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16855_ _16855_/A VGND VGND VPWR VPWR _16855_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15806_ _12867_/A _23331_/Q VGND VGND VPWR VPWR _15808_/B sky130_fd_sc_hd__or2_4
XANTENNA__13136__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21970__B2 _21964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19574_ _19438_/B VGND VGND VPWR VPWR _19703_/A sky130_fd_sc_hd__buf_2
XANTENNA__17831__A _12077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16786_ _16786_/A _16778_/X _16785_/X VGND VGND VPWR VPWR _16787_/C sky130_fd_sc_hd__and3_4
XANTENNA__12040__A _11941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13998_ _13637_/A _24096_/Q VGND VGND VPWR VPWR _13998_/X sky130_fd_sc_hd__or2_4
XANTENNA__22449__A _20658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23218__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18525_ _18506_/X _18513_/Y _18514_/X _18516_/X _18524_/Y VGND VGND VPWR VPWR _18525_/X
+ sky130_fd_sc_hd__a32o_4
X_15737_ _15770_/A _15737_/B VGND VGND VPWR VPWR _15737_/X sky130_fd_sc_hd__or2_4
XFILLER_74_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12949_ _12949_/A _23977_/Q VGND VGND VPWR VPWR _12950_/C sky130_fd_sc_hd__or2_4
XFILLER_45_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12975__A _12975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16447__A _11917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21722__B2 _21717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18456_ _18022_/X _18368_/B _18454_/Y _18027_/X _22979_/B VGND VGND VPWR VPWR _18456_/X
+ sky130_fd_sc_hd__a32o_4
X_15668_ _12273_/A _15668_/B VGND VGND VPWR VPWR _15669_/C sky130_fd_sc_hd__or2_4
X_17407_ _17406_/Y _17280_/B VGND VGND VPWR VPWR _17407_/X sky130_fd_sc_hd__or2_4
X_14619_ _14665_/A VGND VGND VPWR VPWR _14820_/A sky130_fd_sc_hd__buf_2
X_18387_ _17977_/X _18159_/X _17856_/X _18132_/X VGND VGND VPWR VPWR _18387_/X sky130_fd_sc_hd__a2bb2o_4
X_15599_ _15625_/A _15599_/B _15599_/C VGND VGND VPWR VPWR _15600_/C sky130_fd_sc_hd__or3_4
XFILLER_159_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17338_ _17339_/B VGND VGND VPWR VPWR _17340_/B sky130_fd_sc_hd__inv_2
XFILLER_159_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17154__A1 _17153_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22184__A _22184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17278__A _11611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17269_ _17914_/B VGND VGND VPWR VPWR _17269_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19008_ _18987_/X _19006_/X _19007_/Y _18990_/X VGND VGND VPWR VPWR _19008_/X sky130_fd_sc_hd__o22a_4
XFILLER_161_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20280_ _20493_/A VGND VGND VPWR VPWR _20450_/B sky130_fd_sc_hd__buf_2
XANTENNA__22912__A _20218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21789__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18654__A1 _17805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_47_0_HCLK clkbuf_6_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21528__A _21528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17725__B _17407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22202__A2 _22201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15526__A _12258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23970_ _23587_/CLK _21215_/X VGND VGND VPWR VPWR _15487_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14430__A _14430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22921_ _22912_/X VGND VGND VPWR VPWR _22929_/A sky130_fd_sc_hd__buf_2
XFILLER_57_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21961__A1 _21838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18837__A _18837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21961__B2 _21957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13046__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22852_ _22851_/X VGND VGND VPWR VPWR HWDATA[16] sky130_fd_sc_hd__inv_2
XFILLER_25_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22359__A _22366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24143__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21803_ _21598_/X _21798_/X _23638_/Q _21767_/A VGND VGND VPWR VPWR _23638_/D sky130_fd_sc_hd__o22a_4
X_22783_ _22781_/Y _22786_/B _22793_/A VGND VGND VPWR VPWR _22783_/X sky130_fd_sc_hd__and3_4
XFILLER_25_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15261__A _15257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21734_ _21727_/A VGND VGND VPWR VPWR _21734_/X sky130_fd_sc_hd__buf_2
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18590__B1 _18585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22269__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24453_ _23475_/CLK _18812_/X HRESETn VGND VGND VPWR VPWR _24453_/Q sky130_fd_sc_hd__dfrtp_4
X_21665_ _21532_/X _21663_/X _23730_/Q _21660_/X VGND VGND VPWR VPWR _23730_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24293__CLK _24294_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23404_ _23404_/CLK _23404_/D VGND VGND VPWR VPWR _12392_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_71_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20616_ _20444_/X _22737_/A _20308_/A VGND VGND VPWR VPWR _20616_/X sky130_fd_sc_hd__a21o_4
XFILLER_32_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21596_ _21311_/A VGND VGND VPWR VPWR _21596_/X sky130_fd_sc_hd__buf_2
X_24384_ _24445_/CLK _18929_/X HRESETn VGND VGND VPWR VPWR _24384_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22094__A _22106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23335_ _23204_/CLK _22335_/X VGND VGND VPWR VPWR _13148_/B sky130_fd_sc_hd__dfxtp_4
X_20547_ _20267_/X VGND VGND VPWR VPWR _20547_/X sky130_fd_sc_hd__buf_2
XANTENNA__17188__A _17188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16092__A _16110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14605__A _12484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23266_ _23203_/CLK _23266_/D VGND VGND VPWR VPWR _15454_/B sky130_fd_sc_hd__dfxtp_4
X_20478_ _20388_/A _20478_/B VGND VGND VPWR VPWR _20478_/Y sky130_fd_sc_hd__nor2_4
X_22217_ _22161_/X _22215_/X _23417_/Q _22212_/X VGND VGND VPWR VPWR _23417_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22441__A2 _22438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23197_ _23229_/CLK _23197_/D VGND VGND VPWR VPWR _13807_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16820__A _16819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21438__A _21438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22148_ _22146_/X _22147_/X _23455_/Q _22142_/X VGND VGND VPWR VPWR _23455_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11964__A _12108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22079_ _21869_/X _22074_/X _23484_/Q _22078_/X VGND VGND VPWR VPWR _22079_/X sky130_fd_sc_hd__o22a_4
X_14970_ _14970_/A _23862_/Q VGND VGND VPWR VPWR _14970_/X sky130_fd_sc_hd__or2_4
XANTENNA__14340__A _12410_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20204__A1 _19402_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13485__A3 _13454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13921_ _14386_/A _13838_/B VGND VGND VPWR VPWR _13923_/B sky130_fd_sc_hd__or2_4
XFILLER_47_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15155__B _15155_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21952__B2 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20996__B _20996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16640_ _16677_/A _16640_/B VGND VGND VPWR VPWR _16641_/C sky130_fd_sc_hd__or2_4
X_13852_ _11625_/A VGND VGND VPWR VPWR _13853_/A sky130_fd_sc_hd__buf_2
XFILLER_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14994__B _23765_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12803_ _12833_/A _12803_/B VGND VGND VPWR VPWR _12803_/X sky130_fd_sc_hd__or2_4
XANTENNA__21173__A _21152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16571_ _16534_/X _23922_/Q VGND VGND VPWR VPWR _16573_/B sky130_fd_sc_hd__or2_4
XANTENNA__12795__A _13205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13783_ _13692_/Y _13781_/X VGND VGND VPWR VPWR _13784_/A sky130_fd_sc_hd__or2_4
XFILLER_167_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22901__B1 _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18310_ _18310_/A _17605_/D VGND VGND VPWR VPWR _18310_/X sky130_fd_sc_hd__or2_4
XANTENNA__21704__B2 _21667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15522_ _15439_/A _15522_/B VGND VGND VPWR VPWR _15522_/X sky130_fd_sc_hd__or2_4
XFILLER_37_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15171__A _14297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12734_ _12748_/A VGND VGND VPWR VPWR _12738_/A sky130_fd_sc_hd__buf_2
X_19290_ _24292_/Q _19240_/X _19289_/Y VGND VGND VPWR VPWR _24292_/D sky130_fd_sc_hd__o21a_4
XFILLER_37_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21180__A2 _21176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18241_ _17683_/B _18181_/X _17681_/X VGND VGND VPWR VPWR _18241_/X sky130_fd_sc_hd__o21a_4
XFILLER_30_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15453_ _15453_/A VGND VGND VPWR VPWR _15453_/Y sky130_fd_sc_hd__inv_2
X_12665_ _12974_/A _12665_/B VGND VGND VPWR VPWR _12665_/X sky130_fd_sc_hd__or2_4
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14511_/A _24092_/Q VGND VGND VPWR VPWR _14404_/X sky130_fd_sc_hd__or2_4
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _13662_/A VGND VGND VPWR VPWR _11869_/A sky130_fd_sc_hd__buf_2
X_18172_ _17490_/B _18234_/A _17539_/X VGND VGND VPWR VPWR _18172_/X sky130_fd_sc_hd__o21a_4
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15384_ _15384_/A VGND VGND VPWR VPWR _15384_/Y sky130_fd_sc_hd__inv_2
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _12596_/A VGND VGND VPWR VPWR _12597_/A sky130_fd_sc_hd__buf_2
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17123_ _17113_/X _17123_/B VGND VGND VPWR VPWR _17123_/X sky130_fd_sc_hd__or2_4
XANTENNA__17098__A _18485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14335_ _14335_/A VGND VGND VPWR VPWR _14513_/A sky130_fd_sc_hd__buf_2
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18884__A1 _15118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11547_ _24443_/Q IRQ[6] VGND VGND VPWR VPWR _11547_/X sky130_fd_sc_hd__and2_4
XFILLER_144_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14515__A _13229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22680__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20691__A1 _24227_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17054_ _17015_/X _17054_/B VGND VGND VPWR VPWR _17055_/A sky130_fd_sc_hd__or2_4
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14266_ _14266_/A _14266_/B VGND VGND VPWR VPWR _15391_/C sky130_fd_sc_hd__or2_4
XFILLER_171_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16005_ _15959_/A _23822_/Q VGND VGND VPWR VPWR _16006_/C sky130_fd_sc_hd__or2_4
XFILLER_100_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13217_ _13256_/A _13217_/B VGND VGND VPWR VPWR _13217_/X sky130_fd_sc_hd__or2_4
XFILLER_152_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14197_ _14631_/A _14195_/X _14196_/X VGND VGND VPWR VPWR _14202_/B sky130_fd_sc_hd__and3_4
XFILLER_152_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13148_ _13303_/A _13148_/B VGND VGND VPWR VPWR _13148_/X sky130_fd_sc_hd__or2_4
XANTENNA__21348__A _21341_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11874__A _13468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15346__A _15362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13079_ _13088_/A _13012_/B VGND VGND VPWR VPWR _13079_/X sky130_fd_sc_hd__or2_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17956_ _17911_/B _17955_/B _17890_/X VGND VGND VPWR VPWR _17956_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14250__A _13865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22196__B2 _22191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24166__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16907_ _12987_/X _16832_/X VGND VGND VPWR VPWR _16907_/X sky130_fd_sc_hd__or2_4
X_17887_ _17807_/A _17644_/X _18562_/A _17592_/X VGND VGND VPWR VPWR _17887_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17561__A _16383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19626_ _19848_/B VGND VGND VPWR VPWR _19890_/B sky130_fd_sc_hd__buf_2
X_16838_ _16527_/B _16837_/X _16527_/B _16837_/X VGND VGND VPWR VPWR _16838_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22179__A _22208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21083__A _21134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22499__A2 _22494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16769_ _16683_/A _16760_/X _16768_/X VGND VGND VPWR VPWR _16787_/B sky130_fd_sc_hd__and3_4
X_19557_ _19550_/B VGND VGND VPWR VPWR _19557_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15081__A _15081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18508_ _17635_/B _18507_/X VGND VGND VPWR VPWR _18508_/X sky130_fd_sc_hd__or2_4
XFILLER_62_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19488_ _19480_/X _19487_/X HRDATA[11] _19484_/X VGND VGND VPWR VPWR _19539_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21171__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22907__A _22906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18439_ _18485_/A _17393_/X VGND VGND VPWR VPWR _18439_/Y sky130_fd_sc_hd__nor2_4
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16905__A _16905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21450_ _21283_/X _21448_/X _15827_/B _21445_/X VGND VGND VPWR VPWR _23843_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18324__B1 _18060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20401_ _24463_/Q VGND VGND VPWR VPWR _20402_/A sky130_fd_sc_hd__inv_2
Xclkbuf_4_10_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_10_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21381_ _21381_/A VGND VGND VPWR VPWR _21381_/X sky130_fd_sc_hd__buf_2
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20131__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18875__A1 _13945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14425__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20146__B _20145_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23120_ _23728_/CLK _23120_/D VGND VGND VPWR VPWR _16442_/B sky130_fd_sc_hd__dfxtp_4
X_20332_ _20306_/X _20309_/X _20714_/A _20331_/Y VGND VGND VPWR VPWR _20332_/X sky130_fd_sc_hd__a211o_4
XFILLER_31_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14144__B _23135_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23051_ _23051_/A _23051_/B _23050_/X VGND VGND VPWR VPWR _23051_/X sky130_fd_sc_hd__and3_4
X_20263_ _20260_/A VGND VGND VPWR VPWR _20292_/A sky130_fd_sc_hd__inv_2
XFILLER_162_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22002_ _21824_/X _21996_/X _16248_/B _22000_/X VGND VGND VPWR VPWR _22002_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20194_ _20194_/A _20193_/X VGND VGND VPWR VPWR _20195_/B sky130_fd_sc_hd__or2_4
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20162__A IRQ[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19951__A _19950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14160__A _14988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12599__B _12599_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23953_ _23761_/CLK _23953_/D VGND VGND VPWR VPWR _23953_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21934__B2 _21899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22904_ _22742_/A _19953_/A _22738_/A _22904_/D VGND VGND VPWR VPWR _22904_/X sky130_fd_sc_hd__or4_4
XANTENNA__17471__A _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23884_ _23500_/CLK _21387_/X VGND VGND VPWR VPWR _12314_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22835_ _22884_/A VGND VGND VPWR VPWR _22845_/A sky130_fd_sc_hd__buf_2
XANTENNA__16087__A _16016_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22766_ _22766_/A VGND VGND VPWR VPWR _22766_/Y sky130_fd_sc_hd__inv_2
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22817__A _18738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21717_ _21717_/A VGND VGND VPWR VPWR _21717_/X sky130_fd_sc_hd__buf_2
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22697_ _21534_/A _22694_/X _23121_/Q _22691_/X VGND VGND VPWR VPWR _22697_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16815__A _16646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _12194_/A VGND VGND VPWR VPWR _12450_/X sky130_fd_sc_hd__buf_2
X_24436_ _23379_/CLK _18844_/X HRESETn VGND VGND VPWR VPWR _24436_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21648_ _21608_/A VGND VGND VPWR VPWR _21648_/X sky130_fd_sc_hd__buf_2
XANTENNA__20337__A _21528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11959__A _11891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18866__A1 _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ _12978_/A VGND VGND VPWR VPWR _12676_/A sky130_fd_sc_hd__buf_2
X_24367_ _24368_/CLK _24367_/D HRESETn VGND VGND VPWR VPWR _24367_/Q sky130_fd_sc_hd__dfstp_4
X_21579_ _21577_/X _21578_/X _23775_/Q _21573_/X VGND VGND VPWR VPWR _23775_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14335__A _14335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14120_ _14131_/A VGND VGND VPWR VPWR _14148_/A sky130_fd_sc_hd__buf_2
X_23318_ _23671_/CLK _22352_/X VGND VGND VPWR VPWR _14867_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24298_ _24357_/CLK _24298_/D HRESETn VGND VGND VPWR VPWR _19247_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24374__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14051_ _11812_/A VGND VGND VPWR VPWR _15649_/A sky130_fd_sc_hd__buf_2
X_23249_ _23379_/CLK _22497_/X VGND VGND VPWR VPWR _16813_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16550__A _11939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13002_ _12499_/A _23688_/Q VGND VGND VPWR VPWR _13004_/B sky130_fd_sc_hd__or2_4
XFILLER_137_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14989__B _23733_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11587__A2_N _11544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23086__C _23086_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20976__A2 _20967_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_30_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_30_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15166__A _12453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17810_ _17151_/X VGND VGND VPWR VPWR _17810_/X sky130_fd_sc_hd__buf_2
X_18790_ _18790_/A VGND VGND VPWR VPWR _18790_/X sky130_fd_sc_hd__buf_2
XANTENNA__14070__A _11735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22178__B2 _22177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17741_ _17741_/A _17286_/X VGND VGND VPWR VPWR _17758_/A sky130_fd_sc_hd__or2_4
X_14953_ _14916_/X _14951_/X _14952_/X VGND VGND VPWR VPWR _14953_/X sky130_fd_sc_hd__and3_4
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18477__A _16941_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20800__A _22461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21925__A1 _21865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21925__B2 _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13904_ _13916_/A _23677_/Q VGND VGND VPWR VPWR _13904_/X sky130_fd_sc_hd__or2_4
XFILLER_47_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17672_ _17669_/X VGND VGND VPWR VPWR _17672_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14884_ _14881_/A _14884_/B VGND VGND VPWR VPWR _14884_/X sky130_fd_sc_hd__or2_4
XFILLER_130_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16623_ _16656_/A _16621_/X _16623_/C VGND VGND VPWR VPWR _16623_/X sky130_fd_sc_hd__and3_4
X_19411_ _19406_/X VGND VGND VPWR VPWR _19411_/X sky130_fd_sc_hd__buf_2
XFILLER_62_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21088__A2_N _21087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13835_ _14319_/A _24061_/Q VGND VGND VPWR VPWR _13835_/X sky130_fd_sc_hd__or2_4
XFILLER_28_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13414__A _13414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16554_ _12015_/A VGND VGND VPWR VPWR _16554_/X sky130_fd_sc_hd__buf_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19342_ _19340_/X _18066_/X _19340_/X _24271_/Q VGND VGND VPWR VPWR _24271_/D sky130_fd_sc_hd__a2bb2o_4
X_13766_ _13742_/A _13766_/B VGND VGND VPWR VPWR _13766_/X sky130_fd_sc_hd__or2_4
XANTENNA__21153__A2 _21148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15505_ _12626_/A _15505_/B VGND VGND VPWR VPWR _15505_/X sky130_fd_sc_hd__or2_4
XFILLER_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21631__A _21624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12717_ _13339_/A _12692_/X _12699_/X _12708_/X _12716_/X VGND VGND VPWR VPWR _12717_/X
+ sky130_fd_sc_hd__a32o_4
X_19273_ _19250_/B VGND VGND VPWR VPWR _19273_/Y sky130_fd_sc_hd__inv_2
X_16485_ _16166_/X _16409_/B VGND VGND VPWR VPWR _16485_/X sky130_fd_sc_hd__or2_4
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13697_ _13697_/A VGND VGND VPWR VPWR _14543_/A sky130_fd_sc_hd__buf_2
X_18224_ _18282_/A _17469_/A VGND VGND VPWR VPWR _18224_/X sky130_fd_sc_hd__and2_4
X_15436_ _13675_/A _15508_/B VGND VGND VPWR VPWR _15438_/B sky130_fd_sc_hd__or2_4
X_12648_ _12953_/A _12648_/B _12648_/C VGND VGND VPWR VPWR _12649_/C sky130_fd_sc_hd__and3_4
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20247__A _16918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22102__B2 _22094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18155_ _18283_/A _18155_/B _18155_/C _18155_/D VGND VGND VPWR VPWR _18156_/A sky130_fd_sc_hd__or4_4
XANTENNA__11869__A _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15367_ _12580_/A _23864_/Q VGND VGND VPWR VPWR _15367_/X sky130_fd_sc_hd__or2_4
X_12579_ _12955_/A _12579_/B VGND VGND VPWR VPWR _12579_/X sky130_fd_sc_hd__or2_4
XANTENNA__22653__A2 _22651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17106_ _17197_/A VGND VGND VPWR VPWR _17144_/A sky130_fd_sc_hd__buf_2
X_14318_ _15406_/A _23484_/Q VGND VGND VPWR VPWR _14320_/B sky130_fd_sc_hd__or2_4
XFILLER_171_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18086_ _17833_/A _17241_/X _17876_/X _18085_/X VGND VGND VPWR VPWR _18086_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_112_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR _23229_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15298_ _12453_/A _24088_/Q VGND VGND VPWR VPWR _15299_/C sky130_fd_sc_hd__or2_4
XANTENNA__22462__A _22462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17037_ _17048_/A VGND VGND VPWR VPWR _17037_/Y sky130_fd_sc_hd__inv_2
X_14249_ _12336_/A _14249_/B _14248_/X VGND VGND VPWR VPWR _14249_/X sky130_fd_sc_hd__and3_4
XANTENNA__17556__A _16309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15076__A _15076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18988_ _24366_/Q _11540_/B _18981_/Y VGND VGND VPWR VPWR _18988_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_100_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17939_ _18126_/A _17937_/X _17850_/X _17938_/X VGND VGND VPWR VPWR _17940_/A sky130_fd_sc_hd__o22a_4
XFILLER_22_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17291__A _17290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20950_ _20755_/X _20949_/X _11518_/A _20269_/A VGND VGND VPWR VPWR _20950_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21392__A2 _21391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18793__B1 _24466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19609_ HRDATA[27] VGND VGND VPWR VPWR _20380_/B sky130_fd_sc_hd__buf_2
XFILLER_26_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20881_ _20726_/X _20880_/Y _24283_/Q _20347_/X VGND VGND VPWR VPWR _20881_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22620_ _22456_/X _22615_/X _15546_/B _22619_/X VGND VGND VPWR VPWR _23169_/D sky130_fd_sc_hd__o22a_4
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17348__A1 _15252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21144__A2 _21141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18834__B _18888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22551_ _22558_/A VGND VGND VPWR VPWR _22551_/X sky130_fd_sc_hd__buf_2
XFILLER_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16635__A _16635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21502_ _21285_/X _21499_/X _15502_/B _21496_/X VGND VGND VPWR VPWR _23810_/D sky130_fd_sc_hd__o22a_4
XFILLER_167_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22482_ _22482_/A VGND VGND VPWR VPWR _22482_/X sky130_fd_sc_hd__buf_2
XFILLER_50_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20157__A _20157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24221_ _24248_/CLK _19424_/X HRESETn VGND VGND VPWR VPWR _24221_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11779__A _15362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21433_ _21254_/X _21427_/X _16287_/B _21431_/X VGND VGND VPWR VPWR _21433_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19946__A _24129_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18848__A1 _16523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14582__A1 _13689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24152_ _24302_/CLK _20030_/Y HRESETn VGND VGND VPWR VPWR _18190_/A sky130_fd_sc_hd__dfrtp_4
X_21364_ _21307_/X _21362_/X _14736_/B _21359_/X VGND VGND VPWR VPWR _23897_/D sky130_fd_sc_hd__o22a_4
X_20315_ _20315_/A VGND VGND VPWR VPWR _20315_/X sky130_fd_sc_hd__buf_2
X_23103_ _23582_/CLK _23103_/D VGND VGND VPWR VPWR _23103_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14334__A1 _11854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17466__A _17156_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14334__B2 _14333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24083_ _23889_/CLK _24083_/D VGND VGND VPWR VPWR _24083_/Q sky130_fd_sc_hd__dfxtp_4
X_21295_ _20819_/A VGND VGND VPWR VPWR _21295_/X sky130_fd_sc_hd__buf_2
XANTENNA__16370__A _13392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20246_ _20871_/A _20246_/B VGND VGND VPWR VPWR _20247_/D sky130_fd_sc_hd__or2_4
X_23034_ _23007_/X _17703_/A _23019_/X _23033_/X VGND VGND VPWR VPWR _23035_/A sky130_fd_sc_hd__a211o_4
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_17_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20177_ _20157_/Y _20158_/Y _11571_/X _20176_/X VGND VGND VPWR VPWR _20177_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12403__A _12373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24481__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21907__B2 _21906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15714__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11950_ _16116_/A VGND VGND VPWR VPWR _11951_/A sky130_fd_sc_hd__buf_2
X_23936_ _23744_/CLK _23936_/D VGND VGND VPWR VPWR _14035_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21383__A2 _21377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22580__B2 _22576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11881_ _11881_/A VGND VGND VPWR VPWR _13318_/A sky130_fd_sc_hd__buf_2
XANTENNA__20591__B1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23867_ _23515_/CLK _23867_/D VGND VGND VPWR VPWR _14477_/B sky130_fd_sc_hd__dfxtp_4
X_13620_ _15401_/A _13618_/X _13619_/X VGND VGND VPWR VPWR _13620_/X sky130_fd_sc_hd__and3_4
XFILLER_44_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22818_ _22817_/X VGND VGND VPWR VPWR _22818_/X sky130_fd_sc_hd__buf_2
X_23798_ _23862_/CLK _23798_/D VGND VGND VPWR VPWR _14967_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13551_ _13535_/A _13477_/B VGND VGND VPWR VPWR _13552_/C sky130_fd_sc_hd__or2_4
XFILLER_38_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22749_ _22773_/A VGND VGND VPWR VPWR _22749_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16545__A _12001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12502_ _12502_/A VGND VGND VPWR VPWR _12503_/A sky130_fd_sc_hd__buf_2
XFILLER_160_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16270_ _16096_/A _16270_/B VGND VGND VPWR VPWR _16270_/X sky130_fd_sc_hd__or2_4
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13482_ _12874_/A _13478_/X _13482_/C VGND VGND VPWR VPWR _13483_/B sky130_fd_sc_hd__or3_4
XFILLER_9_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15221_ _14631_/A _15221_/B _15220_/X VGND VGND VPWR VPWR _15225_/B sky130_fd_sc_hd__and3_4
XFILLER_139_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12433_ _12433_/A VGND VGND VPWR VPWR _12434_/A sky130_fd_sc_hd__buf_2
X_24419_ _24419_/CLK _24419_/D HRESETn VGND VGND VPWR VPWR _20677_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22635__A2 _22608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14065__A _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15152_ _15022_/A _15152_/B _15151_/X VGND VGND VPWR VPWR _15152_/X sky130_fd_sc_hd__or3_4
X_12364_ _12363_/X _12259_/B VGND VGND VPWR VPWR _12364_/X sky130_fd_sc_hd__or2_4
XANTENNA__24213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19575__B HRDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14103_ _14103_/A _14101_/X _14103_/C VGND VGND VPWR VPWR _14107_/B sky130_fd_sc_hd__and3_4
XFILLER_4_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19960_ _18623_/Y _20150_/A VGND VGND VPWR VPWR _19960_/X sky130_fd_sc_hd__or2_4
X_15083_ _14682_/A _15074_/X _15083_/C VGND VGND VPWR VPWR _15084_/C sky130_fd_sc_hd__and3_4
XFILLER_153_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12295_ _12304_/A VGND VGND VPWR VPWR _13184_/A sky130_fd_sc_hd__buf_2
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22399__B2 _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18911_ _12419_/X _18906_/X _24396_/Q _18907_/X VGND VGND VPWR VPWR _24396_/D sky130_fd_sc_hd__o22a_4
X_14034_ _11680_/A _14024_/X _14034_/C VGND VGND VPWR VPWR _14050_/B sky130_fd_sc_hd__and3_4
X_19891_ _19889_/X _19890_/X _19903_/A VGND VGND VPWR VPWR _19891_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_136_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13409__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21071__B2 _21070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18842_ _18842_/A VGND VGND VPWR VPWR _18843_/A sky130_fd_sc_hd__buf_2
XFILLER_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12313__A _13183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15985_ _15960_/A _24078_/Q VGND VGND VPWR VPWR _15986_/C sky130_fd_sc_hd__or2_4
XFILLER_121_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18773_ _18773_/A _18773_/B _18772_/X VGND VGND VPWR VPWR _18774_/A sky130_fd_sc_hd__and3_4
XANTENNA__20530__A _20530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22020__B1 _15455_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17724_ _18533_/A _17427_/X _17723_/Y VGND VGND VPWR VPWR _17724_/X sky130_fd_sc_hd__a21o_4
X_14936_ _14772_/A VGND VGND VPWR VPWR _14976_/A sky130_fd_sc_hd__buf_2
XFILLER_48_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22571__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14867_ _14108_/A _14867_/B VGND VGND VPWR VPWR _14867_/X sky130_fd_sc_hd__or2_4
X_17655_ _17655_/A _17252_/Y VGND VGND VPWR VPWR _17655_/X sky130_fd_sc_hd__and2_4
XFILLER_91_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13144__A _13164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_37_0_HCLK clkbuf_7_37_0_HCLK/A VGND VGND VPWR VPWR _23761_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16606_ _16606_/A VGND VGND VPWR VPWR _16675_/A sky130_fd_sc_hd__buf_2
XFILLER_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13818_ _13658_/A _13818_/B VGND VGND VPWR VPWR _13818_/X sky130_fd_sc_hd__or2_4
X_17586_ _17140_/Y _18076_/B VGND VGND VPWR VPWR _17586_/X sky130_fd_sc_hd__or2_4
XANTENNA__21126__A2 _21125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14798_ _14691_/A _14798_/B VGND VGND VPWR VPWR _14800_/B sky130_fd_sc_hd__or2_4
XFILLER_44_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22457__A _22433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19325_ _19428_/A VGND VGND VPWR VPWR _19325_/X sky130_fd_sc_hd__buf_2
X_16537_ _11951_/X _16535_/X _16536_/X VGND VGND VPWR VPWR _16542_/B sky130_fd_sc_hd__and3_4
X_13749_ _13229_/A _13749_/B _13749_/C VGND VGND VPWR VPWR _13749_/X sky130_fd_sc_hd__or3_4
XFILLER_56_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12983__A _12914_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20885__A1 _18643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16468_ _16491_/A _16398_/B VGND VGND VPWR VPWR _16468_/X sky130_fd_sc_hd__or2_4
X_19256_ _24307_/Q _19256_/B VGND VGND VPWR VPWR _19258_/A sky130_fd_sc_hd__and2_4
XFILLER_148_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11599__A _17357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24354__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18207_ _18389_/A _18172_/X _18206_/X _18167_/B VGND VGND VPWR VPWR _18207_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22087__B1 _23477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15419_ _11932_/A _15415_/X _15419_/C VGND VGND VPWR VPWR _15419_/X sky130_fd_sc_hd__or3_4
X_19187_ _19149_/B VGND VGND VPWR VPWR _19187_/Y sky130_fd_sc_hd__inv_2
X_16399_ _15998_/X _16399_/B _16399_/C VGND VGND VPWR VPWR _16399_/X sky130_fd_sc_hd__and3_4
XANTENNA__18670__A _18670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__22904__B _19953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18138_ _18138_/A _18137_/X VGND VGND VPWR VPWR _18138_/Y sky130_fd_sc_hd__nand2_4
XFILLER_129_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17502__A1 _13342_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17502__B2 _17501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18069_ _17900_/X _18067_/X _20003_/A _18068_/X VGND VGND VPWR VPWR _24495_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20100_ _18624_/X _18620_/X _20099_/X VGND VGND VPWR VPWR _20100_/X sky130_fd_sc_hd__o21a_4
XFILLER_144_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21080_ _21080_/A VGND VGND VPWR VPWR _21080_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15518__B _15517_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14422__B _14485_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20031_ _19961_/X VGND VGND VPWR VPWR _20031_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21062__B2 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12223__A _12721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20440__A _22110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15534__A _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21982_ _21874_/X _21981_/X _23546_/Q _21978_/X VGND VGND VPWR VPWR _21982_/X sky130_fd_sc_hd__o22a_4
XFILLER_113_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21365__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23721_ _23337_/CLK _21678_/X VGND VGND VPWR VPWR _23721_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20933_ _20639_/A _20921_/X _20779_/X _20932_/Y VGND VGND VPWR VPWR _20933_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15253__B _15253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13054__A _13094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ _23523_/CLK _23652_/D VGND VGND VPWR VPWR _15705_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ _20864_/A VGND VGND VPWR VPWR _20864_/X sky130_fd_sc_hd__buf_2
XANTENNA__21117__A2 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22314__B2 _22312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22603_ _22428_/X _22601_/X _16193_/B _22598_/X VGND VGND VPWR VPWR _23181_/D sky130_fd_sc_hd__o22a_4
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12893__A _12889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23583_ _23582_/CLK _23583_/D VGND VGND VPWR VPWR _23583_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20795_ _20794_/X VGND VGND VPWR VPWR _20795_/Y sky130_fd_sc_hd__inv_2
X_22534_ _22482_/X _22529_/X _23222_/Q _22498_/A VGND VGND VPWR VPWR _22534_/X sky130_fd_sc_hd__o22a_4
X_22465_ _22464_/X _22462_/X _13702_/B _22457_/X VGND VGND VPWR VPWR _22465_/X sky130_fd_sc_hd__o22a_4
XFILLER_124_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20628__A1 _20234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24204_ _23671_/CLK _19701_/X HRESETn VGND VGND VPWR VPWR _11603_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_147_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21416_ _21311_/X _21412_/X _15180_/B _21381_/A VGND VGND VPWR VPWR _23863_/D sky130_fd_sc_hd__o22a_4
XFILLER_33_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22396_ _22156_/X _22390_/X _14495_/B _22394_/X VGND VGND VPWR VPWR _22396_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24135_ _24134_/CLK _24135_/D HRESETn VGND VGND VPWR VPWR _24135_/Q sky130_fd_sc_hd__dfrtp_4
X_21347_ _21278_/X _21341_/X _23909_/Q _21345_/X VGND VGND VPWR VPWR _23909_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15709__A _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24066_ _23587_/CLK _24066_/D VGND VGND VPWR VPWR _15490_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12080_ _12041_/A _23987_/Q VGND VGND VPWR VPWR _12081_/C sky130_fd_sc_hd__or2_4
X_21278_ _21848_/A VGND VGND VPWR VPWR _21278_/X sky130_fd_sc_hd__buf_2
XFILLER_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23871__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21053__B2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13229__A _13229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23017_ _23007_/X _17686_/A _22989_/X _23016_/X VGND VGND VPWR VPWR _23018_/A sky130_fd_sc_hd__a211o_4
X_20229_ _20229_/A VGND VGND VPWR VPWR _20229_/X sky130_fd_sc_hd__buf_2
XFILLER_103_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18770__A1_N _17100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11972__A _11971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15444__A _15444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19549__A2 _19848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23101__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15770_ _15770_/A _23716_/Q VGND VGND VPWR VPWR _15772_/B sky130_fd_sc_hd__or2_4
XANTENNA__24227__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12982_ _12983_/B VGND VGND VPWR VPWR _12982_/X sky130_fd_sc_hd__buf_2
XANTENNA__23083__D _23083_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21356__A2 _21355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22553__B2 _22548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14721_ _12503_/A _14721_/B VGND VGND VPWR VPWR _14722_/C sky130_fd_sc_hd__or2_4
XFILLER_85_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23919_ _23983_/CLK _23919_/D VGND VGND VPWR VPWR _16279_/B sky130_fd_sc_hd__dfxtp_4
X_11933_ _11933_/A VGND VGND VPWR VPWR _12266_/A sky130_fd_sc_hd__buf_2
XANTENNA__15163__B _15227_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17440_ _17436_/B _17438_/X _17439_/X VGND VGND VPWR VPWR _17440_/X sky130_fd_sc_hd__o21a_4
X_14652_ _15625_/A _14646_/X _14651_/X VGND VGND VPWR VPWR _14652_/X sky130_fd_sc_hd__or3_4
X_11864_ _11864_/A VGND VGND VPWR VPWR _13483_/A sky130_fd_sc_hd__buf_2
XANTENNA__22277__A _22284_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _11912_/A VGND VGND VPWR VPWR _15415_/A sky130_fd_sc_hd__buf_2
XPHY_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _17371_/A VGND VGND VPWR VPWR _17375_/A sky130_fd_sc_hd__inv_2
XANTENNA__13899__A _13888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _14278_/A _14583_/B VGND VGND VPWR VPWR _14583_/X sky130_fd_sc_hd__or2_4
XANTENNA__24465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16275__A _11882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11795_ _11836_/A _11795_/B VGND VGND VPWR VPWR _11796_/C sky130_fd_sc_hd__or2_4
XFILLER_25_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16322_ _16195_/A _16257_/B VGND VGND VPWR VPWR _16323_/C sky130_fd_sc_hd__or2_4
X_19110_ _11519_/A _11519_/B _11519_/X VGND VGND VPWR VPWR _19110_/Y sky130_fd_sc_hd__a21boi_4
X_13534_ _13534_/A _23621_/Q VGND VGND VPWR VPWR _13536_/B sky130_fd_sc_hd__or2_4
XFILLER_158_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19041_ _11530_/X VGND VGND VPWR VPWR _19041_/Y sky130_fd_sc_hd__inv_2
X_16253_ _16287_/A _16253_/B VGND VGND VPWR VPWR _16253_/X sky130_fd_sc_hd__or2_4
XANTENNA__22069__B1 _15833_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13465_ _13441_/A _23397_/Q VGND VGND VPWR VPWR _13465_/X sky130_fd_sc_hd__or2_4
XFILLER_146_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15204_ _15198_/X _15147_/B VGND VGND VPWR VPWR _15204_/X sky130_fd_sc_hd__or2_4
X_12416_ _13564_/A _12416_/B _12416_/C VGND VGND VPWR VPWR _12417_/C sky130_fd_sc_hd__and3_4
X_16184_ _16231_/A _23309_/Q VGND VGND VPWR VPWR _16184_/X sky130_fd_sc_hd__or2_4
X_13396_ _13408_/A _23398_/Q VGND VGND VPWR VPWR _13396_/X sky130_fd_sc_hd__or2_4
XFILLER_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15135_ _14994_/A VGND VGND VPWR VPWR _15294_/A sky130_fd_sc_hd__buf_2
X_12347_ _12604_/A VGND VGND VPWR VPWR _13235_/A sky130_fd_sc_hd__buf_2
XFILLER_127_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19943_ _19938_/X _24166_/Q _19939_/X _19773_/X VGND VGND VPWR VPWR _19943_/X sky130_fd_sc_hd__o22a_4
X_15066_ _14841_/A _15058_/X _15065_/X VGND VGND VPWR VPWR _15066_/X sky130_fd_sc_hd__and3_4
X_12278_ _12698_/A _12276_/X _12277_/X VGND VGND VPWR VPWR _12278_/X sky130_fd_sc_hd__and3_4
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19360__A2_N _18450_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14017_ _15369_/A VGND VGND VPWR VPWR _14074_/A sky130_fd_sc_hd__buf_2
XANTENNA__21044__B2 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19874_ _19749_/X _19868_/B _19643_/A _19868_/B VGND VGND VPWR VPWR _19874_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12043__A _16561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18825_ _18789_/A VGND VGND VPWR VPWR _18825_/X sky130_fd_sc_hd__buf_2
XANTENNA__12978__A _12978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11882__A _13318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15354__A _11752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18756_ _18413_/A _18755_/X VGND VGND VPWR VPWR _18756_/Y sky130_fd_sc_hd__nor2_4
X_15968_ _15959_/A VGND VGND VPWR VPWR _15969_/A sky130_fd_sc_hd__buf_2
XANTENNA__21347__A2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14482__B1 _11606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17707_ _17708_/A _17381_/X VGND VGND VPWR VPWR _17711_/A sky130_fd_sc_hd__or2_4
X_14919_ _14919_/A _23734_/Q VGND VGND VPWR VPWR _14920_/C sky130_fd_sc_hd__or2_4
XFILLER_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15899_ _13543_/X _15843_/B VGND VGND VPWR VPWR _15899_/X sky130_fd_sc_hd__or2_4
X_18687_ _18413_/X _17628_/X _18467_/X _17348_/X VGND VGND VPWR VPWR _18687_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_91_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17638_ _17638_/A VGND VGND VPWR VPWR _17638_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22187__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17569_ _17139_/X _18076_/B VGND VGND VPWR VPWR _17569_/X sky130_fd_sc_hd__and2_4
XANTENNA__22278__A2_N _22277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13602__A _14448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19308_ _24283_/Q _19231_/X _19307_/Y VGND VGND VPWR VPWR _19308_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24135__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20580_ _11573_/A VGND VGND VPWR VPWR _20581_/A sky130_fd_sc_hd__inv_2
XFILLER_165_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19239_ _24290_/Q _19295_/A VGND VGND VPWR VPWR _19240_/B sky130_fd_sc_hd__and2_4
XFILLER_143_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12218__A _12218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22250_ _22132_/X _22244_/X _23397_/Q _22248_/X VGND VGND VPWR VPWR _23397_/D sky130_fd_sc_hd__o22a_4
XFILLER_30_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21201_ _20486_/X _21198_/X _23980_/Q _21195_/X VGND VGND VPWR VPWR _21201_/X sky130_fd_sc_hd__o22a_4
X_22181_ _22097_/X _22180_/X _12159_/B _22177_/X VGND VGND VPWR VPWR _23443_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14433__A _12455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21132_ _24020_/Q VGND VGND VPWR VPWR _21132_/Y sky130_fd_sc_hd__inv_2
X_21063_ _21049_/A VGND VGND VPWR VPWR _21063_/X sky130_fd_sc_hd__buf_2
XFILLER_8_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21586__A2 _21578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20014_ _19992_/X _17667_/A _19998_/X _20013_/X VGND VGND VPWR VPWR _20014_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21266__A _20531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17463__B _17481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12888__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11792__A _11768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22535__B2 _22498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21965_ _21845_/X _21960_/X _13297_/B _21964_/X VGND VGND VPWR VPWR _23558_/D sky130_fd_sc_hd__o22a_4
XFILLER_70_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _23770_/CLK _23704_/D VGND VGND VPWR VPWR _15307_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _20894_/X _20915_/X _14598_/B _20861_/X VGND VGND VPWR VPWR _20916_/X sky130_fd_sc_hd__o22a_4
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21896_ _21813_/X _21895_/X _23603_/Q _21892_/X VGND VGND VPWR VPWR _21896_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22097__A _20336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_20_0_HCLK clkbuf_6_10_0_HCLK/X VGND VGND VPWR VPWR _24127_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23889_/CLK _23635_/D VGND VGND VPWR VPWR _23635_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _20847_/A VGND VGND VPWR VPWR _21017_/A sky130_fd_sc_hd__buf_2
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16095__A _12559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14608__A _13655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_83_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR _23864_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20329__B _20329_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23566_ _24078_/CLK _21954_/X VGND VGND VPWR VPWR _23566_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11580_ _24468_/Q IRQ[31] VGND VGND VPWR VPWR _20124_/A sky130_fd_sc_hd__and2_4
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20778_ _20778_/A _20777_/X VGND VGND VPWR VPWR _20778_/X sky130_fd_sc_hd__or2_4
XFILLER_11_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13231__B _23975_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22517_ _22452_/X _22515_/X _15836_/B _22512_/X VGND VGND VPWR VPWR _23235_/D sky130_fd_sc_hd__o22a_4
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23497_ _23561_/CLK _23497_/D VGND VGND VPWR VPWR _23497_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13250_ _12338_/X _13250_/B _13250_/C VGND VGND VPWR VPWR _13251_/C sky130_fd_sc_hd__and3_4
X_22448_ _22447_/X _22438_/X _23269_/Q _22445_/X VGND VGND VPWR VPWR _23269_/D sky130_fd_sc_hd__o22a_4
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12201_ _11881_/A _12201_/B _12201_/C VGND VGND VPWR VPWR _12208_/B sky130_fd_sc_hd__and3_4
XANTENNA__15439__A _15439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13181_ _12741_/A _13181_/B _13181_/C VGND VGND VPWR VPWR _13181_/X sky130_fd_sc_hd__and3_4
XANTENNA__21274__B2 _21264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21425__A2_N _21424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22379_ _22127_/X _22376_/X _13208_/B _22373_/X VGND VGND VPWR VPWR _22379_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14343__A _14519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12132_ _12127_/A _23955_/Q VGND VGND VPWR VPWR _12134_/B sky130_fd_sc_hd__or2_4
X_24118_ _23991_/CLK _24118_/D HRESETn VGND VGND VPWR VPWR _22773_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24049_ _23761_/CLK _24049_/D VGND VGND VPWR VPWR _24049_/Q sky130_fd_sc_hd__dfxtp_4
X_16940_ _16939_/X VGND VGND VPWR VPWR _16940_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12063_ _12058_/A _12142_/B VGND VGND VPWR VPWR _12063_/X sky130_fd_sc_hd__or2_4
XFILLER_81_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14997__B _23285_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21176__A _21136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16871_ _15388_/X VGND VGND VPWR VPWR _16871_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12798__A _13343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18610_ _17980_/X _18130_/Y _17869_/A _18609_/Y VGND VGND VPWR VPWR _18610_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15174__A _13593_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15822_ _12884_/A _15822_/B VGND VGND VPWR VPWR _15824_/B sky130_fd_sc_hd__or2_4
XFILLER_18_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19590_ _24168_/Q _19457_/X HRDATA[20] _19454_/X VGND VGND VPWR VPWR _19590_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21329__A2 _21327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15753_ _12762_/A _15688_/B VGND VGND VPWR VPWR _15754_/C sky130_fd_sc_hd__or2_4
X_18541_ _17435_/Y _18539_/X VGND VGND VPWR VPWR _18541_/X sky130_fd_sc_hd__or2_4
X_12965_ _12941_/A _12965_/B _12965_/C VGND VGND VPWR VPWR _12965_/X sky130_fd_sc_hd__and3_4
XFILLER_166_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18485__A _18485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11916_ _12870_/A VGND VGND VPWR VPWR _12515_/A sky130_fd_sc_hd__buf_2
X_14704_ _14613_/X _14701_/Y VGND VGND VPWR VPWR _14704_/X sky130_fd_sc_hd__and2_4
X_15684_ _12858_/A _15680_/X _15683_/X VGND VGND VPWR VPWR _15684_/X sky130_fd_sc_hd__or3_4
X_18472_ _18458_/X _18463_/Y _18465_/X _18470_/X _18471_/Y VGND VGND VPWR VPWR _18472_/X
+ sky130_fd_sc_hd__a32o_4
X_12896_ _12873_/A _12896_/B _12895_/X VGND VGND VPWR VPWR _12897_/C sky130_fd_sc_hd__and3_4
X_17423_ _17423_/A _17423_/B VGND VGND VPWR VPWR _17635_/A sky130_fd_sc_hd__or2_4
X_14635_ _14635_/A VGND VGND VPWR VPWR _14685_/A sky130_fd_sc_hd__buf_2
X_11847_ _16635_/A _11845_/X _11846_/X VGND VGND VPWR VPWR _11847_/X sky130_fd_sc_hd__and3_4
XFILLER_159_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14518__A _12401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13422__A _13455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20239__B HRDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17019_/X VGND VGND VPWR VPWR _17354_/X sky130_fd_sc_hd__buf_2
X_14566_ _14310_/A _14562_/X _14565_/X VGND VGND VPWR VPWR _14566_/X sky130_fd_sc_hd__or3_4
X_11778_ _11663_/A VGND VGND VPWR VPWR _15362_/A sky130_fd_sc_hd__inv_2
XANTENNA__21501__A2 _21499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13517_ _12971_/A VGND VGND VPWR VPWR _13554_/A sky130_fd_sc_hd__buf_2
X_16305_ _11917_/X _16303_/X _16305_/C VGND VGND VPWR VPWR _16305_/X sky130_fd_sc_hd__and3_4
XFILLER_119_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17285_ _11611_/C VGND VGND VPWR VPWR _17285_/Y sky130_fd_sc_hd__inv_2
X_14497_ _14522_/A _14493_/X _14497_/C VGND VGND VPWR VPWR _14497_/X sky130_fd_sc_hd__or3_4
XANTENNA__16733__A _16561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16236_ _16214_/A _16236_/B _16236_/C VGND VGND VPWR VPWR _16237_/C sky130_fd_sc_hd__or3_4
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19024_ _19024_/A VGND VGND VPWR VPWR _19024_/X sky130_fd_sc_hd__buf_2
XFILLER_173_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13448_ _12886_/A _13446_/X _13447_/X VGND VGND VPWR VPWR _13448_/X sky130_fd_sc_hd__and3_4
XFILLER_174_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20255__A _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21265__B2 _21264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16167_ _16166_/X _16167_/B VGND VGND VPWR VPWR _16168_/C sky130_fd_sc_hd__or2_4
XFILLER_155_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13379_ _13379_/A _13297_/B VGND VGND VPWR VPWR _13380_/C sky130_fd_sc_hd__or2_4
XANTENNA__14253__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15118_ _14983_/A VGND VGND VPWR VPWR _15118_/X sky130_fd_sc_hd__buf_2
XFILLER_173_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16098_ _16108_/A _23373_/Q VGND VGND VPWR VPWR _16103_/B sky130_fd_sc_hd__or2_4
XFILLER_141_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15068__B _23573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19926_ _24179_/Q _19921_/X _20246_/B _19925_/X VGND VGND VPWR VPWR _24179_/D sky130_fd_sc_hd__o22a_4
X_15049_ _14771_/A VGND VGND VPWR VPWR _15078_/A sky130_fd_sc_hd__buf_2
XANTENNA__22214__B1 _14463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21086__A _21101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19857_ _19899_/A _19857_/B VGND VGND VPWR VPWR _19857_/X sky130_fd_sc_hd__or2_4
XANTENNA__15084__A _11674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18808_ _13262_/X _18803_/X _11573_/A _18804_/X VGND VGND VPWR VPWR _18808_/X sky130_fd_sc_hd__o22a_4
X_19788_ _19788_/A _19807_/A VGND VGND VPWR VPWR _19788_/X sky130_fd_sc_hd__and2_4
XFILLER_56_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22517__B2 _22512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21814__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18739_ _18738_/X VGND VGND VPWR VPWR _22846_/B sky130_fd_sc_hd__inv_2
XFILLER_23_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15812__A _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21750_ _21592_/X _21748_/X _14720_/B _21745_/X VGND VGND VPWR VPWR _21750_/X sky130_fd_sc_hd__o22a_4
XFILLER_92_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21740__A2 _21734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20701_ _20641_/X _20700_/X _20639_/X VGND VGND VPWR VPWR _20701_/Y sky130_fd_sc_hd__o21ai_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21681_ _21674_/A VGND VGND VPWR VPWR _21681_/X sky130_fd_sc_hd__buf_2
XANTENNA__14428__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23420_ _23772_/CLK _23420_/D VGND VGND VPWR VPWR _14392_/B sky130_fd_sc_hd__dfxtp_4
X_20632_ _20632_/A VGND VGND VPWR VPWR _21848_/A sky130_fd_sc_hd__buf_2
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23351_ _23511_/CLK _23351_/D VGND VGND VPWR VPWR _15125_/B sky130_fd_sc_hd__dfxtp_4
X_20563_ _24424_/Q _20427_/X _24456_/Q _20471_/X VGND VGND VPWR VPWR _20563_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22302_ _22134_/X _22301_/X _15660_/B _22298_/X VGND VGND VPWR VPWR _22302_/X sky130_fd_sc_hd__o22a_4
XFILLER_109_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19449__A1 HRDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23282_ _23537_/CLK _23282_/D VGND VGND VPWR VPWR _16609_/B sky130_fd_sc_hd__dfxtp_4
X_20494_ _20494_/A _20494_/B VGND VGND VPWR VPWR _20494_/X sky130_fd_sc_hd__or2_4
XANTENNA__22453__B1 _15789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11787__A _11742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15259__A _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22233_ _22103_/X _22230_/X _16798_/B _22227_/X VGND VGND VPWR VPWR _23409_/D sky130_fd_sc_hd__o22a_4
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14163__A _13791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22164_ _22163_/X _22159_/X _23448_/Q _22154_/X VGND VGND VPWR VPWR _23448_/D sky130_fd_sc_hd__o22a_4
XFILLER_133_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22380__A _22358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21115_ _21101_/A VGND VGND VPWR VPWR _21115_/X sky130_fd_sc_hd__buf_2
XFILLER_161_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22095_ _20298_/A VGND VGND VPWR VPWR _22095_/X sky130_fd_sc_hd__buf_2
XANTENNA__21559__A2 _21554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21046_ _20441_/X _21045_/X _24078_/Q _21042_/X VGND VGND VPWR VPWR _24078_/D sky130_fd_sc_hd__o22a_4
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21724__A _21724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22997_ _22978_/X _22995_/X _22997_/C VGND VGND VPWR VPWR _22997_/X sky130_fd_sc_hd__and3_4
XFILLER_28_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16818__A _16684_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12750_ _11864_/A _12749_/X VGND VGND VPWR VPWR _12750_/X sky130_fd_sc_hd__and2_4
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21948_ _21817_/X _21946_/X _23570_/Q _21943_/X VGND VGND VPWR VPWR _21948_/X sky130_fd_sc_hd__o22a_4
XFILLER_83_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11701_/A VGND VGND VPWR VPWR _13367_/A sky130_fd_sc_hd__buf_2
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12681_ _12574_/X _12679_/Y VGND VGND VPWR VPWR _12682_/A sky130_fd_sc_hd__or2_4
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21879_ _20959_/A VGND VGND VPWR VPWR _21879_/X sky130_fd_sc_hd__buf_2
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14338__A _14377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13242__A _12338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/A _14484_/B VGND VGND VPWR VPWR _14420_/X sky130_fd_sc_hd__or2_4
X_11632_ _11631_/X VGND VGND VPWR VPWR _11632_/X sky130_fd_sc_hd__buf_2
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _23587_/CLK _23618_/D VGND VGND VPWR VPWR _15489_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19688__A1 _19797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _12401_/A _14349_/X _14350_/X VGND VGND VPWR VPWR _14351_/X sky130_fd_sc_hd__and3_4
XANTENNA__21495__B2 _21489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23549_ _23679_/CLK _23549_/D VGND VGND VPWR VPWR _13819_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ _20159_/A IRQ[15] _11562_/X VGND VGND VPWR VPWR _11563_/X sky130_fd_sc_hd__a21o_4
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13276_/A _13302_/B _13301_/X VGND VGND VPWR VPWR _13302_/X sky130_fd_sc_hd__and3_4
XFILLER_128_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11983__A1 _11868_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17070_ _17070_/A _17070_/B _17069_/X VGND VGND VPWR VPWR _17070_/X sky130_fd_sc_hd__and3_4
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _13601_/A _14355_/B VGND VGND VPWR VPWR _14282_/X sky130_fd_sc_hd__or2_4
X_16021_ _16031_/A VGND VGND VPWR VPWR _16061_/A sky130_fd_sc_hd__buf_2
XFILLER_137_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13233_ _13252_/A _23623_/Q VGND VGND VPWR VPWR _13233_/X sky130_fd_sc_hd__or2_4
XANTENNA__15169__A _14295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11697__A _11697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21994__A2_N _21993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18190__D _18148_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14073__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13164_ _13164_/A _23623_/Q VGND VGND VPWR VPWR _13166_/B sky130_fd_sc_hd__or2_4
XFILLER_83_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20803__A HRDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12115_ _16080_/A VGND VGND VPWR VPWR _16775_/A sky130_fd_sc_hd__buf_2
XFILLER_2_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17384__A _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13095_ _13095_/A _23976_/Q VGND VGND VPWR VPWR _13096_/C sky130_fd_sc_hd__or2_4
X_17972_ _17793_/X _17972_/B _17970_/Y _17972_/D VGND VGND VPWR VPWR _17973_/A sky130_fd_sc_hd__or4_4
XANTENNA__22747__B2 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19711_ _19711_/A VGND VGND VPWR VPWR _19712_/B sky130_fd_sc_hd__inv_2
X_16923_ _16915_/X _16920_/X _16922_/X VGND VGND VPWR VPWR _16925_/B sky130_fd_sc_hd__and3_4
X_12046_ _11941_/A VGND VGND VPWR VPWR _16724_/A sky130_fd_sc_hd__buf_2
XFILLER_78_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13417__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19642_ _19642_/A VGND VGND VPWR VPWR _19642_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12321__A _11659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16854_ _13271_/X _16839_/X _13271_/X _16839_/X VGND VGND VPWR VPWR _16858_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21970__A2 _21967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15805_ _12889_/A _15803_/X _15805_/C VGND VGND VPWR VPWR _15805_/X sky130_fd_sc_hd__and3_4
XANTENNA__21634__A _21620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19573_ _19573_/A VGND VGND VPWR VPWR _19573_/X sky130_fd_sc_hd__buf_2
XFILLER_19_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24480__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16785_ _16606_/A _16785_/B _16784_/X VGND VGND VPWR VPWR _16785_/X sky130_fd_sc_hd__or3_4
X_13997_ _13627_/A _23488_/Q VGND VGND VPWR VPWR _13999_/B sky130_fd_sc_hd__or2_4
XANTENNA__18179__B2 _18178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18524_ _18523_/X VGND VGND VPWR VPWR _18524_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15632__A _15616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12948_ _12948_/A _23913_/Q VGND VGND VPWR VPWR _12948_/X sky130_fd_sc_hd__or2_4
X_15736_ _12766_/X _15734_/X _15736_/C VGND VGND VPWR VPWR _15736_/X sky130_fd_sc_hd__and3_4
XFILLER_34_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21722__A2 _21720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18455_ _18367_/A _16981_/X _18433_/Y VGND VGND VPWR VPWR _22979_/B sky130_fd_sc_hd__a21oi_4
X_12879_ _12906_/A _23465_/Q VGND VGND VPWR VPWR _12880_/C sky130_fd_sc_hd__or2_4
X_15667_ _12727_/A _24036_/Q VGND VGND VPWR VPWR _15667_/X sky130_fd_sc_hd__or2_4
XFILLER_61_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17406_ _17251_/A VGND VGND VPWR VPWR _17406_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14618_ _14819_/A _14618_/B VGND VGND VPWR VPWR _14621_/B sky130_fd_sc_hd__or2_4
X_18386_ _18386_/A VGND VGND VPWR VPWR _18411_/B sky130_fd_sc_hd__inv_2
X_15598_ _15612_/A _15596_/X _15597_/X VGND VGND VPWR VPWR _15599_/C sky130_fd_sc_hd__and3_4
XFILLER_159_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21486__B2 _21482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22683__B1 _15162_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17337_ _15117_/Y _17025_/A _17025_/Y _17336_/X VGND VGND VPWR VPWR _17339_/B sky130_fd_sc_hd__o22a_4
X_14549_ _14547_/X VGND VGND VPWR VPWR _14549_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12991__A _12875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18351__B2 _18350_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17268_ _17266_/X _17913_/B VGND VGND VPWR VPWR _17914_/B sky130_fd_sc_hd__or2_4
XFILLER_140_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19007_ _19007_/A VGND VGND VPWR VPWR _19007_/Y sky130_fd_sc_hd__inv_2
X_16219_ _16219_/A _16219_/B VGND VGND VPWR VPWR _16220_/C sky130_fd_sc_hd__or2_4
XANTENNA__15079__A _15103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17199_ _16821_/B _17197_/X _15382_/B _17198_/X VGND VGND VPWR VPWR _17199_/X sky130_fd_sc_hd__o22a_4
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21789__A2 _21784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15807__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14711__A _14297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19909_ _22846_/B VGND VGND VPWR VPWR _19909_/X sky130_fd_sc_hd__buf_2
XFILLER_29_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13327__A _13327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22920_ _23086_/A _22920_/B VGND VGND VPWR VPWR HADDR[3] sky130_fd_sc_hd__nor2_4
XFILLER_111_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21410__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12231__A _12273_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21961__A2 _21960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22851_ _17491_/Y _22847_/X _22884_/A _22850_/X VGND VGND VPWR VPWR _22851_/X sky130_fd_sc_hd__a211o_4
XFILLER_72_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16638__A _16672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15542__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21802_ _21596_/X _21798_/X _15173_/B _21767_/A VGND VGND VPWR VPWR _23639_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22782_ _22781_/A _22781_/B VGND VGND VPWR VPWR _22786_/B sky130_fd_sc_hd__or2_4
XFILLER_83_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13651__A1 _14480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21733_ _21563_/X _21727_/X _23685_/Q _21731_/X VGND VGND VPWR VPWR _23685_/D sky130_fd_sc_hd__o22a_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15261__B _23768_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14158__A _14272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13062__A _13091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24452_ _23475_/CLK _24452_/D HRESETn VGND VGND VPWR VPWR _20159_/A sky130_fd_sc_hd__dfrtp_4
X_21664_ _21528_/X _21663_/X _23731_/Q _21660_/X VGND VGND VPWR VPWR _21664_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23403_ _23558_/CLK _22242_/X VGND VGND VPWR VPWR _12655_/B sky130_fd_sc_hd__dfxtp_4
X_20615_ _20533_/X _20613_/X _24102_/Q _20614_/X VGND VGND VPWR VPWR _20615_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24383_ _24445_/CLK _18930_/X HRESETn VGND VGND VPWR VPWR _19078_/A sky130_fd_sc_hd__dfstp_4
X_21595_ _21594_/X _21590_/X _23768_/Q _21585_/X VGND VGND VPWR VPWR _21595_/X sky130_fd_sc_hd__o22a_4
X_23334_ _23558_/CLK _23334_/D VGND VGND VPWR VPWR _13296_/B sky130_fd_sc_hd__dfxtp_4
X_20546_ _20490_/X _20545_/Y _19246_/A _20323_/X VGND VGND VPWR VPWR _20546_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17188__B _17187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21229__B2 _21223_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23265_ _23203_/CLK _22458_/X VGND VGND VPWR VPWR _15522_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12406__A _15894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20477_ _20343_/X _20476_/X _19153_/A _20352_/X VGND VGND VPWR VPWR _20478_/B sky130_fd_sc_hd__o22a_4
X_22216_ _22158_/X _22215_/X _23418_/Q _22212_/X VGND VGND VPWR VPWR _22216_/X sky130_fd_sc_hd__o22a_4
XFILLER_156_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23196_ _24096_/CLK _23196_/D VGND VGND VPWR VPWR _14349_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22147_ _22147_/A VGND VGND VPWR VPWR _22147_/X sky130_fd_sc_hd__buf_2
XFILLER_161_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22078_ _22057_/A VGND VGND VPWR VPWR _22078_/X sky130_fd_sc_hd__buf_2
XFILLER_94_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20204__A2 _17005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21401__B2 _21395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21029_ _21081_/A _17415_/Y _21234_/B VGND VGND VPWR VPWR _21030_/A sky130_fd_sc_hd__or3_4
X_13920_ _14348_/A _13920_/B _13920_/C VGND VGND VPWR VPWR _13928_/B sky130_fd_sc_hd__or3_4
XANTENNA__24238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21952__A2 _21946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13851_ _11933_/A _13847_/X _13850_/X VGND VGND VPWR VPWR _13851_/X sky130_fd_sc_hd__or3_4
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12802_ _13562_/A _12800_/X _12802_/C VGND VGND VPWR VPWR _12806_/B sky130_fd_sc_hd__and3_4
XANTENNA__11980__A _11951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13782_ _13692_/Y _13781_/X VGND VGND VPWR VPWR _13782_/X sky130_fd_sc_hd__and2_4
X_16570_ _11868_/X _16542_/X _16550_/X _16561_/X _16569_/X VGND VGND VPWR VPWR _16570_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_167_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21704__A2 _21677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22901__B2 _20665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12733_ _12708_/A _12729_/X _12732_/X VGND VGND VPWR VPWR _12733_/X sky130_fd_sc_hd__or3_4
XANTENNA__18030__B1 _18027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15521_ _15518_/X _15520_/Y VGND VGND VPWR VPWR _15521_/X sky130_fd_sc_hd__or2_4
XFILLER_167_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24397__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18581__A1 _17109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18240_ _18064_/X VGND VGND VPWR VPWR _18240_/X sky130_fd_sc_hd__buf_2
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15452_ _11854_/A _11628_/A _15421_/X _11605_/A _15451_/X VGND VGND VPWR VPWR _15453_/A
+ sky130_fd_sc_hd__a32o_4
X_12664_ _12973_/A _12664_/B VGND VGND VPWR VPWR _12664_/X sky130_fd_sc_hd__or2_4
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14510_/A _23484_/Q VGND VGND VPWR VPWR _14405_/B sky130_fd_sc_hd__or2_4
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_53_0_HCLK clkbuf_6_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11928_/A VGND VGND VPWR VPWR _13662_/A sky130_fd_sc_hd__buf_2
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17379__A _17358_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15383_ _15382_/A _15381_/A _15185_/X _15252_/A VGND VGND VPWR VPWR _15384_/A sky130_fd_sc_hd__o22a_4
X_18171_ _17490_/A _18170_/X _17538_/Y VGND VGND VPWR VPWR _18234_/A sky130_fd_sc_hd__o21a_4
XANTENNA__21468__B2 _21431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23805__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12595_ _12659_/A _12585_/X _12595_/C VGND VGND VPWR VPWR _12595_/X sky130_fd_sc_hd__or3_4
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19530__B1 HRDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17122_ _17114_/X _17117_/X _17119_/X _17121_/X VGND VGND VPWR VPWR _17123_/B sky130_fd_sc_hd__o22a_4
XANTENNA__13700__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14334_ _11854_/A _11628_/A _14303_/X _11605_/A _14333_/X VGND VGND VPWR VPWR _14334_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _24442_/Q IRQ[5] _20169_/A VGND VGND VPWR VPWR _11549_/A sky130_fd_sc_hd__a21o_4
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17053_ _12112_/Y _17024_/X _17031_/X _17052_/Y VGND VGND VPWR VPWR _17054_/B sky130_fd_sc_hd__o22a_4
X_14265_ _14263_/A _14262_/X _14264_/Y VGND VGND VPWR VPWR _14266_/B sky130_fd_sc_hd__a21o_4
XFILLER_167_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12316__A _13045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16004_ _15956_/A _23118_/Q VGND VGND VPWR VPWR _16006_/B sky130_fd_sc_hd__or2_4
X_13216_ _13252_/A _13216_/B VGND VGND VPWR VPWR _13216_/X sky130_fd_sc_hd__or2_4
XFILLER_174_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14196_ _14196_/A _23775_/Q VGND VGND VPWR VPWR _14196_/X sky130_fd_sc_hd__or2_4
XANTENNA__20533__A _20533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13147_ _11887_/A VGND VGND VPWR VPWR _13303_/A sky130_fd_sc_hd__buf_2
XFILLER_135_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21640__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14531__A _14519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13078_ _13067_/A VGND VGND VPWR VPWR _13088_/A sky130_fd_sc_hd__buf_2
X_17955_ _17911_/B _17955_/B VGND VGND VPWR VPWR _17955_/Y sky130_fd_sc_hd__nand2_4
XFILLER_97_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22196__A2 _22194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13147__A _11887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16906_ _16825_/Y _16906_/B VGND VGND VPWR VPWR _16911_/C sky130_fd_sc_hd__nor2_4
X_12029_ _11876_/X VGND VGND VPWR VPWR _16561_/A sky130_fd_sc_hd__buf_2
XFILLER_65_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17886_ _17807_/X _18711_/B _17870_/X _17885_/X VGND VGND VPWR VPWR _17886_/X sky130_fd_sc_hd__a211o_4
X_19625_ _19834_/A _19660_/A VGND VGND VPWR VPWR _19848_/B sky130_fd_sc_hd__or2_4
X_16837_ _16527_/A _16836_/X _16384_/X VGND VGND VPWR VPWR _16837_/X sky130_fd_sc_hd__o21a_4
XFILLER_47_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23335__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15362__A _15362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19556_ _19889_/A VGND VGND VPWR VPWR _19556_/X sky130_fd_sc_hd__buf_2
XANTENNA__21083__B _21370_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16768_ _16768_/A _16768_/B _16767_/X VGND VGND VPWR VPWR _16768_/X sky130_fd_sc_hd__or3_4
XFILLER_34_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18507_ _17635_/D _17617_/Y _17613_/Y VGND VGND VPWR VPWR _18507_/X sky130_fd_sc_hd__o21a_4
X_15719_ _12758_/A _15657_/B VGND VGND VPWR VPWR _15719_/X sky130_fd_sc_hd__or2_4
XANTENNA__19769__A HRDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19487_ _24175_/Q _19481_/X HRDATA[27] _19482_/X VGND VGND VPWR VPWR _19487_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16699_ _16588_/A _16699_/B _16699_/C VGND VGND VPWR VPWR _16703_/B sky130_fd_sc_hd__and3_4
XFILLER_55_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18438_ _18376_/A _17448_/B VGND VGND VPWR VPWR _18438_/Y sky130_fd_sc_hd__nor2_4
XFILLER_94_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22656__B1 _12548_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17289__A _14701_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18369_ _18402_/A _18368_/X _17903_/A VGND VGND VPWR VPWR _18370_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__14706__A _14295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20400_ _24431_/Q _20318_/B VGND VGND VPWR VPWR _20400_/Y sky130_fd_sc_hd__nand2_4
X_21380_ _21249_/X _21377_/X _23889_/Q _21374_/X VGND VGND VPWR VPWR _23889_/D sky130_fd_sc_hd__o22a_4
X_20331_ _20331_/A VGND VGND VPWR VPWR _20331_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20682__A2 _20681_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12226__A _13045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23050_ _18101_/X _23055_/B VGND VGND VPWR VPWR _23050_/X sky130_fd_sc_hd__or2_4
X_20262_ _20261_/X VGND VGND VPWR VPWR _20262_/X sky130_fd_sc_hd__buf_2
XANTENNA__19824__A1 _19705_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22001_ _21821_/X _21996_/X _16388_/B _22000_/X VGND VGND VPWR VPWR _22001_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20193_ _20118_/Y _20192_/X VGND VGND VPWR VPWR _20193_/X sky130_fd_sc_hd__and2_4
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13057__A _13103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23952_ _24080_/CLK _23952_/D VGND VGND VPWR VPWR _16412_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24331__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21934__A2 _21930_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22903_ _22884_/A _22902_/X VGND VGND VPWR VPWR HWDATA[31] sky130_fd_sc_hd__nor2_4
XFILLER_84_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23883_ _24074_/CLK _23883_/D VGND VGND VPWR VPWR _12665_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12896__A _12873_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15272__A _14272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22834_ _22814_/X _22834_/B VGND VGND VPWR VPWR HWDATA[12] sky130_fd_sc_hd__nor2_4
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24260__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16087__B _16085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18012__B1 _17014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22895__B1 _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22765_ SYSTICKCLKDIV[5] VGND VGND VPWR VPWR _22765_/Y sky130_fd_sc_hd__inv_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22817__B _18774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19760__B1 _17816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21716_ _21534_/X _21713_/X _23697_/Q _21710_/X VGND VGND VPWR VPWR _23697_/D sky130_fd_sc_hd__o22a_4
XFILLER_25_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22696_ _21532_/A _22694_/X _23122_/Q _22691_/X VGND VGND VPWR VPWR _22696_/X sky130_fd_sc_hd__o22a_4
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24435_ _24428_/CLK _24435_/D HRESETn VGND VGND VPWR VPWR _20318_/A sky130_fd_sc_hd__dfrtp_4
X_21647_ _21587_/X _21641_/X _14488_/B _21645_/X VGND VGND VPWR VPWR _23739_/D sky130_fd_sc_hd__o22a_4
XFILLER_138_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14616__A _14616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12380_ _13530_/A _12353_/X _12379_/X VGND VGND VPWR VPWR _12380_/X sky130_fd_sc_hd__or3_4
X_24366_ _24360_/CLK _24366_/D HRESETn VGND VGND VPWR VPWR _24366_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21578_ _21523_/A VGND VGND VPWR VPWR _21578_/X sky130_fd_sc_hd__buf_2
XFILLER_123_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23317_ _23456_/CLK _23317_/D VGND VGND VPWR VPWR _15003_/B sky130_fd_sc_hd__dfxtp_4
X_20529_ _24234_/Q _20420_/X _20528_/Y VGND VGND VPWR VPWR _20530_/A sky130_fd_sc_hd__o21a_4
XFILLER_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24297_ _24357_/CLK _24297_/D HRESETn VGND VGND VPWR VPWR _19246_/A sky130_fd_sc_hd__dfrtp_4
X_14050_ _11674_/A _14050_/B _14050_/C VGND VGND VPWR VPWR _14084_/B sky130_fd_sc_hd__or3_4
X_23248_ _24080_/CLK _22499_/X VGND VGND VPWR VPWR _16438_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_107_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13001_ _12881_/A _12997_/X _13001_/C VGND VGND VPWR VPWR _13001_/X sky130_fd_sc_hd__or3_4
XFILLER_97_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15447__A _15447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23179_ _24012_/CLK _23179_/D VGND VGND VPWR VPWR _12520_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21622__B2 _21617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14351__A _12401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23086__D _23084_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20976__A3 _20974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19579__B1 HRDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18758__A _18744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17740_ _17740_/A VGND VGND VPWR VPWR _17741_/A sky130_fd_sc_hd__buf_2
XFILLER_48_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14952_ _14919_/A _23958_/Q VGND VGND VPWR VPWR _14952_/X sky130_fd_sc_hd__or2_4
XANTENNA__20189__A1 _24466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13863__A1 _11854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21925__A2 _21923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13903_ _14348_/A _13898_/X _13902_/X VGND VGND VPWR VPWR _13903_/X sky130_fd_sc_hd__or3_4
X_17671_ _17671_/A _17671_/B VGND VGND VPWR VPWR _17779_/C sky130_fd_sc_hd__nor2_4
XFILLER_130_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14883_ _14127_/A _23606_/Q VGND VGND VPWR VPWR _14883_/X sky130_fd_sc_hd__or2_4
XFILLER_169_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19410_ _19407_/X _18309_/X _19407_/X _24231_/Q VGND VGND VPWR VPWR _19410_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15182__A _15029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16622_ _16662_/A _23794_/Q VGND VGND VPWR VPWR _16623_/C sky130_fd_sc_hd__or2_4
X_13834_ _12497_/A _23613_/Q VGND VGND VPWR VPWR _13834_/X sky130_fd_sc_hd__or2_4
XFILLER_29_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19341_ _19340_/X _18016_/X _19340_/X _24272_/Q VGND VGND VPWR VPWR _19341_/X sky130_fd_sc_hd__a2bb2o_4
X_13765_ _13753_/A _13765_/B VGND VGND VPWR VPWR _13767_/B sky130_fd_sc_hd__or2_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22886__B1 _17425_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16553_ _16558_/A _23698_/Q VGND VGND VPWR VPWR _16556_/B sky130_fd_sc_hd__or2_4
XFILLER_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15910__A _13564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15504_ _13053_/A _23714_/Q VGND VGND VPWR VPWR _15506_/B sky130_fd_sc_hd__or2_4
X_12716_ _11970_/A _12715_/X VGND VGND VPWR VPWR _12716_/X sky130_fd_sc_hd__and2_4
X_19272_ _19250_/A _19250_/B _19271_/Y VGND VGND VPWR VPWR _19272_/X sky130_fd_sc_hd__o21a_4
XFILLER_71_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16484_ _16164_/X _22326_/A VGND VGND VPWR VPWR _16486_/B sky130_fd_sc_hd__or2_4
X_13696_ _13696_/A VGND VGND VPWR VPWR _13697_/A sky130_fd_sc_hd__buf_2
XFILLER_94_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20528__A _20438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18223_ _18335_/A _17467_/X VGND VGND VPWR VPWR _18225_/C sky130_fd_sc_hd__and2_4
X_12647_ _12632_/A _12647_/B VGND VGND VPWR VPWR _12648_/C sky130_fd_sc_hd__or2_4
X_15435_ _15412_/A _15435_/B _15434_/X VGND VGND VPWR VPWR _15435_/X sky130_fd_sc_hd__or3_4
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14526__A _14519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20247__B _16922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22102__A2 _22099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13430__A _13462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18154_ _18282_/A _18154_/B VGND VGND VPWR VPWR _18155_/D sky130_fd_sc_hd__and2_4
X_15366_ _13699_/A _15307_/B VGND VGND VPWR VPWR _15368_/B sky130_fd_sc_hd__or2_4
X_12578_ _12578_/A VGND VGND VPWR VPWR _12659_/A sky130_fd_sc_hd__buf_2
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22743__A _22736_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14245__B _23807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17105_ _17105_/A VGND VGND VPWR VPWR _17105_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14317_ _14292_/A _14317_/B _14316_/X VGND VGND VPWR VPWR _14317_/X sky130_fd_sc_hd__or3_4
X_11529_ _19053_/A _19054_/A VGND VGND VPWR VPWR _11530_/B sky130_fd_sc_hd__or2_4
XFILLER_129_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15297_ _14574_/A _23480_/Q VGND VGND VPWR VPWR _15299_/B sky130_fd_sc_hd__or2_4
X_18085_ _17812_/X _17862_/X _17812_/X _17854_/Y VGND VGND VPWR VPWR _18085_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21861__B2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12046__A _11941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16741__A _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17036_ _18782_/B _17251_/B VGND VGND VPWR VPWR _17036_/X sky130_fd_sc_hd__and2_4
X_14248_ _14248_/A _23871_/Q VGND VGND VPWR VPWR _14248_/X sky130_fd_sc_hd__or2_4
XANTENNA__21359__A _21338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24133__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11885__A _16116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15357__A _11654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14179_ _15325_/A VGND VGND VPWR VPWR _14229_/A sky130_fd_sc_hd__buf_2
XANTENNA__14261__A _14261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18987_ _18987_/A VGND VGND VPWR VPWR _18987_/X sky130_fd_sc_hd__buf_2
XFILLER_140_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17938_ _17819_/X _17216_/X _17230_/X _17195_/X VGND VGND VPWR VPWR _17938_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24283__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17045__A1 _17037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21094__A _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17869_ _17869_/A VGND VGND VPWR VPWR _17869_/X sky130_fd_sc_hd__buf_2
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18793__A1 _17255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13605__A _12477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19608_ _19571_/X _19577_/X _19606_/X _17398_/A _19607_/X VGND VGND VPWR VPWR _19608_/X
+ sky130_fd_sc_hd__a32o_4
X_20880_ _20880_/A VGND VGND VPWR VPWR _20880_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21822__A _21809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19539_ _19539_/A VGND VGND VPWR VPWR _19687_/C sky130_fd_sc_hd__buf_2
XFILLER_81_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16916__A _17060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15820__A _12848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22550_ _22423_/X _22544_/X _16256_/B _22548_/X VGND VGND VPWR VPWR _23215_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18834__C _18834_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24380__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20438__A _20438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21501_ _21283_/X _21499_/X _15841_/B _21496_/X VGND VGND VPWR VPWR _23811_/D sky130_fd_sc_hd__o22a_4
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22481_ _22480_/X _22474_/X _15122_/B _22421_/A VGND VGND VPWR VPWR _23255_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14436__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24220_ _24182_/CLK _24220_/D HRESETn VGND VGND VPWR VPWR _24220_/Q sky130_fd_sc_hd__dfrtp_4
X_21432_ _21251_/X _21427_/X _16429_/B _21431_/X VGND VGND VPWR VPWR _23856_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20655__A2 _20643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24151_ _24302_/CLK _20035_/Y HRESETn VGND VGND VPWR VPWR _24151_/Q sky130_fd_sc_hd__dfrtp_4
X_21363_ _21304_/X _21362_/X _14583_/B _21359_/X VGND VGND VPWR VPWR _21363_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21852__B2 _21846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16651__A _16675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23102_ _23229_/CLK _22724_/X VGND VGND VPWR VPWR _13765_/B sky130_fd_sc_hd__dfxtp_4
X_20314_ _20287_/A VGND VGND VPWR VPWR _20754_/A sky130_fd_sc_hd__buf_2
XANTENNA__21269__A _21269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24082_ _23922_/CLK _21040_/X VGND VGND VPWR VPWR _24082_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21294_ _21292_/X _21293_/X _23935_/Q _21288_/X VGND VGND VPWR VPWR _23935_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11795__A _11836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23033_ _23008_/X _23030_/Y _23033_/C VGND VGND VPWR VPWR _23033_/X sky130_fd_sc_hd__and3_4
XFILLER_118_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20245_ _20864_/A HRDATA[15] VGND VGND VPWR VPWR _20247_/C sky130_fd_sc_hd__or2_4
XANTENNA__22801__B1 _16918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19962__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14171__A _14171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20176_ _20159_/Y _20160_/Y _11562_/X _20175_/X VGND VGND VPWR VPWR _20176_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12403__B _23724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21368__B1 _23893_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21907__A2 _21902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23935_ _23582_/CLK _23935_/D VGND VGND VPWR VPWR _23935_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13515__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11880_ _11880_/A VGND VGND VPWR VPWR _11881_/A sky130_fd_sc_hd__buf_2
X_23866_ _23391_/CLK _21413_/X VGND VGND VPWR VPWR _14688_/B sky130_fd_sc_hd__dfxtp_4
X_22817_ _18738_/X _18774_/X VGND VGND VPWR VPWR _22817_/X sky130_fd_sc_hd__or2_4
XFILLER_72_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23797_ _23392_/CLK _21519_/X VGND VGND VPWR VPWR _15038_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18536__A1 _18111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13550_ _13534_/A _13476_/B VGND VGND VPWR VPWR _13552_/B sky130_fd_sc_hd__or2_4
XANTENNA__15730__A _12783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22748_ _19920_/X _22736_/X _23086_/B _22743_/Y VGND VGND VPWR VPWR _24126_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12501_ _12501_/A VGND VGND VPWR VPWR _12502_/A sky130_fd_sc_hd__buf_2
X_13481_ _12515_/A _13481_/B _13480_/X VGND VGND VPWR VPWR _13482_/C sky130_fd_sc_hd__and3_4
X_22679_ _22672_/A VGND VGND VPWR VPWR _22679_/X sky130_fd_sc_hd__buf_2
XFILLER_139_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14346__A _14512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13250__A _12338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15220_ _14196_/A _15156_/B VGND VGND VPWR VPWR _15220_/X sky130_fd_sc_hd__or2_4
XFILLER_139_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12432_ _14108_/A VGND VGND VPWR VPWR _12433_/A sky130_fd_sc_hd__buf_2
X_24418_ _23475_/CLK _24418_/D HRESETn VGND VGND VPWR VPWR _24418_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22096__B2 _22094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24156__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15151_ _13954_/A _15151_/B _15150_/X VGND VGND VPWR VPWR _15151_/X sky130_fd_sc_hd__and3_4
X_12363_ _12923_/A VGND VGND VPWR VPWR _12363_/X sky130_fd_sc_hd__buf_2
X_24349_ _24382_/CLK _24349_/D HRESETn VGND VGND VPWR VPWR _11523_/A sky130_fd_sc_hd__dfstp_4
XFILLER_154_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16561__A _16561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14102_ _14138_/A _23775_/Q VGND VGND VPWR VPWR _14103_/C sky130_fd_sc_hd__or2_4
XFILLER_10_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15082_ _15106_/A _15082_/B _15082_/C VGND VGND VPWR VPWR _15083_/C sky130_fd_sc_hd__or3_4
X_12294_ _12294_/A VGND VGND VPWR VPWR _12304_/A sky130_fd_sc_hd__buf_2
XFILLER_49_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22399__A2 _22397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18910_ _16240_/X _18906_/X _24397_/Q _18907_/X VGND VGND VPWR VPWR _24397_/D sky130_fd_sc_hd__o22a_4
X_14033_ _11753_/A _14027_/X _14032_/X VGND VGND VPWR VPWR _14034_/C sky130_fd_sc_hd__or3_4
XANTENNA__15177__A _15017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19890_ _19890_/A _19890_/B VGND VGND VPWR VPWR _19890_/X sky130_fd_sc_hd__and2_4
XANTENNA__14081__A _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21071__A2 _21066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18841_ _18838_/X VGND VGND VPWR VPWR _18842_/A sky130_fd_sc_hd__inv_2
XFILLER_171_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12313__B _23724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18772_ _18772_/A _18762_/Y _18411_/A _18771_/X VGND VGND VPWR VPWR _18772_/X sky130_fd_sc_hd__or4_4
XFILLER_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15984_ _15957_/A _16057_/B VGND VGND VPWR VPWR _15986_/B sky130_fd_sc_hd__or2_4
XFILLER_0_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17723_ _17723_/A VGND VGND VPWR VPWR _17723_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22020__B2 _22014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14935_ _14916_/X _14933_/X _14934_/X VGND VGND VPWR VPWR _14935_/X sky130_fd_sc_hd__and3_4
XANTENNA__13425__A _13468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18775__B2 _16943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19972__B1 _17919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17654_ _16945_/A _17052_/Y _16945_/A _17052_/Y VGND VGND VPWR VPWR _17654_/X sky130_fd_sc_hd__a2bb2o_4
X_14866_ _12425_/A _14864_/X _14866_/C VGND VGND VPWR VPWR _14866_/X sky130_fd_sc_hd__and3_4
XFILLER_1_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16605_ _11694_/X VGND VGND VPWR VPWR _16606_/A sky130_fd_sc_hd__buf_2
X_13817_ _15404_/A _13814_/X _13817_/C VGND VGND VPWR VPWR _13821_/B sky130_fd_sc_hd__and3_4
XFILLER_91_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17585_ _16240_/X _18114_/B VGND VGND VPWR VPWR _17585_/Y sky130_fd_sc_hd__nand2_4
X_14797_ _14667_/A _14795_/X _14797_/C VGND VGND VPWR VPWR _14797_/X sky130_fd_sc_hd__and3_4
XFILLER_56_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19324_ _19324_/A VGND VGND VPWR VPWR _19428_/A sky130_fd_sc_hd__buf_2
XANTENNA__15640__A _14335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16536_ _12106_/A _23538_/Q VGND VGND VPWR VPWR _16536_/X sky130_fd_sc_hd__or2_4
X_13748_ _12616_/A _13740_/X _13748_/C VGND VGND VPWR VPWR _13749_/C sky130_fd_sc_hd__and3_4
XFILLER_32_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20258__A _20257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19255_ _24306_/Q _19255_/B VGND VGND VPWR VPWR _19256_/B sky130_fd_sc_hd__and2_4
X_16467_ _16490_/A _16397_/B VGND VGND VPWR VPWR _16467_/X sky130_fd_sc_hd__or2_4
X_13679_ _13676_/A _13776_/B VGND VGND VPWR VPWR _13680_/C sky130_fd_sc_hd__or2_4
XANTENNA__14256__A _15595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18206_ _17249_/X VGND VGND VPWR VPWR _18206_/X sky130_fd_sc_hd__buf_2
X_15418_ _11878_/A _15416_/X _15418_/C VGND VGND VPWR VPWR _15419_/C sky130_fd_sc_hd__and3_4
X_19186_ _19149_/A _19149_/B _19185_/Y VGND VGND VPWR VPWR _24328_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_5_23_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22087__B2 _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16398_ _16009_/X _16398_/B VGND VGND VPWR VPWR _16399_/C sky130_fd_sc_hd__or2_4
XANTENNA__22473__A _22158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18137_ _17594_/X _17640_/X _18095_/A _17545_/X VGND VGND VPWR VPWR _18137_/X sky130_fd_sc_hd__o22a_4
X_15349_ _15319_/A _23960_/Q VGND VGND VPWR VPWR _15349_/X sky130_fd_sc_hd__or2_4
XANTENNA__16471__A _11684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17502__A2 _17020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21089__A _21118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18068_ _17900_/A VGND VGND VPWR VPWR _18068_/X sky130_fd_sc_hd__buf_2
XFILLER_171_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17019_ _17018_/X VGND VGND VPWR VPWR _17019_/X sky130_fd_sc_hd__buf_2
XANTENNA__15087__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12504__A _12504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21062__A2 _21059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20030_ _20029_/X VGND VGND VPWR VPWR _20030_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20721__A HRDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22011__A1 _21838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22011__B2 _22007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21981_ _21941_/A VGND VGND VPWR VPWR _21981_/X sky130_fd_sc_hd__buf_2
XFILLER_6_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23720_ _23337_/CLK _21679_/X VGND VGND VPWR VPWR _23720_/Q sky130_fd_sc_hd__dfxtp_4
X_20932_ _20931_/X VGND VGND VPWR VPWR _20932_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22648__A _22648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23651_ _23939_/CLK _21786_/X VGND VGND VPWR VPWR _15837_/B sky130_fd_sc_hd__dfxtp_4
X_20863_ _20863_/A VGND VGND VPWR VPWR _20943_/A sky130_fd_sc_hd__buf_2
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16646__A _16646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22314__A2 _22308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22602_ _22425_/X _22601_/X _16041_/B _22598_/X VGND VGND VPWR VPWR _23182_/D sky130_fd_sc_hd__o22a_4
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15550__A _14450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23582_ _23582_/CLK _23582_/D VGND VGND VPWR VPWR _13733_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20794_ _18548_/X _20675_/X _20780_/X _20793_/Y VGND VGND VPWR VPWR _20794_/X sky130_fd_sc_hd__a211o_4
XANTENNA__20168__A IRQ[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24179__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22533_ _22480_/X _22529_/X _15172_/B _22498_/A VGND VGND VPWR VPWR _22533_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14166__A _14131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22464_ _20818_/A VGND VGND VPWR VPWR _22464_/X sky130_fd_sc_hd__buf_2
XANTENNA__22383__A _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24203_ _23671_/CLK _19720_/X HRESETn VGND VGND VPWR VPWR _11965_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20628__A2 _20616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21415_ _21309_/X _21412_/X _23864_/Q _21409_/X VGND VGND VPWR VPWR _23864_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21825__B2 _21822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17477__A _17145_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22395_ _22153_/X _22390_/X _14355_/B _22394_/X VGND VGND VPWR VPWR _22395_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16381__A _16380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24134_ _24134_/CLK _24134_/D HRESETn VGND VGND VPWR VPWR _16970_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_162_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21346_ _21275_/X _21341_/X _13309_/B _21345_/X VGND VGND VPWR VPWR _23910_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12318__A1 _12882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24065_ _23908_/CLK _24065_/D VGND VGND VPWR VPWR _24065_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_162_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21277_ _21275_/X _21269_/X _13364_/B _21276_/X VGND VGND VPWR VPWR _23942_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12414__A _13542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23016_ _23008_/X _23016_/B _23015_/X VGND VGND VPWR VPWR _23016_/X sky130_fd_sc_hd__and3_4
XANTENNA__21053__A2 _21052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_43_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR _23438_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21727__A _21727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20228_ _20216_/D _17033_/A VGND VGND VPWR VPWR _20229_/A sky130_fd_sc_hd__or2_4
XANTENNA__22250__B2 _22248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15725__A _13091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20159_ _20159_/A VGND VGND VPWR VPWR _20159_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22002__B2 _22000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12981_ _12980_/X VGND VGND VPWR VPWR _12983_/B sky130_fd_sc_hd__inv_2
XFILLER_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18757__A1 _17980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22553__A2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19954__B1 _23086_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14720_ _13666_/A _14720_/B VGND VGND VPWR VPWR _14722_/B sky130_fd_sc_hd__or2_4
X_23918_ _23918_/CLK _23918_/D VGND VGND VPWR VPWR _16054_/B sky130_fd_sc_hd__dfxtp_4
X_11932_ _11932_/A VGND VGND VPWR VPWR _11933_/A sky130_fd_sc_hd__buf_2
XFILLER_131_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22558__A _22558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21462__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11863_ _13046_/A VGND VGND VPWR VPWR _11864_/A sky130_fd_sc_hd__buf_2
X_14651_ _14647_/X _14649_/X _14650_/X VGND VGND VPWR VPWR _14651_/X sky130_fd_sc_hd__and3_4
X_23849_ _24073_/CLK _21442_/X VGND VGND VPWR VPWR _23849_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15460__A _12587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13602_ _14448_/A _13597_/X _13601_/X VGND VGND VPWR VPWR _13602_/X sky130_fd_sc_hd__and3_4
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _17170_/Y _17372_/A VGND VGND VPWR VPWR _17371_/A sky130_fd_sc_hd__or2_4
XPHY_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _11772_/X VGND VGND VPWR VPWR _11836_/A sky130_fd_sc_hd__buf_2
X_14582_ _13689_/A _14559_/X _14566_/X _14573_/X _14581_/X VGND VGND VPWR VPWR _14582_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16321_ _16192_/A _16256_/B VGND VGND VPWR VPWR _16323_/B sky130_fd_sc_hd__or2_4
X_13533_ _12402_/X _13533_/B _13532_/X VGND VGND VPWR VPWR _13533_/X sky130_fd_sc_hd__and3_4
XFILLER_13_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14076__A _12581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19040_ _24357_/Q VGND VGND VPWR VPWR _19040_/Y sky130_fd_sc_hd__inv_2
X_13464_ _13474_/A _13464_/B _13463_/X VGND VGND VPWR VPWR _13464_/X sky130_fd_sc_hd__and3_4
X_16252_ _16099_/X VGND VGND VPWR VPWR _16287_/A sky130_fd_sc_hd__buf_2
XANTENNA__22069__B2 _22064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12415_ _15887_/A _12409_/X _12415_/C VGND VGND VPWR VPWR _12416_/C sky130_fd_sc_hd__or3_4
X_15203_ _14235_/A _15146_/B VGND VGND VPWR VPWR _15205_/B sky130_fd_sc_hd__or2_4
X_16183_ _13379_/A VGND VGND VPWR VPWR _16231_/A sky130_fd_sc_hd__buf_2
X_13395_ _13376_/A _13393_/X _13395_/C VGND VGND VPWR VPWR _13399_/B sky130_fd_sc_hd__and3_4
XFILLER_138_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21816__B2 _21810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12346_ _11739_/A _12346_/B _12346_/C VGND VGND VPWR VPWR _12352_/B sky130_fd_sc_hd__and3_4
X_15134_ _15267_/A _15134_/B VGND VGND VPWR VPWR _15137_/B sky130_fd_sc_hd__or2_4
XFILLER_154_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14523__B _14523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19942_ _19938_/X _24167_/Q _19939_/X _20561_/B VGND VGND VPWR VPWR _24167_/D sky130_fd_sc_hd__o22a_4
X_15065_ _15091_/A _15065_/B _15064_/X VGND VGND VPWR VPWR _15065_/X sky130_fd_sc_hd__or3_4
X_12277_ _12273_/A _12390_/B VGND VGND VPWR VPWR _12277_/X sky130_fd_sc_hd__or2_4
XFILLER_114_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12324__A _13230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14016_ _11750_/A VGND VGND VPWR VPWR _15369_/A sky130_fd_sc_hd__buf_2
XFILLER_49_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21044__A2 _21038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19873_ _19752_/B _19752_/D VGND VGND VPWR VPWR _19873_/X sky130_fd_sc_hd__or2_4
XFILLER_110_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18824_ _18786_/A VGND VGND VPWR VPWR _18824_/X sky130_fd_sc_hd__buf_2
XFILLER_49_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_0_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18755_ _17100_/A _18754_/Y _18383_/Y VGND VGND VPWR VPWR _18755_/X sky130_fd_sc_hd__o21a_4
X_15967_ _15967_/A _16048_/B VGND VGND VPWR VPWR _15967_/X sky130_fd_sc_hd__or2_4
XANTENNA__14482__A1 _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14482__B2 _14481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13155__A _13183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19945__B1 _22745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17706_ _17705_/X VGND VGND VPWR VPWR _17706_/Y sky130_fd_sc_hd__inv_2
X_14918_ _14922_/A _14852_/B VGND VGND VPWR VPWR _14918_/X sky130_fd_sc_hd__or2_4
X_18686_ _18670_/X _11639_/A _18685_/Y _24473_/Q _18625_/X VGND VGND VPWR VPWR _18686_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_48_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15898_ _13521_/X _15896_/X _15897_/X VGND VGND VPWR VPWR _15898_/X sky130_fd_sc_hd__and3_4
XANTENNA__21752__B1 _15139_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22468__A _20859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21372__A _21405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17637_ _17384_/X _17637_/B _17637_/C _17637_/D VGND VGND VPWR VPWR _17638_/A sky130_fd_sc_hd__or4_4
XANTENNA__24321__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14849_ _12188_/A _14912_/B VGND VGND VPWR VPWR _14849_/X sky130_fd_sc_hd__or2_4
XANTENNA__12994__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16466__A _13367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15370__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17568_ _16016_/Y _17024_/A _17024_/A _17567_/X VGND VGND VPWR VPWR _18076_/B sky130_fd_sc_hd__a2bb2o_4
X_19307_ _19233_/B VGND VGND VPWR VPWR _19307_/Y sky130_fd_sc_hd__inv_2
X_16519_ _11684_/X _16519_/B _16519_/C VGND VGND VPWR VPWR _16519_/X sky130_fd_sc_hd__and3_4
X_17499_ _18290_/A VGND VGND VPWR VPWR _17499_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17184__B1 _17339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19238_ _24289_/Q _19237_/X VGND VGND VPWR VPWR _19295_/A sky130_fd_sc_hd__and2_4
XANTENNA__24471__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20716__A _20857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19169_ _19158_/B VGND VGND VPWR VPWR _19169_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14714__A _14296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21200_ _20464_/X _21198_/X _23981_/Q _21195_/X VGND VGND VPWR VPWR _21200_/X sky130_fd_sc_hd__o22a_4
XFILLER_173_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22180_ _22194_/A VGND VGND VPWR VPWR _22180_/X sky130_fd_sc_hd__buf_2
XANTENNA__18684__B1 _18019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22931__A _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21131_ _21024_/X _21104_/A _24021_/Q _21086_/X VGND VGND VPWR VPWR _21131_/X sky130_fd_sc_hd__o22a_4
XFILLER_99_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21062_ _20719_/X _21059_/X _15490_/B _21056_/X VGND VGND VPWR VPWR _24066_/D sky130_fd_sc_hd__o22a_4
XFILLER_87_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22232__B2 _22227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20013_ _18143_/X _20007_/X _20012_/Y _19994_/X VGND VGND VPWR VPWR _20013_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15545__A _13687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20794__A1 _18548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22535__A2 _22508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21964_ _21957_/A VGND VGND VPWR VPWR _21964_/X sky130_fd_sc_hd__buf_2
XFILLER_39_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23703_ _23770_/CLK _21702_/X VGND VGND VPWR VPWR _15179_/B sky130_fd_sc_hd__dfxtp_4
X_20915_ _21304_/A VGND VGND VPWR VPWR _20915_/X sky130_fd_sc_hd__buf_2
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21895_ _21909_/A VGND VGND VPWR VPWR _21895_/X sky130_fd_sc_hd__buf_2
XFILLER_27_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23569__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15280__A _15022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23634_ _23922_/CLK _21818_/X VGND VGND VPWR VPWR _23634_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22299__B2 _22298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _20244_/X _20845_/X _20639_/X VGND VGND VPWR VPWR _20846_/Y sky130_fd_sc_hd__o21ai_4
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23565_ _23501_/CLK _21955_/X VGND VGND VPWR VPWR _16203_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20777_ _20664_/A _20777_/B _20777_/C VGND VGND VPWR VPWR _20777_/X sky130_fd_sc_hd__and3_4
XFILLER_11_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17714__A2 _17389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18911__A1 _12419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22516_ _22449_/X _22515_/X _15704_/B _22512_/X VGND VGND VPWR VPWR _22516_/X sky130_fd_sc_hd__o22a_4
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23496_ _23496_/CLK _23496_/D VGND VGND VPWR VPWR _23496_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23002__A _22910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22447_ _20632_/A VGND VGND VPWR VPWR _22447_/X sky130_fd_sc_hd__buf_2
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12200_ _12569_/A _23532_/Q VGND VGND VPWR VPWR _12201_/C sky130_fd_sc_hd__or2_4
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13180_ _11902_/A _23655_/Q VGND VGND VPWR VPWR _13181_/C sky130_fd_sc_hd__or2_4
XANTENNA__21274__A2 _21269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22378_ _22125_/X _22376_/X _12999_/B _22373_/X VGND VGND VPWR VPWR _22378_/X sky130_fd_sc_hd__o22a_4
XFILLER_135_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15439__B _15511_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12131_ _11686_/X _12123_/X _12131_/C VGND VGND VPWR VPWR _12147_/B sky130_fd_sc_hd__and3_4
X_24117_ _23544_/CLK _24117_/D HRESETn VGND VGND VPWR VPWR _18948_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_163_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21329_ _21247_/X _21327_/X _23922_/Q _21324_/X VGND VGND VPWR VPWR _23922_/D sky130_fd_sc_hd__o22a_4
XFILLER_2_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24048_ _23662_/CLK _21095_/X VGND VGND VPWR VPWR _16397_/B sky130_fd_sc_hd__dfxtp_4
X_12062_ _11963_/A VGND VGND VPWR VPWR _16732_/A sky130_fd_sc_hd__buf_2
XFILLER_104_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20234__B1 _20233_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16870_ _16869_/X VGND VGND VPWR VPWR _16873_/C sky130_fd_sc_hd__inv_2
XFILLER_49_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15821_ _12886_/A _15819_/X _15820_/X VGND VGND VPWR VPWR _15821_/X sky130_fd_sc_hd__and3_4
XFILLER_65_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24344__CLK _24342_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18540_ _17435_/Y _18539_/X VGND VGND VPWR VPWR _18540_/Y sky130_fd_sc_hd__nand2_4
X_15752_ _12758_/A _23908_/Q VGND VGND VPWR VPWR _15754_/B sky130_fd_sc_hd__or2_4
X_12964_ _12940_/A _12964_/B VGND VGND VPWR VPWR _12965_/C sky130_fd_sc_hd__or2_4
XFILLER_92_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14703_ _14703_/A VGND VGND VPWR VPWR _14705_/A sky130_fd_sc_hd__inv_2
X_11915_ _11915_/A VGND VGND VPWR VPWR _12870_/A sky130_fd_sc_hd__buf_2
X_18471_ _17396_/B _18469_/X _18176_/A VGND VGND VPWR VPWR _18471_/Y sky130_fd_sc_hd__a21oi_4
X_15683_ _12745_/A _15681_/X _15682_/X VGND VGND VPWR VPWR _15683_/X sky130_fd_sc_hd__and3_4
X_12895_ _12895_/A _23433_/Q VGND VGND VPWR VPWR _12895_/X sky130_fd_sc_hd__or2_4
X_17422_ _17421_/X VGND VGND VPWR VPWR _17423_/B sky130_fd_sc_hd__inv_2
XANTENNA__24494__CLK _24306_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14634_ _14667_/A _14632_/X _14633_/X VGND VGND VPWR VPWR _14641_/B sky130_fd_sc_hd__and3_4
X_11846_ _11836_/A _23668_/Q VGND VGND VPWR VPWR _11846_/X sky130_fd_sc_hd__or2_4
XPHY_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _15582_/X VGND VGND VPWR VPWR _17353_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21920__A _21906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11777_ _11686_/X _11749_/X _11776_/X VGND VGND VPWR VPWR _11777_/X sky130_fd_sc_hd__and3_4
X_14565_ _15394_/A _14565_/B _14564_/X VGND VGND VPWR VPWR _14565_/X sky130_fd_sc_hd__and3_4
XPHY_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18902__A1 _12180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16304_ _11903_/X _16304_/B VGND VGND VPWR VPWR _16305_/C sky130_fd_sc_hd__or2_4
X_13516_ _13515_/X _13449_/B VGND VGND VPWR VPWR _13516_/X sky130_fd_sc_hd__or2_4
XANTENNA__15716__A1 _13307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17284_ _14613_/X VGND VGND VPWR VPWR _17284_/Y sky130_fd_sc_hd__inv_2
X_14496_ _14509_/A _14494_/X _14495_/X VGND VGND VPWR VPWR _14497_/C sky130_fd_sc_hd__and3_4
XANTENNA__16913__B1 _16905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_HCLK_A clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19023_ _19010_/X _19022_/X _19010_/X _11535_/A VGND VGND VPWR VPWR _24361_/D sky130_fd_sc_hd__a2bb2o_4
X_16235_ _16185_/A _16233_/X _16234_/X VGND VGND VPWR VPWR _16236_/C sky130_fd_sc_hd__and3_4
X_13447_ _12885_/A _13447_/B VGND VGND VPWR VPWR _13447_/X sky130_fd_sc_hd__or2_4
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14534__A _14510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21265__A2 _21257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13378_ _13378_/A _13296_/B VGND VGND VPWR VPWR _13378_/X sky130_fd_sc_hd__or2_4
X_16166_ _13397_/A VGND VGND VPWR VPWR _16166_/X sky130_fd_sc_hd__buf_2
XFILLER_115_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15117_ _14911_/X VGND VGND VPWR VPWR _15117_/Y sky130_fd_sc_hd__inv_2
X_12329_ _12329_/A VGND VGND VPWR VPWR _12625_/A sky130_fd_sc_hd__buf_2
X_16097_ _16112_/A VGND VGND VPWR VPWR _16108_/A sky130_fd_sc_hd__buf_2
XANTENNA__12054__A _16592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18681__A3 _18677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19925_ _22745_/A VGND VGND VPWR VPWR _19925_/X sky130_fd_sc_hd__buf_2
X_15048_ _15047_/Y VGND VGND VPWR VPWR _15048_/X sky130_fd_sc_hd__buf_2
XANTENNA__22214__B2 _22212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20271__A _20270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12989__A _12854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15365__A _13695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19856_ _19823_/B _19848_/B _19849_/B _19725_/A VGND VGND VPWR VPWR _19856_/X sky130_fd_sc_hd__o22a_4
XFILLER_69_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18807_ _13266_/X _18803_/X _24456_/Q _18804_/X VGND VGND VPWR VPWR _24456_/D sky130_fd_sc_hd__o22a_4
XFILLER_96_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19787_ _19787_/A _19787_/B VGND VGND VPWR VPWR _19807_/A sky130_fd_sc_hd__or2_4
X_16999_ _16945_/A _16999_/B VGND VGND VPWR VPWR _16999_/X sky130_fd_sc_hd__or2_4
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17580__A _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18738_ _18409_/A _18730_/Y _18731_/X _18008_/A _18737_/X VGND VGND VPWR VPWR _18738_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_114_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21725__B1 _12500_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22198__A _22176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18669_ _11511_/A VGND VGND VPWR VPWR _18670_/A sky130_fd_sc_hd__buf_2
XFILLER_58_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16196__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14709__A _13596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20700_ _20700_/A _20700_/B _20699_/X VGND VGND VPWR VPWR _20700_/X sky130_fd_sc_hd__and3_4
XANTENNA__13613__A _15018_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21680_ _21558_/X _21677_/X _23719_/Q _21674_/X VGND VGND VPWR VPWR _21680_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22926__A _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14428__B _14423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20631_ _24229_/Q _20534_/X _20630_/X VGND VGND VPWR VPWR _20632_/A sky130_fd_sc_hd__o21a_4
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23861__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12229__A _12727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22150__B1 _13738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23350_ _23095_/CLK _22320_/X VGND VGND VPWR VPWR _14852_/B sky130_fd_sc_hd__dfxtp_4
X_20562_ _20251_/A _20561_/X _20306_/X VGND VGND VPWR VPWR _20562_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_137_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22301_ _22294_/A VGND VGND VPWR VPWR _22301_/X sky130_fd_sc_hd__buf_2
XFILLER_20_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23281_ _23281_/CLK _23281_/D VGND VGND VPWR VPWR _16751_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_165_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20493_ _20493_/A VGND VGND VPWR VPWR _20494_/B sky130_fd_sc_hd__buf_2
XANTENNA__14444__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24217__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22232_ _22101_/X _22230_/X _16664_/B _22227_/X VGND VGND VPWR VPWR _22232_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18657__B1 _18009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22453__B2 _22445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22163_ _20958_/A VGND VGND VPWR VPWR _22163_/X sky130_fd_sc_hd__buf_2
XFILLER_132_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21114_ _20719_/X _21111_/X _15465_/B _21108_/X VGND VGND VPWR VPWR _21114_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23241__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22094_ _22106_/A VGND VGND VPWR VPWR _22094_/X sky130_fd_sc_hd__buf_2
XANTENNA__12899__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21045_ _21045_/A VGND VGND VPWR VPWR _21045_/X sky130_fd_sc_hd__buf_2
XANTENNA__15275__A _14131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_HCLK_A clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22996_ _18394_/X _22973_/B VGND VGND VPWR VPWR _22997_/C sky130_fd_sc_hd__or2_4
XFILLER_83_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21947_ _21813_/X _21946_/X _23571_/Q _21943_/X VGND VGND VPWR VPWR _21947_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21192__B2 _21188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11700_ _13223_/A VGND VGND VPWR VPWR _11701_/A sky130_fd_sc_hd__buf_2
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12679_/Y VGND VGND VPWR VPWR _12680_/X sky130_fd_sc_hd__buf_2
XFILLER_42_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21878_ _21877_/X _21875_/X _14739_/B _21870_/X VGND VGND VPWR VPWR _23609_/D sky130_fd_sc_hd__o22a_4
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A VGND VGND VPWR VPWR _11631_/X sky130_fd_sc_hd__buf_2
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _20828_/X VGND VGND VPWR VPWR _20829_/Y sky130_fd_sc_hd__inv_2
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23617_ _23617_/CLK _21859_/X VGND VGND VPWR VPWR _15555_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21495__A2 _21492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _24451_/Q IRQ[14] VGND VGND VPWR VPWR _11562_/X sky130_fd_sc_hd__and2_4
X_14350_ _14517_/A _23772_/Q VGND VGND VPWR VPWR _14350_/X sky130_fd_sc_hd__or2_4
XFILLER_156_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23548_ _23323_/CLK _21979_/X VGND VGND VPWR VPWR _23548_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22692__B2 _22691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13301_ _13301_/A _13365_/B VGND VGND VPWR VPWR _13301_/X sky130_fd_sc_hd__or2_4
XFILLER_128_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14281_ _14311_/A _24028_/Q VGND VGND VPWR VPWR _14283_/B sky130_fd_sc_hd__or2_4
X_23479_ _23864_/CLK _22085_/X VGND VGND VPWR VPWR _15169_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16020_ _16056_/A VGND VGND VPWR VPWR _16066_/A sky130_fd_sc_hd__buf_2
X_13232_ _13232_/A _13230_/X _13231_/X VGND VGND VPWR VPWR _13232_/X sky130_fd_sc_hd__and3_4
XFILLER_40_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18648__B1 _17805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13163_ _13276_/A _13161_/X _13162_/X VGND VGND VPWR VPWR _13163_/X sky130_fd_sc_hd__and3_4
XFILLER_83_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24357__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12114_ _16608_/A _12114_/B VGND VGND VPWR VPWR _12114_/X sky130_fd_sc_hd__or2_4
XANTENNA__21187__A _21202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13094_ _13094_/A _13018_/B VGND VGND VPWR VPWR _13096_/B sky130_fd_sc_hd__or2_4
X_17971_ _17801_/X _17971_/B VGND VGND VPWR VPWR _17972_/D sky130_fd_sc_hd__and2_4
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19710_ _19494_/A _19848_/A _19677_/A VGND VGND VPWR VPWR _19711_/A sky130_fd_sc_hd__o21a_4
X_16922_ _16915_/C _16915_/A _16922_/C _16914_/A VGND VGND VPWR VPWR _16922_/X sky130_fd_sc_hd__or4_4
XFILLER_46_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12045_ _16704_/A _12124_/B VGND VGND VPWR VPWR _12045_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_13_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_13_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19641_ _19446_/A _19640_/X HRDATA[2] _19461_/X VGND VGND VPWR VPWR _19642_/A sky130_fd_sc_hd__o22a_4
X_16853_ _15933_/X _16246_/B _15933_/X _16246_/B VGND VGND VPWR VPWR _16853_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15804_ _12885_/A _15804_/B VGND VGND VPWR VPWR _15805_/C sky130_fd_sc_hd__or2_4
XFILLER_133_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19572_ HRDATA[28] VGND VGND VPWR VPWR _20364_/B sky130_fd_sc_hd__buf_2
XFILLER_65_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15913__A _15912_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16784_ _16759_/A _16782_/X _16783_/X VGND VGND VPWR VPWR _16784_/X sky130_fd_sc_hd__and3_4
X_13996_ _13663_/A _13996_/B _13996_/C VGND VGND VPWR VPWR _13996_/X sky130_fd_sc_hd__or3_4
XFILLER_19_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18523_ _17421_/X _18520_/X _17890_/X _18522_/X VGND VGND VPWR VPWR _18523_/X sky130_fd_sc_hd__a211o_4
X_15735_ _12783_/X _15735_/B VGND VGND VPWR VPWR _15736_/C sky130_fd_sc_hd__or2_4
X_12947_ _12641_/A _12947_/B _12947_/C VGND VGND VPWR VPWR _12979_/B sky130_fd_sc_hd__or3_4
XFILLER_46_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13433__A _13330_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18454_ _18367_/A _18366_/X VGND VGND VPWR VPWR _18454_/Y sky130_fd_sc_hd__nand2_4
X_15666_ _12722_/A _15664_/X _15665_/X VGND VGND VPWR VPWR _15666_/X sky130_fd_sc_hd__and3_4
X_12878_ _12878_/A _12935_/B VGND VGND VPWR VPWR _12880_/B sky130_fd_sc_hd__or2_4
XANTENNA__19128__A1 _18948_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17405_ _17404_/X VGND VGND VPWR VPWR _17436_/A sky130_fd_sc_hd__buf_2
X_14617_ _14235_/A VGND VGND VPWR VPWR _14819_/A sky130_fd_sc_hd__buf_2
XFILLER_159_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18385_ _18200_/X _18381_/X _18382_/X _18383_/Y _18384_/Y VGND VGND VPWR VPWR _18386_/A
+ sky130_fd_sc_hd__a32o_4
X_11829_ _12168_/A _11827_/X _11828_/X VGND VGND VPWR VPWR _11829_/X sky130_fd_sc_hd__and3_4
X_15597_ _15611_/A _15533_/B VGND VGND VPWR VPWR _15597_/X sky130_fd_sc_hd__or2_4
XANTENNA__12049__A _16595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17336_ _12570_/A _17297_/X _21081_/A _17039_/A VGND VGND VPWR VPWR _17336_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21486__A2 _21485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14548_ _14547_/X VGND VGND VPWR VPWR _14548_/X sky130_fd_sc_hd__buf_2
XANTENNA__22683__B2 _22648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17267_ _17266_/X _17913_/B VGND VGND VPWR VPWR _17915_/B sky130_fd_sc_hd__and2_4
XFILLER_147_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14479_ _14292_/A _14475_/X _14478_/X VGND VGND VPWR VPWR _14479_/X sky130_fd_sc_hd__or3_4
X_19006_ _19004_/Y _19005_/Y _11538_/B VGND VGND VPWR VPWR _19006_/X sky130_fd_sc_hd__o21a_4
X_16218_ _16202_/A _16142_/B VGND VGND VPWR VPWR _16218_/X sky130_fd_sc_hd__or2_4
XFILLER_134_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19774__B HRDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17198_ _17198_/A VGND VGND VPWR VPWR _17198_/X sky130_fd_sc_hd__buf_2
XANTENNA__23264__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16149_ _16142_/A _16149_/B VGND VGND VPWR VPWR _16151_/B sky130_fd_sc_hd__or2_4
XANTENNA__17575__A _11608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20997__A1 _22846_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21097__A _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19908_ _19908_/A VGND VGND VPWR VPWR _20871_/A sky130_fd_sc_hd__buf_2
XANTENNA__13608__A _13823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12512__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21410__A2 _21405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19839_ _19839_/A _19815_/B _19849_/B VGND VGND VPWR VPWR _19839_/X sky130_fd_sc_hd__and3_4
XANTENNA__12231__B _24012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15823__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22850_ _15048_/X _22848_/X _22849_/X VGND VGND VPWR VPWR _22850_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21801_ _21594_/X _21798_/X _23640_/Q _21795_/X VGND VGND VPWR VPWR _23640_/D sky130_fd_sc_hd__o22a_4
X_22781_ _22781_/A _22781_/B VGND VGND VPWR VPWR _22781_/Y sky130_fd_sc_hd__nand2_4
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21174__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14439__A _12537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13343__A _13343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21732_ _21560_/X _21727_/X _23686_/Q _21731_/X VGND VGND VPWR VPWR _23686_/D sky130_fd_sc_hd__o22a_4
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21663_ _21677_/A VGND VGND VPWR VPWR _21663_/X sky130_fd_sc_hd__buf_2
XFILLER_12_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24451_ _23475_/CLK _18814_/X HRESETn VGND VGND VPWR VPWR _24451_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20614_ _20510_/A VGND VGND VPWR VPWR _20614_/X sky130_fd_sc_hd__buf_2
X_23402_ _23404_/CLK _23402_/D VGND VGND VPWR VPWR _12819_/B sky130_fd_sc_hd__dfxtp_4
X_24382_ _24382_/CLK _24382_/D HRESETn VGND VGND VPWR VPWR _24382_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22674__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21594_ _20959_/A VGND VGND VPWR VPWR _21594_/X sky130_fd_sc_hd__buf_2
XANTENNA__23607__CLK _23864_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23333_ _23557_/CLK _23333_/D VGND VGND VPWR VPWR _22337_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__11798__A _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19965__A _17801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20545_ _20545_/A VGND VGND VPWR VPWR _20545_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21229__A2 _21226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23264_ _23203_/CLK _23264_/D VGND VGND VPWR VPWR _23264_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20476_ _20344_/X _20474_/X _11538_/A _20475_/X VGND VGND VPWR VPWR _20476_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12914__A1 _11857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22215_ _22208_/A VGND VGND VPWR VPWR _22215_/X sky130_fd_sc_hd__buf_2
XFILLER_105_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12914__B2 _12913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17485__A _12680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23195_ _24096_/CLK _22578_/X VGND VGND VPWR VPWR _14491_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22146_ _22461_/A VGND VGND VPWR VPWR _22146_/X sky130_fd_sc_hd__buf_2
XFILLER_160_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22077_ _21867_/X _22074_/X _13845_/B _22071_/X VGND VGND VPWR VPWR _22077_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17066__C1 _17017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21028_ _21028_/A VGND VGND VPWR VPWR _21134_/B sky130_fd_sc_hd__buf_2
XANTENNA__21401__A2 _21398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15733__A _13123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13850_ _11879_/A _13850_/B _13849_/X VGND VGND VPWR VPWR _13850_/X sky130_fd_sc_hd__and3_4
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12801_ _12801_/A _24010_/Q VGND VGND VPWR VPWR _12802_/C sky130_fd_sc_hd__or2_4
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13781_ _15517_/A _13749_/X _13781_/C VGND VGND VPWR VPWR _13781_/X sky130_fd_sc_hd__and3_4
XANTENNA__24278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21165__B2 _21159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22979_ _22961_/A _22979_/B VGND VGND VPWR VPWR _22981_/B sky130_fd_sc_hd__nand2_4
XANTENNA__18030__A1 _18022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15520_ _15519_/X VGND VGND VPWR VPWR _15520_/Y sky130_fd_sc_hd__inv_2
X_12732_ _12298_/A _12730_/X _12731_/X VGND VGND VPWR VPWR _12732_/X sky130_fd_sc_hd__and3_4
XFILLER_71_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15451_ _11969_/A _15428_/X _15435_/X _15442_/X _15450_/X VGND VGND VPWR VPWR _15451_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_31_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12663_ _12953_/A _12661_/X _12662_/X VGND VGND VPWR VPWR _12667_/B sky130_fd_sc_hd__and3_4
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16564__A _12001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _14372_/A _14398_/X _14401_/X VGND VGND VPWR VPWR _14402_/X sky130_fd_sc_hd__or3_4
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_4_0_HCLK clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_11614_ _11965_/A VGND VGND VPWR VPWR _11625_/A sky130_fd_sc_hd__buf_2
X_18170_ _18169_/Y _17527_/X _17535_/X VGND VGND VPWR VPWR _18170_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21468__A2 _21441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _15382_/A _15382_/B VGND VGND VPWR VPWR _15382_/X sky130_fd_sc_hd__and2_4
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12670_/A _12590_/X _12593_/X VGND VGND VPWR VPWR _12595_/C sky130_fd_sc_hd__and3_4
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23287__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ _14845_/Y _17115_/X _17120_/Y _17116_/X VGND VGND VPWR VPWR _17121_/X sky130_fd_sc_hd__o22a_4
X_14333_ _14450_/A _14310_/X _14317_/X _14324_/X _14332_/X VGND VGND VPWR VPWR _14333_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11545_ _20923_/A IRQ[4] VGND VGND VPWR VPWR _20169_/A sky130_fd_sc_hd__and2_4
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14084__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ _17036_/X _17047_/X _17051_/X VGND VGND VPWR VPWR _17052_/Y sky130_fd_sc_hd__o21ai_4
X_14264_ _14263_/X VGND VGND VPWR VPWR _14264_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22417__B2 _22409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16003_ _16003_/A _15997_/X _16003_/C VGND VGND VPWR VPWR _16003_/X sky130_fd_sc_hd__or3_4
XANTENNA__20428__B1 _24462_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13215_ _12372_/A VGND VGND VPWR VPWR _13252_/A sky130_fd_sc_hd__buf_2
XFILLER_152_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14195_ _14225_/A _23199_/Q VGND VGND VPWR VPWR _14195_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13146_ _13290_/A _13146_/B _13146_/C VGND VGND VPWR VPWR _13151_/B sky130_fd_sc_hd__and3_4
XANTENNA__21640__A2 _21634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13428__A _13327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13077_ _13051_/A VGND VGND VPWR VPWR _13099_/A sky130_fd_sc_hd__buf_2
X_17954_ _18411_/A _17591_/X _17807_/A _17643_/Y VGND VGND VPWR VPWR _17955_/B sky130_fd_sc_hd__o22a_4
XFILLER_39_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16905_ _16905_/A _16905_/B VGND VGND VPWR VPWR _16906_/B sky130_fd_sc_hd__or2_4
X_12028_ _11868_/X VGND VGND VPWR VPWR _12028_/X sky130_fd_sc_hd__buf_2
XANTENNA__21645__A _21624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17885_ _18562_/A _17885_/B VGND VGND VPWR VPWR _17885_/X sky130_fd_sc_hd__and2_4
XANTENNA__16739__A _12061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15643__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19624_ _19624_/A _19624_/B VGND VGND VPWR VPWR _19660_/A sky130_fd_sc_hd__or2_4
X_16836_ _15933_/X _16528_/A _16529_/Y VGND VGND VPWR VPWR _16836_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19555_ _19465_/A VGND VGND VPWR VPWR _19889_/A sky130_fd_sc_hd__buf_2
X_16767_ _16767_/A _16767_/B _16766_/X VGND VGND VPWR VPWR _16767_/X sky130_fd_sc_hd__and3_4
XANTENNA__21083__C _21184_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14259__A _11812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13979_ _12467_/A _13979_/B _13979_/C VGND VGND VPWR VPWR _13980_/C sky130_fd_sc_hd__and3_4
XFILLER_94_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21156__B2 _21152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13163__A _13276_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18506_ _18506_/A VGND VGND VPWR VPWR _18506_/X sky130_fd_sc_hd__buf_2
X_15718_ _15717_/X VGND VGND VPWR VPWR _15785_/A sky130_fd_sc_hd__inv_2
XFILLER_94_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19486_ _19823_/A VGND VGND VPWR VPWR _19525_/A sky130_fd_sc_hd__inv_2
X_16698_ _16691_/A _23793_/Q VGND VGND VPWR VPWR _16699_/C sky130_fd_sc_hd__or2_4
XFILLER_34_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22476__A _20937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18437_ _18483_/A _17609_/D VGND VGND VPWR VPWR _18437_/X sky130_fd_sc_hd__or2_4
XFILLER_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15649_ _15649_/A _15633_/X _15649_/C VGND VGND VPWR VPWR _15649_/X sky130_fd_sc_hd__or3_4
X_18368_ _18368_/A _18368_/B VGND VGND VPWR VPWR _18368_/X sky130_fd_sc_hd__or2_4
XANTENNA__22656__B2 _22655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17319_ _15382_/A VGND VGND VPWR VPWR _17319_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18299_ _18279_/X _18284_/Y _18289_/X _18297_/X _18298_/Y VGND VGND VPWR VPWR _18299_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_174_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12507__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20330_ _17650_/X _20847_/A _20638_/A _20329_/Y VGND VGND VPWR VPWR _20331_/A sky130_fd_sc_hd__a211o_4
XFILLER_31_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23081__A1 _19953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20261_ _20233_/Y VGND VGND VPWR VPWR _20261_/X sky130_fd_sc_hd__buf_2
XANTENNA__14722__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22000_ _22000_/A VGND VGND VPWR VPWR _22000_/X sky130_fd_sc_hd__buf_2
XFILLER_143_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20192_ _20192_/A _20191_/X VGND VGND VPWR VPWR _20192_/X sky130_fd_sc_hd__or2_4
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13338__A _13338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12242__A _12294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21919__B1 _15471_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23951_ _23983_/CLK _21255_/X VGND VGND VPWR VPWR _16270_/B sky130_fd_sc_hd__dfxtp_4
X_22902_ _12021_/Y _22849_/X _19909_/X _22901_/X VGND VGND VPWR VPWR _22902_/X sky130_fd_sc_hd__o22a_4
XFILLER_56_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23882_ _23531_/CLK _21390_/X VGND VGND VPWR VPWR _12747_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24405__CLK _23409_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22833_ _17353_/Y _22816_/X _22818_/X _22832_/X VGND VGND VPWR VPWR _22834_/B sky130_fd_sc_hd__o22a_4
XANTENNA__21147__B2 _21145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14169__A _14169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13073__A _12977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22764_ SYSTICKCLKDIV[6] _22763_/A _22762_/Y _22763_/Y VGND VGND VPWR VPWR _22768_/C
+ sky130_fd_sc_hd__o22a_4
XANTENNA__22895__B2 _20665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21715_ _21532_/X _21713_/X _23698_/Q _21710_/X VGND VGND VPWR VPWR _23698_/D sky130_fd_sc_hd__o22a_4
XFILLER_13_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22695_ _21528_/A _22694_/X _23123_/Q _22691_/X VGND VGND VPWR VPWR _23123_/D sky130_fd_sc_hd__o22a_4
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16384__A _16309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13801__A _15394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24434_ _23409_/CLK _24434_/D HRESETn VGND VGND VPWR VPWR _24434_/Q sky130_fd_sc_hd__dfrtp_4
X_21646_ _21584_/X _21641_/X _14345_/B _21645_/X VGND VGND VPWR VPWR _23740_/D sky130_fd_sc_hd__o22a_4
XFILLER_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22647__B2 _22641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21577_ _20801_/A VGND VGND VPWR VPWR _21577_/X sky130_fd_sc_hd__buf_2
X_24365_ _24368_/CLK _18999_/X HRESETn VGND VGND VPWR VPWR _18994_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__12417__A _12676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20528_ _20438_/A _20527_/X VGND VGND VPWR VPWR _20528_/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23316_ _23476_/CLK _23316_/D VGND VGND VPWR VPWR _11774_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_153_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24296_ _24357_/CLK _19282_/X HRESETn VGND VGND VPWR VPWR _24296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15728__A _13090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23010__A _18325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23247_ _23119_/CLK _23247_/D VGND VGND VPWR VPWR _16296_/B sky130_fd_sc_hd__dfxtp_4
X_20459_ _20398_/X _20445_/X _20714_/A _20458_/Y VGND VGND VPWR VPWR _20459_/X sky130_fd_sc_hd__a211o_4
XFILLER_137_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13000_ _12472_/A _13000_/B _12999_/X VGND VGND VPWR VPWR _13001_/C sky130_fd_sc_hd__and3_4
XFILLER_122_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21622__A2 _21620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23178_ _23852_/CLK _23178_/D VGND VGND VPWR VPWR _12794_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_79_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22129_ _20612_/A VGND VGND VPWR VPWR _22129_/X sky130_fd_sc_hd__buf_2
XANTENNA__13248__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18758__B _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14951_ _14922_/A _14880_/B VGND VGND VPWR VPWR _14951_/X sky130_fd_sc_hd__or2_4
XFILLER_134_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20189__A2 IRQ[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21386__B2 _21381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22583__B1 _15129_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11991__A _11943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13902_ _13697_/A _13900_/X _13901_/X VGND VGND VPWR VPWR _13902_/X sky130_fd_sc_hd__and3_4
XFILLER_130_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17670_ _17666_/X _17668_/Y _17669_/X VGND VGND VPWR VPWR _17671_/B sky130_fd_sc_hd__o21ai_4
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14882_ _14094_/A _14880_/X _14881_/X VGND VGND VPWR VPWR _14882_/X sky130_fd_sc_hd__and3_4
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16621_ _16621_/A _16621_/B VGND VGND VPWR VPWR _16621_/X sky130_fd_sc_hd__or2_4
X_13833_ _13657_/A _13831_/X _13833_/C VGND VGND VPWR VPWR _13837_/B sky130_fd_sc_hd__and3_4
XFILLER_169_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14079__A _12329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19340_ _19340_/A VGND VGND VPWR VPWR _19340_/X sky130_fd_sc_hd__buf_2
XFILLER_44_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16552_ _16593_/A VGND VGND VPWR VPWR _16558_/A sky130_fd_sc_hd__buf_2
X_13764_ _12616_/A _13764_/B _13763_/X VGND VGND VPWR VPWR _13764_/X sky130_fd_sc_hd__and3_4
XANTENNA__21689__A2 _21684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15503_ _12621_/X _15501_/X _15502_/X VGND VGND VPWR VPWR _15503_/X sky130_fd_sc_hd__and3_4
X_12715_ _12266_/A _12715_/B _12714_/X VGND VGND VPWR VPWR _12715_/X sky130_fd_sc_hd__or3_4
X_19271_ _19251_/B VGND VGND VPWR VPWR _19271_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16483_ _16507_/A _16480_/X _16482_/X VGND VGND VPWR VPWR _16483_/X sky130_fd_sc_hd__and3_4
XFILLER_31_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13695_ _13695_/A VGND VGND VPWR VPWR _13696_/A sky130_fd_sc_hd__buf_2
X_18222_ _18222_/A _17467_/B VGND VGND VPWR VPWR _18225_/B sky130_fd_sc_hd__and2_4
X_15434_ _15411_/A _15432_/X _15434_/C VGND VGND VPWR VPWR _15434_/X sky130_fd_sc_hd__and3_4
X_12646_ _12646_/A _12646_/B VGND VGND VPWR VPWR _12648_/B sky130_fd_sc_hd__or2_4
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14526__B _14462_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18153_ _18545_/A VGND VGND VPWR VPWR _18282_/A sky130_fd_sc_hd__buf_2
X_15365_ _13695_/A _15365_/B _15364_/X VGND VGND VPWR VPWR _15365_/X sky130_fd_sc_hd__and3_4
X_12577_ _12367_/A VGND VGND VPWR VPWR _12578_/A sky130_fd_sc_hd__buf_2
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21310__B2 _21300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17104_ _17089_/X _17095_/X _17099_/Y _17104_/D VGND VGND VPWR VPWR _17105_/A sky130_fd_sc_hd__or4_4
X_14316_ _11914_/A _14316_/B _14316_/C VGND VGND VPWR VPWR _14316_/X sky130_fd_sc_hd__and3_4
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11528_ _11528_/A _11528_/B VGND VGND VPWR VPWR _19054_/A sky130_fd_sc_hd__or2_4
X_18084_ _17876_/X _18081_/Y _17833_/A _18083_/Y VGND VGND VPWR VPWR _18084_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15296_ _13788_/A _15292_/X _15295_/X VGND VGND VPWR VPWR _15296_/X sky130_fd_sc_hd__or3_4
XANTENNA__21861__A2 _21851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14879__A1 _14012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17035_ _17035_/A VGND VGND VPWR VPWR _17251_/B sky130_fd_sc_hd__buf_2
X_14247_ _14254_/A _23711_/Q VGND VGND VPWR VPWR _14249_/B sky130_fd_sc_hd__or2_4
XANTENNA__15638__A _13885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14178_ _13694_/A VGND VGND VPWR VPWR _14616_/A sky130_fd_sc_hd__buf_2
XFILLER_124_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13158__A _12858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13129_ _12698_/A _13129_/B _13129_/C VGND VGND VPWR VPWR _13129_/X sky130_fd_sc_hd__and3_4
XANTENNA__18490__A1 _17805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12062__A _11963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18986_ _19016_/A VGND VGND VPWR VPWR _18987_/A sky130_fd_sc_hd__buf_2
XFILLER_112_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17937_ _17825_/X _17209_/X _17814_/X _17213_/X VGND VGND VPWR VPWR _17937_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12997__A _12877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22574__B1 _13721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15373__A _11659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17868_ _18265_/A VGND VGND VPWR VPWR _17869_/A sky130_fd_sc_hd__buf_2
XANTENNA__24129__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19607_ _19719_/A VGND VGND VPWR VPWR _19607_/X sky130_fd_sc_hd__buf_2
X_16819_ _11671_/X _16819_/B _16818_/X VGND VGND VPWR VPWR _16819_/X sky130_fd_sc_hd__and3_4
XFILLER_54_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17799_ _18335_/A _17258_/A VGND VGND VPWR VPWR _17799_/X sky130_fd_sc_hd__and2_4
XANTENNA__21129__B2 _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19538_ _19538_/A VGND VGND VPWR VPWR _19883_/A sky130_fd_sc_hd__buf_2
XFILLER_35_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19469_ _19700_/A VGND VGND VPWR VPWR _19469_/X sky130_fd_sc_hd__buf_2
XFILLER_59_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14717__A _13823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21500_ _21280_/X _21499_/X _23812_/Q _21496_/X VGND VGND VPWR VPWR _23812_/D sky130_fd_sc_hd__o22a_4
XFILLER_167_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22480_ _22480_/A VGND VGND VPWR VPWR _22480_/X sky130_fd_sc_hd__buf_2
XFILLER_148_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21431_ _21431_/A VGND VGND VPWR VPWR _21431_/X sky130_fd_sc_hd__buf_2
XFILLER_148_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16308__A1 _16130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21301__B2 _21300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24150_ _24302_/CLK _24150_/D HRESETn VGND VGND VPWR VPWR _24150_/Q sky130_fd_sc_hd__dfrtp_4
X_21362_ _21322_/A VGND VGND VPWR VPWR _21362_/X sky130_fd_sc_hd__buf_2
XANTENNA__21852__A2 _21851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20313_ _20257_/X VGND VGND VPWR VPWR _20313_/X sky130_fd_sc_hd__buf_2
X_23101_ _23101_/CLK _23101_/D VGND VGND VPWR VPWR _13929_/B sky130_fd_sc_hd__dfxtp_4
X_24081_ _23761_/CLK _21041_/X VGND VGND VPWR VPWR _24081_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15548__A _12427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21293_ _21238_/A VGND VGND VPWR VPWR _21293_/X sky130_fd_sc_hd__buf_2
XANTENNA__14334__A3 _14303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14452__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21065__B1 _24064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23032_ _18210_/X _23055_/B VGND VGND VPWR VPWR _23033_/C sky130_fd_sc_hd__or2_4
XFILLER_89_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20244_ _20863_/A _20244_/B VGND VGND VPWR VPWR _20244_/X sky130_fd_sc_hd__and2_4
XFILLER_118_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22801__A1 _18738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18481__A1 _18111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20175_ _20161_/Y _20162_/Y _11560_/X _20174_/X VGND VGND VPWR VPWR _20175_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16379__A _13416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21368__B2 _21331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23934_ _23582_/CLK _23934_/D VGND VGND VPWR VPWR _13732_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23865_ _23641_/CLK _21414_/X VGND VGND VPWR VPWR _14761_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20591__A2 _20577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22317__B1 _14779_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22816_ _22815_/X VGND VGND VPWR VPWR _22816_/X sky130_fd_sc_hd__buf_2
X_23796_ _23668_/CLK _23796_/D VGND VGND VPWR VPWR _23796_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22747_ _23086_/A _22746_/X _22945_/A _19402_/X VGND VGND VPWR VPWR _22747_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21540__B2 _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12500_ _12871_/A _12500_/B VGND VGND VPWR VPWR _12500_/X sky130_fd_sc_hd__or2_4
X_13480_ _12514_/A _13480_/B VGND VGND VPWR VPWR _13480_/X sky130_fd_sc_hd__or2_4
XFILLER_125_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_66_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR _23126_/CLK sky130_fd_sc_hd__clkbuf_1
X_22678_ _22471_/X _22672_/X _14523_/B _22676_/X VGND VGND VPWR VPWR _22678_/X sky130_fd_sc_hd__o22a_4
X_12431_ _14905_/A VGND VGND VPWR VPWR _14108_/A sky130_fd_sc_hd__buf_2
X_24417_ _24419_/CLK _24417_/D HRESETn VGND VGND VPWR VPWR _20727_/A sky130_fd_sc_hd__dfrtp_4
X_21629_ _21556_/X _21627_/X _23752_/Q _21624_/X VGND VGND VPWR VPWR _23752_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19497__B1 HRDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12147__A _16053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15150_ _14994_/A _15150_/B VGND VGND VPWR VPWR _15150_/X sky130_fd_sc_hd__or2_4
X_12362_ _12362_/A VGND VGND VPWR VPWR _12923_/A sky130_fd_sc_hd__buf_2
X_24348_ _24382_/CLK _24348_/D HRESETn VGND VGND VPWR VPWR _11522_/A sky130_fd_sc_hd__dfstp_4
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14101_ _11623_/A _23199_/Q VGND VGND VPWR VPWR _14101_/X sky130_fd_sc_hd__or2_4
XFILLER_126_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11986__A _16742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12293_ _12735_/A _12293_/B VGND VGND VPWR VPWR _12293_/X sky130_fd_sc_hd__or2_4
X_15081_ _15081_/A _15081_/B _15081_/C VGND VGND VPWR VPWR _15082_/C sky130_fd_sc_hd__and3_4
X_24279_ _24292_/CLK _24279_/D HRESETn VGND VGND VPWR VPWR _19228_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14032_ _13696_/A _14032_/B _14031_/X VGND VGND VPWR VPWR _14032_/X sky130_fd_sc_hd__and3_4
XANTENNA__15177__B _15177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18840_ _18840_/A VGND VGND VPWR VPWR _18840_/X sky130_fd_sc_hd__buf_2
XFILLER_110_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21195__A _21195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18771_ _19973_/A _18769_/X _19962_/B _18770_/X VGND VGND VPWR VPWR _18771_/X sky130_fd_sc_hd__o22a_4
X_15983_ _15993_/A _15981_/X _15983_/C VGND VGND VPWR VPWR _15983_/X sky130_fd_sc_hd__and3_4
XFILLER_121_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22556__B1 _12599_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17722_ _17721_/A _17427_/X VGND VGND VPWR VPWR _17723_/A sky130_fd_sc_hd__or2_4
XANTENNA__15193__A _14773_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22020__A2 _22017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13706__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14934_ _14967_/A _14934_/B VGND VGND VPWR VPWR _14934_/X sky130_fd_sc_hd__or2_4
XFILLER_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12610__A _12610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18775__A2 _18774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19972__A1 _17974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17653_ _17652_/X VGND VGND VPWR VPWR _17653_/X sky130_fd_sc_hd__buf_2
XANTENNA__21923__A _21923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14865_ _14881_/A _23990_/Q VGND VGND VPWR VPWR _14866_/C sky130_fd_sc_hd__or2_4
XFILLER_29_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16604_ _11686_/X VGND VGND VPWR VPWR _16683_/A sky130_fd_sc_hd__buf_2
XANTENNA__22738__B _22737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13816_ _14319_/A _23997_/Q VGND VGND VPWR VPWR _13817_/C sky130_fd_sc_hd__or2_4
X_17584_ _17551_/B VGND VGND VPWR VPWR _17968_/B sky130_fd_sc_hd__inv_2
X_14796_ _14675_/A _14728_/B VGND VGND VPWR VPWR _14797_/C sky130_fd_sc_hd__or2_4
XFILLER_91_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19323_ _19957_/A VGND VGND VPWR VPWR _19324_/A sky130_fd_sc_hd__buf_2
XFILLER_90_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16535_ _16534_/X _16609_/B VGND VGND VPWR VPWR _16535_/X sky130_fd_sc_hd__or2_4
X_13747_ _12578_/A _13747_/B _13747_/C VGND VGND VPWR VPWR _13748_/C sky130_fd_sc_hd__or3_4
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13441__A _13441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21531__B2 _21525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19254_ _24305_/Q _19254_/B VGND VGND VPWR VPWR _19255_/B sky130_fd_sc_hd__and2_4
X_16466_ _13367_/A VGND VGND VPWR VPWR _16507_/A sky130_fd_sc_hd__buf_2
X_13678_ _15439_/A _13775_/B VGND VGND VPWR VPWR _13678_/X sky130_fd_sc_hd__or2_4
X_18205_ _18198_/X _18202_/Y _17224_/X _18204_/X VGND VGND VPWR VPWR _18205_/X sky130_fd_sc_hd__a211o_4
X_15417_ _14329_/A _15474_/B VGND VGND VPWR VPWR _15418_/C sky130_fd_sc_hd__or2_4
X_12629_ _12976_/A _12620_/X _12629_/C VGND VGND VPWR VPWR _12640_/B sky130_fd_sc_hd__or3_4
XFILLER_129_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19488__B1 HRDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19185_ _19185_/A VGND VGND VPWR VPWR _19185_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22087__A2 _22060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16397_ _16007_/X _16397_/B VGND VGND VPWR VPWR _16399_/B sky130_fd_sc_hd__or2_4
XANTENNA__22754__A1_N SYSTICKCLKDIV[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18136_ _17111_/X _18130_/Y _17224_/X _18135_/Y VGND VGND VPWR VPWR _18136_/X sky130_fd_sc_hd__a211o_4
X_15348_ _15318_/A _23896_/Q VGND VGND VPWR VPWR _15348_/X sky130_fd_sc_hd__or2_4
XANTENNA__22904__D _22904_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18160__B1 _17811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18067_ _18020_/X _18063_/X _18065_/X _18066_/X VGND VGND VPWR VPWR _18067_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15368__A _11735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15279_ _14897_/X _15279_/B _15278_/X VGND VGND VPWR VPWR _15279_/X sky130_fd_sc_hd__and3_4
XANTENNA__14272__A _14272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24250__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17018_ _17025_/A VGND VGND VPWR VPWR _17018_/X sky130_fd_sc_hd__buf_2
XFILLER_99_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18969_ _18963_/X _18965_/X _18966_/Y _18968_/X VGND VGND VPWR VPWR _18969_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13616__A _13990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22011__A2 _22010_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12520__A _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21980_ _21872_/X _21974_/X _14440_/B _21978_/X VGND VGND VPWR VPWR _23547_/D sky130_fd_sc_hd__o22a_4
XFILLER_2_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22929__A _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13335__B _23718_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20931_ _18681_/X _20313_/X _20780_/X _20930_/Y VGND VGND VPWR VPWR _20931_/X sky130_fd_sc_hd__a211o_4
XFILLER_6_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20862_ _20772_/X _20860_/X _24092_/Q _20861_/X VGND VGND VPWR VPWR _20862_/X sky130_fd_sc_hd__o22a_4
X_23650_ _23650_/CLK _23650_/D VGND VGND VPWR VPWR _15512_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22601_ _22608_/A VGND VGND VPWR VPWR _22601_/X sky130_fd_sc_hd__buf_2
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12263__A1 _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20793_ _20930_/A _20792_/X VGND VGND VPWR VPWR _20793_/Y sky130_fd_sc_hd__nor2_4
X_23581_ _23582_/CLK _23581_/D VGND VGND VPWR VPWR _13897_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14447__A _13601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22532_ _22478_/X _22529_/X _15300_/B _22526_/X VGND VGND VPWR VPWR _23224_/D sky130_fd_sc_hd__o22a_4
XFILLER_23_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14166__B _23807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22463_ _22461_/X _22462_/X _23263_/Q _22457_/X VGND VGND VPWR VPWR _22463_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21286__B1 _15470_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20089__B2 _19951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24202_ _24182_/CLK _24202_/D HRESETn VGND VGND VPWR VPWR _11928_/A sky130_fd_sc_hd__dfrtp_4
X_21414_ _21307_/X _21412_/X _14761_/B _21409_/X VGND VGND VPWR VPWR _21414_/X sky130_fd_sc_hd__o22a_4
XFILLER_159_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21825__A2 _21815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22394_ _22358_/A VGND VGND VPWR VPWR _22394_/X sky130_fd_sc_hd__buf_2
XFILLER_163_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21345_ _21338_/A VGND VGND VPWR VPWR _21345_/X sky130_fd_sc_hd__buf_2
X_24133_ _24471_/CLK _24133_/D HRESETn VGND VGND VPWR VPWR _16971_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15278__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21276_ _21264_/A VGND VGND VPWR VPWR _21276_/X sky130_fd_sc_hd__buf_2
XFILLER_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24064_ _23587_/CLK _24064_/D VGND VGND VPWR VPWR _24064_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20912__A _20977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_HCLK clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23015_ _18299_/X _23003_/B VGND VGND VPWR VPWR _23015_/X sky130_fd_sc_hd__or2_4
X_20227_ _20226_/X VGND VGND VPWR VPWR _20358_/A sky130_fd_sc_hd__buf_2
XANTENNA__22250__A2 _22244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20158_ IRQ[17] VGND VGND VPWR VPWR _20158_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22002__A2 _21996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19403__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12980_ _12979_/X VGND VGND VPWR VPWR _12980_/X sky130_fd_sc_hd__buf_2
X_20089_ _18593_/X _20079_/X _20088_/Y _19951_/X VGND VGND VPWR VPWR _20089_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12430__A _13792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23917_ _24045_/CLK _21336_/X VGND VGND VPWR VPWR _16132_/B sky130_fd_sc_hd__dfxtp_4
X_11931_ _11931_/A VGND VGND VPWR VPWR _11932_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15741__A _13067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21761__B2 _21760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14650_ _14658_/A _23450_/Q VGND VGND VPWR VPWR _14650_/X sky130_fd_sc_hd__or2_4
X_23848_ _23592_/CLK _23848_/D VGND VGND VPWR VPWR _23848_/Q sky130_fd_sc_hd__dfxtp_4
X_11862_ _13689_/A VGND VGND VPWR VPWR _13046_/A sky130_fd_sc_hd__buf_2
XFILLER_33_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _13601_/A _13707_/B VGND VGND VPWR VPWR _13601_/X sky130_fd_sc_hd__or2_4
XANTENNA__24123__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14581_ _14302_/A _14580_/X VGND VGND VPWR VPWR _14581_/X sky130_fd_sc_hd__and2_4
XPHY_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23779_ _23111_/CLK _21569_/X VGND VGND VPWR VPWR _15797_/B sky130_fd_sc_hd__dfxtp_4
X_11793_ _11792_/X _11793_/B VGND VGND VPWR VPWR _11793_/X sky130_fd_sc_hd__or2_4
XFILLER_14_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16320_ _13407_/A _16320_/B _16319_/X VGND VGND VPWR VPWR _16328_/B sky130_fd_sc_hd__or3_4
XANTENNA__13261__A _15517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13532_ _13532_/A _23973_/Q VGND VGND VPWR VPWR _13532_/X sky130_fd_sc_hd__or2_4
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14076__B _24096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16251_ _16282_/A _16251_/B VGND VGND VPWR VPWR _16251_/X sky130_fd_sc_hd__or2_4
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13463_ _13431_/X _23845_/Q VGND VGND VPWR VPWR _13463_/X sky130_fd_sc_hd__or2_4
XFILLER_158_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22069__A2 _22067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15202_ _14614_/A _15202_/B _15201_/X VGND VGND VPWR VPWR _15202_/X sky130_fd_sc_hd__and3_4
X_12414_ _13542_/A _12412_/X _12413_/X VGND VGND VPWR VPWR _12415_/C sky130_fd_sc_hd__and3_4
X_16182_ _16181_/X _24045_/Q VGND VGND VPWR VPWR _16185_/B sky130_fd_sc_hd__or2_4
XANTENNA__21816__A2 _21815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13394_ _13385_/A _23846_/Q VGND VGND VPWR VPWR _13395_/C sky130_fd_sc_hd__or2_4
XANTENNA__20094__A _20093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14804__B _14721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15133_ _14169_/A VGND VGND VPWR VPWR _15267_/A sky130_fd_sc_hd__buf_2
XANTENNA__15188__A _14771_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12345_ _12829_/A _23788_/Q VGND VGND VPWR VPWR _12346_/C sky130_fd_sc_hd__or2_4
XFILLER_5_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14092__A _14003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12605__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19941_ _19938_/X _24168_/Q _19939_/X _20917_/B VGND VGND VPWR VPWR _24168_/D sky130_fd_sc_hd__o22a_4
X_15064_ _15078_/A _15064_/B _15063_/X VGND VGND VPWR VPWR _15064_/X sky130_fd_sc_hd__and3_4
X_12276_ _12727_/A _12389_/B VGND VGND VPWR VPWR _12276_/X sky130_fd_sc_hd__or2_4
XANTENNA__20822__A _21007_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18499__A _18019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14015_ _14014_/X VGND VGND VPWR VPWR _14086_/A sky130_fd_sc_hd__inv_2
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17248__A2 _18734_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15916__A _15912_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19872_ _19871_/X VGND VGND VPWR VPWR _19872_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20252__A1 _18780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18823_ _17272_/X _18817_/X _24444_/Q _18818_/X VGND VGND VPWR VPWR _24444_/D sky130_fd_sc_hd__o22a_4
XFILLER_95_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13436__A _13462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15966_ _15956_/A VGND VGND VPWR VPWR _15967_/A sky130_fd_sc_hd__buf_2
X_18754_ _17809_/A _11633_/X VGND VGND VPWR VPWR _18754_/Y sky130_fd_sc_hd__nor2_4
XFILLER_23_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21201__B1 _23980_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14482__A2 _11629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19945__A1 _19920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17705_ _17770_/A _17701_/Y _17702_/X _17704_/Y VGND VGND VPWR VPWR _17705_/X sky130_fd_sc_hd__a211o_4
XANTENNA__19945__B2 _22737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14917_ _14772_/A VGND VGND VPWR VPWR _14922_/A sky130_fd_sc_hd__buf_2
X_15897_ _13496_/A _15841_/B VGND VGND VPWR VPWR _15897_/X sky130_fd_sc_hd__or2_4
X_18685_ _18684_/X VGND VGND VPWR VPWR _18685_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20555__A2 _20443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17956__B1 _17890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16747__A _12108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21752__B2 _21717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14848_ _14847_/X VGND VGND VPWR VPWR _14848_/Y sky130_fd_sc_hd__inv_2
X_17636_ _17636_/A _17636_/B VGND VGND VPWR VPWR _17637_/D sky130_fd_sc_hd__nor2_4
XFILLER_24_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17567_ _17047_/A _17566_/X _17050_/X VGND VGND VPWR VPWR _17567_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14779_ _14674_/A _14779_/B VGND VGND VPWR VPWR _14781_/B sky130_fd_sc_hd__or2_4
XANTENNA__18962__A _20192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14267__A _14267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21504__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13171__A _13303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16518_ _16370_/X _16514_/X _16518_/C VGND VGND VPWR VPWR _16519_/C sky130_fd_sc_hd__or3_4
X_19306_ _24284_/Q _19233_/B _19305_/Y VGND VGND VPWR VPWR _24284_/D sky130_fd_sc_hd__o21a_4
XFILLER_149_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20712__C1 _20711_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17498_ _17496_/Y _17497_/X VGND VGND VPWR VPWR _18290_/A sky130_fd_sc_hd__or2_4
XANTENNA__17184__A1 _17015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22484__A _22169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16449_ _11865_/X _16448_/X VGND VGND VPWR VPWR _16449_/X sky130_fd_sc_hd__and2_4
X_19237_ _19237_/A _19237_/B VGND VGND VPWR VPWR _19237_/X sky130_fd_sc_hd__and2_4
XFILLER_20_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17578__A _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19168_ _19158_/A _19158_/B _19167_/Y VGND VGND VPWR VPWR _24337_/D sky130_fd_sc_hd__o21a_4
XFILLER_173_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18119_ _17095_/X _18119_/B _18119_/C _18119_/D VGND VGND VPWR VPWR _18120_/A sky130_fd_sc_hd__or4_4
XANTENNA__18684__A1 _18064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15098__A _15106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19099_ _19099_/A VGND VGND VPWR VPWR _19099_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12515__A _12515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21130_ _21004_/X _21125_/X _14859_/B _21086_/X VGND VGND VPWR VPWR _21130_/X sky130_fd_sc_hd__o22a_4
XFILLER_132_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15826__A _12884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21061_ _20693_/X _21059_/X _15823_/B _21056_/X VGND VGND VPWR VPWR _21061_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22232__A2 _22230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24144__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20012_ _20012_/A VGND VGND VPWR VPWR _20012_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13346__A _12834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24146__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19936__B2 _20844_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21963_ _21843_/X _21960_/X _23559_/Q _21957_/X VGND VGND VPWR VPWR _23559_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20546__A2 _20545_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21743__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15561__A _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23702_ _23194_/CLK _23702_/D VGND VGND VPWR VPWR _23702_/Q sky130_fd_sc_hd__dfxtp_4
X_20914_ _22158_/A VGND VGND VPWR VPWR _21304_/A sky130_fd_sc_hd__buf_2
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21894_ _21923_/A VGND VGND VPWR VPWR _21909_/A sky130_fd_sc_hd__buf_2
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23633_ _23761_/CLK _23633_/D VGND VGND VPWR VPWR _23633_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22299__A2 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20845_/A _20843_/X _20844_/X VGND VGND VPWR VPWR _20845_/X sky130_fd_sc_hd__and3_4
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14177__A _15321_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23170__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24296__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23564_ _23500_/CLK _21956_/X VGND VGND VPWR VPWR _12376_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20776_ _20776_/A _20671_/A VGND VGND VPWR VPWR _20777_/C sky130_fd_sc_hd__or2_4
XFILLER_50_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22394__A _22358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22515_ _22508_/A VGND VGND VPWR VPWR _22515_/X sky130_fd_sc_hd__buf_2
XFILLER_167_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23495_ _24039_/CLK _22063_/X VGND VGND VPWR VPWR _23495_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16392__A _16011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22446_ _22444_/X _22438_/X _13273_/B _22445_/X VGND VGND VPWR VPWR _22446_/X sky130_fd_sc_hd__o22a_4
XFILLER_164_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22377_ _22122_/X _22376_/X _23305_/Q _22373_/X VGND VGND VPWR VPWR _22377_/X sky130_fd_sc_hd__o22a_4
XFILLER_136_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24116_ _23668_/CLK _24116_/D VGND VGND VPWR VPWR _24116_/Q sky130_fd_sc_hd__dfxtp_4
X_12130_ _11760_/X _12126_/X _12130_/C VGND VGND VPWR VPWR _12131_/C sky130_fd_sc_hd__or3_4
X_21328_ _21243_/X _21327_/X _23923_/Q _21324_/X VGND VGND VPWR VPWR _23923_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21738__A _21724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21259_ _20464_/A VGND VGND VPWR VPWR _21259_/X sky130_fd_sc_hd__buf_2
XFILLER_151_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24047_ _23119_/CLK _21096_/X VGND VGND VPWR VPWR _16259_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15736__A _12766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12061_ _12061_/A _12061_/B _12061_/C VGND VGND VPWR VPWR _12067_/B sky130_fd_sc_hd__and3_4
XANTENNA__18427__B2 _18426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20234__A1 _16915_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15455__B _15455_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15820_ _12848_/A _15820_/B VGND VGND VPWR VPWR _15820_/X sky130_fd_sc_hd__or2_4
XANTENNA__13256__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21982__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15751_ _12641_/A _15751_/B _15750_/X VGND VGND VPWR VPWR _15783_/B sky130_fd_sc_hd__or3_4
XANTENNA__19927__B2 _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21473__A _21506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12963_ _12951_/A _12963_/B VGND VGND VPWR VPWR _12965_/B sky130_fd_sc_hd__or2_4
XFILLER_46_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16567__A _11951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14702_ _14613_/X _14701_/Y VGND VGND VPWR VPWR _14703_/A sky130_fd_sc_hd__or2_4
X_11914_ _11914_/A VGND VGND VPWR VPWR _11915_/A sky130_fd_sc_hd__buf_2
X_18470_ _17396_/B _18469_/X VGND VGND VPWR VPWR _18470_/X sky130_fd_sc_hd__or2_4
X_15682_ _12311_/A _15682_/B VGND VGND VPWR VPWR _15682_/X sky130_fd_sc_hd__or2_4
X_12894_ _12894_/A _23401_/Q VGND VGND VPWR VPWR _12896_/B sky130_fd_sc_hd__or2_4
XANTENNA__22492__A2_N _22491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17421_ _14084_/X _17421_/B VGND VGND VPWR VPWR _17421_/X sky130_fd_sc_hd__or2_4
X_14633_ _14820_/A _14633_/B VGND VGND VPWR VPWR _14633_/X sky130_fd_sc_hd__or2_4
X_11845_ _11792_/X _11845_/B VGND VGND VPWR VPWR _11845_/X sky130_fd_sc_hd__or2_4
XPHY_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18782__A _17048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _17272_/X _17306_/A _17312_/Y _17351_/X VGND VGND VPWR VPWR _18418_/A sky130_fd_sc_hd__a211o_4
XPHY_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14564_ _12454_/A _14564_/B VGND VGND VPWR VPWR _14564_/X sky130_fd_sc_hd__or2_4
XPHY_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _12138_/A _11765_/X _11775_/X VGND VGND VPWR VPWR _11776_/X sky130_fd_sc_hd__or3_4
XANTENNA__17166__A1 _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _11889_/X _16303_/B VGND VGND VPWR VPWR _16303_/X sky130_fd_sc_hd__or2_4
XFILLER_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13515_ _12970_/A VGND VGND VPWR VPWR _13515_/X sky130_fd_sc_hd__buf_2
XANTENNA__23663__CLK _23246_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17398__A _17398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17283_ _14549_/Y _17303_/B VGND VGND VPWR VPWR _18603_/B sky130_fd_sc_hd__or2_4
X_14495_ _14378_/A _14495_/B VGND VGND VPWR VPWR _14495_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_36_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_72_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19022_ _19016_/X _19019_/X _19020_/Y _19021_/X VGND VGND VPWR VPWR _19022_/X sky130_fd_sc_hd__o22a_4
X_16234_ _16219_/A _16150_/B VGND VGND VPWR VPWR _16234_/X sky130_fd_sc_hd__or2_4
XFILLER_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13446_ _12863_/A _13512_/B VGND VGND VPWR VPWR _13446_/X sky130_fd_sc_hd__or2_4
XFILLER_70_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16165_ _16164_/X _16090_/B VGND VGND VPWR VPWR _16165_/X sky130_fd_sc_hd__or2_4
X_13377_ _13377_/A VGND VGND VPWR VPWR _13398_/A sky130_fd_sc_hd__buf_2
XFILLER_127_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15116_ _11666_/X _15084_/X _15116_/C VGND VGND VPWR VPWR _15116_/X sky130_fd_sc_hd__and3_4
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21648__A _21608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12328_ _12580_/A VGND VGND VPWR VPWR _12329_/A sky130_fd_sc_hd__buf_2
XFILLER_86_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16096_ _16096_/A VGND VGND VPWR VPWR _16112_/A sky130_fd_sc_hd__buf_2
XFILLER_114_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19924_ _19924_/A VGND VGND VPWR VPWR _22745_/A sky130_fd_sc_hd__buf_2
X_15047_ _15047_/A VGND VGND VPWR VPWR _15047_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15646__A _13923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12259_ _12702_/A _12259_/B VGND VGND VPWR VPWR _12259_/X sky130_fd_sc_hd__or2_4
XANTENNA__22214__A2 _22208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18022__A _18148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14550__A _14482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24169__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19855_ _19854_/X VGND VGND VPWR VPWR _19855_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21973__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18806_ _12980_/X _18803_/X _11556_/A _18804_/X VGND VGND VPWR VPWR _24457_/D sky130_fd_sc_hd__o22a_4
XFILLER_95_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12070__A _11963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19786_ _19788_/A _19811_/B _19743_/Y VGND VGND VPWR VPWR _19786_/X sky130_fd_sc_hd__a21o_4
X_16998_ _17655_/A _17008_/A VGND VGND VPWR VPWR _16999_/B sky130_fd_sc_hd__or2_4
XFILLER_23_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18737_ _18461_/A _17624_/Y _18733_/X _18736_/Y VGND VGND VPWR VPWR _18737_/X sky130_fd_sc_hd__a211o_4
X_15949_ _11917_/X VGND VGND VPWR VPWR _15952_/A sky130_fd_sc_hd__buf_2
XANTENNA__16477__A _16163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21725__B2 _21724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18668_ _18574_/X _18666_/X _24474_/Q _18667_/X VGND VGND VPWR VPWR _18668_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14709__B _14779_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19788__A _19788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17619_ _17315_/Y _18651_/B _17292_/X VGND VGND VPWR VPWR _17620_/B sky130_fd_sc_hd__o21a_4
Xclkbuf_7_118_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR _23997_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18599_ _17618_/Y _18599_/B VGND VGND VPWR VPWR _18599_/X sky130_fd_sc_hd__or2_4
X_20630_ _20535_/X _20629_/X VGND VGND VPWR VPWR _20630_/X sky130_fd_sc_hd__or2_4
XANTENNA__17157__A1 _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22150__B2 _22142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20561_ _20307_/X _20561_/B VGND VGND VPWR VPWR _20561_/X sky130_fd_sc_hd__and2_4
XANTENNA__14725__A _11913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22300_ _22132_/X _22294_/X _23365_/Q _22298_/X VGND VGND VPWR VPWR _22300_/X sky130_fd_sc_hd__o22a_4
X_23280_ _23760_/CLK _22422_/X VGND VGND VPWR VPWR _16387_/B sky130_fd_sc_hd__dfxtp_4
X_20492_ _11554_/A VGND VGND VPWR VPWR _20494_/A sky130_fd_sc_hd__inv_2
XANTENNA__22942__A _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22231_ _22097_/X _22230_/X _12158_/B _22227_/X VGND VGND VPWR VPWR _23411_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12245__A _13301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24325__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19854__B1 _21370_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22162_ _22161_/X _22159_/X _14731_/B _22154_/X VGND VGND VPWR VPWR _22162_/X sky130_fd_sc_hd__o22a_4
XFILLER_156_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21113_ _20693_/X _21111_/X _15799_/B _21108_/X VGND VGND VPWR VPWR _21113_/X sky130_fd_sc_hd__o22a_4
X_22093_ _22118_/A VGND VGND VPWR VPWR _22106_/A sky130_fd_sc_hd__buf_2
XANTENNA__14460__A _12455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21044_ _20416_/X _21038_/X _16283_/B _21042_/X VGND VGND VPWR VPWR _24079_/D sky130_fd_sc_hd__o22a_4
XFILLER_8_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21293__A _21238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22995_ _17906_/A _17906_/B _22949_/A _18248_/C VGND VGND VPWR VPWR _22995_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21716__B2 _21710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15291__A _14269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13804__A _12485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21946_ _21960_/A VGND VGND VPWR VPWR _21946_/X sky130_fd_sc_hd__buf_2
XFILLER_27_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21192__A2 _21191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21877_ _20938_/A VGND VGND VPWR VPWR _21877_/X sky130_fd_sc_hd__buf_2
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11630_/A VGND VGND VPWR VPWR _11631_/A sky130_fd_sc_hd__buf_2
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _24096_/CLK _23616_/D VGND VGND VPWR VPWR _23616_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ _20676_/X _20825_/Y _20827_/X _19090_/Y _20731_/X VGND VGND VPWR VPWR _20828_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20637__A _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23547_ _23323_/CLK _23547_/D VGND VGND VPWR VPWR _14440_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _20161_/A IRQ[13] _11560_/X VGND VGND VPWR VPWR _11561_/X sky130_fd_sc_hd__a21o_4
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20759_ _20644_/X _20757_/X _19237_/A _20758_/X VGND VGND VPWR VPWR _20759_/X sky130_fd_sc_hd__o22a_4
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14635__A _14635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13300_ _13300_/A _13364_/B VGND VGND VPWR VPWR _13302_/B sky130_fd_sc_hd__or2_4
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ _14280_/A _14278_/X _14280_/C VGND VGND VPWR VPWR _14284_/B sky130_fd_sc_hd__and3_4
XFILLER_11_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23478_ _23864_/CLK _23478_/D VGND VGND VPWR VPWR _23478_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14354__B _24028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13231_ _13200_/X _23975_/Q VGND VGND VPWR VPWR _13231_/X sky130_fd_sc_hd__or2_4
X_22429_ _22428_/X _22426_/X _16090_/B _22421_/X VGND VGND VPWR VPWR _22429_/X sky130_fd_sc_hd__o22a_4
XFILLER_136_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18648__A1 _17980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13162_ _13279_/A _23975_/Q VGND VGND VPWR VPWR _13162_/X sky130_fd_sc_hd__or2_4
XFILLER_152_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24311__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11994__A _11990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12113_ _16079_/A VGND VGND VPWR VPWR _16608_/A sky130_fd_sc_hd__buf_2
XFILLER_123_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13093_ _12641_/A _13093_/B _13093_/C VGND VGND VPWR VPWR _13125_/B sky130_fd_sc_hd__or3_4
XANTENNA__14370__A _12583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17970_ _18407_/A _17554_/B VGND VGND VPWR VPWR _17970_/Y sky130_fd_sc_hd__nor2_4
XFILLER_111_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20207__B2 _19951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16921_ _16921_/A VGND VGND VPWR VPWR _16922_/C sky130_fd_sc_hd__buf_2
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12044_ _16568_/A VGND VGND VPWR VPWR _16592_/A sky130_fd_sc_hd__buf_2
XFILLER_46_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12602__B _23787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21955__B2 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19640_ _24166_/Q _19457_/X HRDATA[18] _19454_/X VGND VGND VPWR VPWR _19640_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18820__A1 _14261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16852_ _16852_/A _16846_/X _16850_/X _16852_/D VGND VGND VPWR VPWR _16852_/X sky130_fd_sc_hd__and4_4
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15803_ _12863_/A _15803_/B VGND VGND VPWR VPWR _15803_/X sky130_fd_sc_hd__or2_4
XFILLER_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19571_ _19439_/A VGND VGND VPWR VPWR _19571_/X sky130_fd_sc_hd__buf_2
X_16783_ _16611_/A _23569_/Q VGND VGND VPWR VPWR _16783_/X sky130_fd_sc_hd__or2_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13995_ _11912_/A _13993_/X _13995_/C VGND VGND VPWR VPWR _13996_/C sky130_fd_sc_hd__and3_4
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15734_ _12780_/X _23940_/Q VGND VGND VPWR VPWR _15734_/X sky130_fd_sc_hd__or2_4
X_18522_ _18565_/A _17423_/A VGND VGND VPWR VPWR _18522_/X sky130_fd_sc_hd__and2_4
X_12946_ _12962_/A _12946_/B _12946_/C VGND VGND VPWR VPWR _12947_/C sky130_fd_sc_hd__and3_4
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15665_ _12690_/A _23780_/Q VGND VGND VPWR VPWR _15665_/X sky130_fd_sc_hd__or2_4
X_18453_ _18399_/X VGND VGND VPWR VPWR _18453_/X sky130_fd_sc_hd__buf_2
X_12877_ _12877_/A _12877_/B _12877_/C VGND VGND VPWR VPWR _12877_/X sky130_fd_sc_hd__and3_4
X_17404_ _17401_/X _18557_/A VGND VGND VPWR VPWR _17404_/X sky130_fd_sc_hd__and2_4
X_14616_ _14616_/A VGND VGND VPWR VPWR _14676_/A sky130_fd_sc_hd__buf_2
X_18384_ _11633_/X _17188_/A _17848_/A VGND VGND VPWR VPWR _18384_/Y sky130_fd_sc_hd__a21oi_4
X_11828_ _11833_/A _11828_/B VGND VGND VPWR VPWR _11828_/X sky130_fd_sc_hd__or2_4
X_15596_ _15610_/A _24033_/Q VGND VGND VPWR VPWR _15596_/X sky130_fd_sc_hd__or2_4
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20547__A _20267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _22039_/A VGND VGND VPWR VPWR _21081_/A sky130_fd_sc_hd__inv_2
X_14547_ _15517_/A _14547_/B _14547_/C VGND VGND VPWR VPWR _14547_/X sky130_fd_sc_hd__and3_4
X_11759_ _16214_/A VGND VGND VPWR VPWR _11759_/X sky130_fd_sc_hd__buf_2
XANTENNA__22683__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14545__A _11681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20694__A1 _20635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20694__B2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17266_ _16819_/X VGND VGND VPWR VPWR _17266_/X sky130_fd_sc_hd__buf_2
X_14478_ _11914_/A _14476_/X _14477_/X VGND VGND VPWR VPWR _14478_/X sky130_fd_sc_hd__and3_4
XFILLER_105_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22762__A SYSTICKCLKDIV[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23409__CLK _23409_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16217_ _16163_/X _16215_/X _16216_/X VGND VGND VPWR VPWR _16221_/B sky130_fd_sc_hd__and3_4
X_19005_ _11537_/B VGND VGND VPWR VPWR _19005_/Y sky130_fd_sc_hd__inv_2
X_13429_ _12891_/A VGND VGND VPWR VPWR _13462_/A sky130_fd_sc_hd__buf_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17197_ _17197_/A VGND VGND VPWR VPWR _17197_/X sky130_fd_sc_hd__buf_2
XANTENNA__12065__A _12064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16148_ _16148_/A _16148_/B _16148_/C VGND VGND VPWR VPWR _16152_/B sky130_fd_sc_hd__and3_4
XANTENNA__17575__B _17251_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20282__A _20282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20997__A2 _20313_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15376__A _11752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16079_ _16079_/A _16000_/B VGND VGND VPWR VPWR _16081_/B sky130_fd_sc_hd__or2_4
XANTENNA__14280__A _14280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22199__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19907_ _20237_/A VGND VGND VPWR VPWR _19908_/A sky130_fd_sc_hd__inv_2
XFILLER_123_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19838_ _19553_/X _19837_/X _16922_/C _19553_/X VGND VGND VPWR VPWR _19838_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19769_ HRDATA[19] VGND VGND VPWR VPWR _20561_/B sky130_fd_sc_hd__buf_2
XFILLER_37_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13624__A _12504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21800_ _21592_/X _21798_/X _14754_/B _21795_/X VGND VGND VPWR VPWR _23641_/D sky130_fd_sc_hd__o22a_4
XFILLER_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16000__A _15967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22780_ _22780_/A _22781_/B _22793_/A VGND VGND VPWR VPWR _22780_/X sky130_fd_sc_hd__and3_4
XANTENNA__22371__A1 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21174__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22937__A _23079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22371__B2 _22366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21731_ _21724_/A VGND VGND VPWR VPWR _21731_/X sky130_fd_sc_hd__buf_2
XFILLER_25_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19949__C _18834_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24450_ _23475_/CLK _24450_/D HRESETn VGND VGND VPWR VPWR _20161_/A sky130_fd_sc_hd__dfrtp_4
X_21662_ _21658_/A VGND VGND VPWR VPWR _21677_/A sky130_fd_sc_hd__buf_2
X_23401_ _23561_/CLK _22245_/X VGND VGND VPWR VPWR _23401_/Q sky130_fd_sc_hd__dfxtp_4
X_20613_ _21560_/A VGND VGND VPWR VPWR _20613_/X sky130_fd_sc_hd__buf_2
XFILLER_162_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24363__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24381_ _24445_/CLK _24381_/D HRESETn VGND VGND VPWR VPWR _19090_/A sky130_fd_sc_hd__dfstp_4
XFILLER_71_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14455__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21593_ _21592_/X _21590_/X _14788_/B _21585_/X VGND VGND VPWR VPWR _23769_/D sky130_fd_sc_hd__o22a_4
XFILLER_32_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23332_ _23588_/CLK _23332_/D VGND VGND VPWR VPWR _15746_/B sky130_fd_sc_hd__dfxtp_4
X_20544_ _20447_/X _20541_/Y _20543_/X _19020_/Y _20495_/X VGND VGND VPWR VPWR _20545_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22672__A _22672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17550__A1 _16452_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24334__CLK _24294_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23263_ _23229_/CLK _22463_/X VGND VGND VPWR VPWR _23263_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20475_ _20269_/A VGND VGND VPWR VPWR _20475_/X sky130_fd_sc_hd__buf_2
XFILLER_152_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22214_ _22156_/X _22208_/X _14463_/B _22212_/X VGND VGND VPWR VPWR _22214_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21288__A _21264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23194_ _23194_/CLK _22580_/X VGND VGND VPWR VPWR _14560_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20192__A _20192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22145_ _22144_/X _22135_/X _14039_/B _22142_/X VGND VGND VPWR VPWR _23456_/D sky130_fd_sc_hd__o22a_4
XFILLER_134_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12703__A _13279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24484__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22076_ _21865_/X _22074_/X _13772_/B _22071_/X VGND VGND VPWR VPWR _22076_/X sky130_fd_sc_hd__o22a_4
XFILLER_126_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21027_ _22687_/A VGND VGND VPWR VPWR _21184_/A sky130_fd_sc_hd__buf_2
XANTENNA__18802__A1 _12678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23008__A _22912_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12800_ _12800_/A _23690_/Q VGND VGND VPWR VPWR _12800_/X sky130_fd_sc_hd__or2_4
X_13780_ _11813_/A _13764_/X _13779_/X VGND VGND VPWR VPWR _13781_/C sky130_fd_sc_hd__or3_4
X_22978_ _22912_/X VGND VGND VPWR VPWR _22978_/X sky130_fd_sc_hd__buf_2
XANTENNA__17369__A1 _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21165__A2 _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17369__B2 _17368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18566__B1 _17890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14349__B _14349_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12731_ _13301_/A _12731_/B VGND VGND VPWR VPWR _12731_/X sky130_fd_sc_hd__or2_4
XFILLER_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21929_ _21872_/X _21923_/X _14500_/B _21927_/X VGND VGND VPWR VPWR _23579_/D sky130_fd_sc_hd__o22a_4
XFILLER_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15450_ _15450_/A _15449_/X VGND VGND VPWR VPWR _15450_/X sky130_fd_sc_hd__and2_4
X_12662_ _12632_/A _12565_/B VGND VGND VPWR VPWR _12662_/X sky130_fd_sc_hd__or2_4
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22114__A1 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_101_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR _24096_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22114__B2 _22106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14401_ _13752_/A _14399_/X _14400_/X VGND VGND VPWR VPWR _14401_/X sky130_fd_sc_hd__and3_4
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11610_/X _18888_/B VGND VGND VPWR VPWR _20095_/D sky130_fd_sc_hd__or2_4
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15381_/A VGND VGND VPWR VPWR _15382_/B sky130_fd_sc_hd__buf_2
XANTENNA__18869__A1 _15651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12971_/A _23755_/Q VGND VGND VPWR VPWR _12593_/X sky130_fd_sc_hd__or2_4
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ _16523_/B VGND VGND VPWR VPWR _17120_/Y sky130_fd_sc_hd__inv_2
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _15450_/A _14332_/B VGND VGND VPWR VPWR _14332_/X sky130_fd_sc_hd__and2_4
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ _24370_/Q _18964_/A _11544_/C _11544_/D VGND VGND VPWR VPWR _11544_/X sky130_fd_sc_hd__or4_4
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17051_ _17050_/X VGND VGND VPWR VPWR _17051_/X sky130_fd_sc_hd__buf_2
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _14263_/A _14263_/B VGND VGND VPWR VPWR _14263_/X sky130_fd_sc_hd__or2_4
XFILLER_156_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22417__A2 _22414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16002_ _16110_/A _16000_/X _16001_/X VGND VGND VPWR VPWR _16003_/C sky130_fd_sc_hd__and3_4
XFILLER_104_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21625__B1 _23755_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13214_ _13232_/A _13212_/X _13214_/C VGND VGND VPWR VPWR _13214_/X sky130_fd_sc_hd__and3_4
XANTENNA__23701__CLK _23456_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21198__A _21198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14194_ _15324_/A VGND VGND VPWR VPWR _14631_/A sky130_fd_sc_hd__buf_2
XFILLER_48_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13145_ _13145_/A _24007_/Q VGND VGND VPWR VPWR _13146_/C sky130_fd_sc_hd__or2_4
XANTENNA__13709__A _12634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12613__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13076_ _13096_/A _13076_/B _13076_/C VGND VGND VPWR VPWR _13083_/B sky130_fd_sc_hd__and3_4
X_17953_ _18413_/A VGND VGND VPWR VPWR _18411_/A sky130_fd_sc_hd__buf_2
XFILLER_151_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21928__A1 _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21928__B2 _21927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19597__A2 _19724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16904_ _12025_/B _12183_/X VGND VGND VPWR VPWR _16904_/Y sky130_fd_sc_hd__nor2_4
X_12027_ _11858_/X VGND VGND VPWR VPWR _12027_/X sky130_fd_sc_hd__buf_2
XFILLER_66_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17884_ _17875_/X _17881_/X _17883_/X VGND VGND VPWR VPWR _17885_/B sky130_fd_sc_hd__o21ai_4
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19623_ _19623_/A VGND VGND VPWR VPWR _19834_/A sky130_fd_sc_hd__buf_2
X_16835_ _12423_/X _16834_/X _12423_/X _16834_/X VGND VGND VPWR VPWR _16897_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13444__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24207__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19554_ _19515_/X _19551_/X _18782_/B _19553_/X VGND VGND VPWR VPWR _19554_/X sky130_fd_sc_hd__a2bb2o_4
X_16766_ _16757_/X _16766_/B VGND VGND VPWR VPWR _16766_/X sky130_fd_sc_hd__or2_4
XFILLER_53_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13978_ _12501_/A _14039_/B VGND VGND VPWR VPWR _13979_/C sky130_fd_sc_hd__or2_4
XANTENNA__21156__A2 _21155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18505_ _17648_/X VGND VGND VPWR VPWR _18506_/A sky130_fd_sc_hd__buf_2
XFILLER_59_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12929_ _12941_/A _12929_/B _12929_/C VGND VGND VPWR VPWR _12930_/C sky130_fd_sc_hd__and3_4
X_15717_ _11856_/A _11630_/A _15686_/X _12264_/X _15716_/X VGND VGND VPWR VPWR _15717_/X
+ sky130_fd_sc_hd__a32o_4
X_19485_ _19480_/X _19483_/X HRDATA[12] _19484_/X VGND VGND VPWR VPWR _19823_/A sky130_fd_sc_hd__o22a_4
X_16697_ _16586_/A _16761_/B VGND VGND VPWR VPWR _16699_/B sky130_fd_sc_hd__or2_4
XANTENNA__16755__A _11768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18436_ _18435_/X VGND VGND VPWR VPWR _18436_/Y sky130_fd_sc_hd__inv_2
X_15648_ _13894_/A _15640_/X _15647_/X VGND VGND VPWR VPWR _15649_/C sky130_fd_sc_hd__and3_4
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24357__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11899__A _14421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22656__A2 _22651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18367_ _18367_/A _18366_/X VGND VGND VPWR VPWR _18368_/B sky130_fd_sc_hd__or2_4
X_15579_ _15449_/A _15575_/X _15579_/C VGND VGND VPWR VPWR _15579_/X sky130_fd_sc_hd__or3_4
XANTENNA__14275__A _14280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17318_ _17318_/A VGND VGND VPWR VPWR _17630_/A sky130_fd_sc_hd__inv_2
XANTENNA__21864__B1 _23615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18298_ _17517_/Y _18296_/X _18176_/X VGND VGND VPWR VPWR _18298_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12507__B _12632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17586__A _17140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17249_ _18538_/A VGND VGND VPWR VPWR _17249_/X sky130_fd_sc_hd__buf_2
XFILLER_128_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23381__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20260_ _20260_/A VGND VGND VPWR VPWR _20260_/X sky130_fd_sc_hd__buf_2
XFILLER_115_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13619__A _15423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21092__B2 _21087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20191_ _20156_/Y _20191_/B VGND VGND VPWR VPWR _20191_/X sky130_fd_sc_hd__and2_4
XANTENNA__12523__A _12881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21836__A _20531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21919__B2 _21913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23950_ _23918_/CLK _23950_/D VGND VGND VPWR VPWR _16038_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22901_ _19915_/X _22843_/X _15785_/A _20665_/X VGND VGND VPWR VPWR _22901_/X sky130_fd_sc_hd__o22a_4
XFILLER_69_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22592__B2 _22591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23881_ _24073_/CLK _23881_/D VGND VGND VPWR VPWR _23881_/Q sky130_fd_sc_hd__dfxtp_4
X_22832_ _22819_/X _14767_/Y VGND VGND VPWR VPWR _22832_/X sky130_fd_sc_hd__or2_4
XFILLER_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21147__A2 _21141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14169__B _23711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18548__B1 _18543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22763_ _22763_/A VGND VGND VPWR VPWR _22763_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21714_ _21528_/X _21713_/X _23699_/Q _21710_/X VGND VGND VPWR VPWR _21714_/X sky130_fd_sc_hd__o22a_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22694_ _22708_/A VGND VGND VPWR VPWR _22694_/X sky130_fd_sc_hd__buf_2
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24433_ _23379_/CLK _18847_/X HRESETn VGND VGND VPWR VPWR _24433_/Q sky130_fd_sc_hd__dfrtp_4
X_21645_ _21624_/A VGND VGND VPWR VPWR _21645_/X sky130_fd_sc_hd__buf_2
XFILLER_123_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24340__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14185__A _14616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22647__A2 _22644_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24364_ _24360_/CLK _24364_/D HRESETn VGND VGND VPWR VPWR _11538_/A sky130_fd_sc_hd__dfstp_4
XFILLER_166_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21576_ _21575_/X _21566_/X _23776_/Q _21573_/X VGND VGND VPWR VPWR _21576_/X sky130_fd_sc_hd__o22a_4
XFILLER_165_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23315_ _23379_/CLK _23315_/D VGND VGND VPWR VPWR _12128_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_138_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20527_ _20466_/X _20513_/Y _20525_/X _20526_/Y _20481_/X VGND VGND VPWR VPWR _20527_/X
+ sky130_fd_sc_hd__a32o_4
X_24295_ _24357_/CLK _19284_/X HRESETn VGND VGND VPWR VPWR _24295_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23246_ _23246_/CLK _23246_/D VGND VGND VPWR VPWR _16000_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20458_ _20457_/X VGND VGND VPWR VPWR _20458_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14632__B _14560_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13529__A _13529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23177_ _23337_/CLK _22609_/X VGND VGND VPWR VPWR _12935_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20389_ _18011_/X _20260_/X _20341_/X _20388_/Y VGND VGND VPWR VPWR _20389_/X sky130_fd_sc_hd__a211o_4
XFILLER_134_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22128_ _22127_/X _22123_/X _13217_/B _22118_/X VGND VGND VPWR VPWR _23463_/D sky130_fd_sc_hd__o22a_4
XFILLER_47_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_26_0_HCLK clkbuf_6_13_0_HCLK/X VGND VGND VPWR VPWR _24360_/CLK sky130_fd_sc_hd__clkbuf_1
X_14950_ _11673_/A _14932_/X _14949_/X VGND VGND VPWR VPWR _14950_/X sky130_fd_sc_hd__or3_4
XFILLER_48_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22059_ _21836_/X _22053_/X _12833_/B _22057_/X VGND VGND VPWR VPWR _22059_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_89_0_HCLK clkbuf_7_89_0_HCLK/A VGND VGND VPWR VPWR _23294_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_88_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21386__A2 _21384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22583__B2 _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13901_ _13706_/A _13901_/B VGND VGND VPWR VPWR _13901_/X sky130_fd_sc_hd__or2_4
XANTENNA__15463__B _23778_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14881_ _14881_/A _23958_/Q VGND VGND VPWR VPWR _14881_/X sky130_fd_sc_hd__or2_4
XANTENNA__21184__C _21184_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13264__A _13192_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16620_ _11760_/X VGND VGND VPWR VPWR _16682_/A sky130_fd_sc_hd__buf_2
X_13832_ _15423_/A _23965_/Q VGND VGND VPWR VPWR _13833_/C sky130_fd_sc_hd__or2_4
XFILLER_75_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24499__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14079__B _23648_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16551_ _11891_/X VGND VGND VPWR VPWR _16593_/A sky130_fd_sc_hd__buf_2
X_13763_ _14372_/A _13759_/X _13763_/C VGND VGND VPWR VPWR _13763_/X sky130_fd_sc_hd__or3_4
XANTENNA__16014__A1 _16130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17211__B1 _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15502_ _15502_/A _15502_/B VGND VGND VPWR VPWR _15502_/X sky130_fd_sc_hd__or2_4
X_12714_ _12745_/A _12714_/B _12713_/X VGND VGND VPWR VPWR _12714_/X sky130_fd_sc_hd__and3_4
XFILLER_71_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16482_ _16481_/X _16406_/B VGND VGND VPWR VPWR _16482_/X sky130_fd_sc_hd__or2_4
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19270_ _24302_/Q _19251_/B _19269_/Y VGND VGND VPWR VPWR _24302_/D sky130_fd_sc_hd__o21a_4
X_13694_ _13694_/A VGND VGND VPWR VPWR _13695_/A sky130_fd_sc_hd__buf_2
XFILLER_70_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20097__A NMI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15433_ _12198_/A _15497_/B VGND VGND VPWR VPWR _15434_/C sky130_fd_sc_hd__or2_4
X_18221_ _18405_/A _18165_/B VGND VGND VPWR VPWR _18221_/X sky130_fd_sc_hd__or2_4
X_12645_ _12972_/A _12643_/X _12645_/C VGND VGND VPWR VPWR _12645_/X sky130_fd_sc_hd__and3_4
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14095__A _12473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15364_ _15328_/A _15305_/B VGND VGND VPWR VPWR _15364_/X sky130_fd_sc_hd__or2_4
X_18152_ _18407_/A _17478_/B VGND VGND VPWR VPWR _18155_/C sky130_fd_sc_hd__nor2_4
X_12576_ _12576_/A VGND VGND VPWR VPWR _12977_/A sky130_fd_sc_hd__buf_2
XFILLER_157_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21310__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17103_ _17103_/A _18440_/A VGND VGND VPWR VPWR _17104_/D sky130_fd_sc_hd__and2_4
X_14315_ _13656_/A _14392_/B VGND VGND VPWR VPWR _14316_/C sky130_fd_sc_hd__or2_4
XFILLER_7_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _19063_/A _11526_/X VGND VGND VPWR VPWR _11528_/B sky130_fd_sc_hd__or2_4
X_18083_ _18083_/A VGND VGND VPWR VPWR _18083_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15295_ _14272_/A _15293_/X _15294_/X VGND VGND VPWR VPWR _15295_/X sky130_fd_sc_hd__and3_4
XFILLER_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17034_ _17481_/B VGND VGND VPWR VPWR _17035_/A sky130_fd_sc_hd__buf_2
XFILLER_156_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14246_ _14201_/A _14244_/X _14245_/X VGND VGND VPWR VPWR _14246_/X sky130_fd_sc_hd__and3_4
XANTENNA__13439__A _12873_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21074__B2 _21070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14177_ _15321_/A VGND VGND VPWR VPWR _14615_/A sky130_fd_sc_hd__buf_2
XANTENNA__12343__A _11689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13128_ _12690_/A _23527_/Q VGND VGND VPWR VPWR _13129_/C sky130_fd_sc_hd__or2_4
X_18985_ _18978_/X _18984_/X _18978_/X _24367_/Q VGND VGND VPWR VPWR _24367_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15654__A _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13059_ _13094_/A _12991_/B VGND VGND VPWR VPWR _13059_/X sky130_fd_sc_hd__or2_4
X_17936_ _17824_/X _17932_/Y _17933_/X _17935_/Y VGND VGND VPWR VPWR _17936_/X sky130_fd_sc_hd__o22a_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22574__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17867_ _17867_/A VGND VGND VPWR VPWR _18711_/B sky130_fd_sc_hd__inv_2
XFILLER_39_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13174__A _13338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19606_ _19510_/X _19601_/X _19603_/X _19605_/X VGND VGND VPWR VPWR _19606_/X sky130_fd_sc_hd__a211o_4
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16818_ _16684_/A _16818_/B _16818_/C VGND VGND VPWR VPWR _16818_/X sky130_fd_sc_hd__or3_4
XFILLER_4_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21129__A2 _21125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17798_ _17798_/A VGND VGND VPWR VPWR _18335_/A sky130_fd_sc_hd__buf_2
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21391__A _21391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19537_ _19623_/A _19537_/B VGND VGND VPWR VPWR _19538_/A sky130_fd_sc_hd__or2_4
XFILLER_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16749_ _11984_/X _16726_/X _16733_/X _16740_/X _16748_/X VGND VGND VPWR VPWR _16749_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13902__A _13697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19468_ _19439_/A VGND VGND VPWR VPWR _19700_/A sky130_fd_sc_hd__buf_2
XANTENNA__14717__B _14717_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18419_ _18418_/Y _17437_/B _17443_/X VGND VGND VPWR VPWR _18419_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12518__A _12487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19399_ _19428_/A VGND VGND VPWR VPWR _19399_/X sky130_fd_sc_hd__buf_2
XFILLER_33_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21430_ _21249_/X _21427_/X _23857_/Q _21424_/X VGND VGND VPWR VPWR _23857_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21301__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15829__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21361_ _21302_/X _21355_/X _14452_/B _21359_/X VGND VGND VPWR VPWR _23899_/D sky130_fd_sc_hd__o22a_4
X_23100_ _23515_/CLK _22727_/X VGND VGND VPWR VPWR _14396_/B sky130_fd_sc_hd__dfxtp_4
X_20312_ _20233_/Y VGND VGND VPWR VPWR _20638_/A sky130_fd_sc_hd__buf_2
X_24080_ _24080_/CLK _21043_/X VGND VGND VPWR VPWR _16425_/B sky130_fd_sc_hd__dfxtp_4
X_21292_ _20801_/A VGND VGND VPWR VPWR _21292_/X sky130_fd_sc_hd__buf_2
XANTENNA__14452__B _14452_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22950__A _18590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13349__A _13349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23031_ _22910_/X VGND VGND VPWR VPWR _23055_/B sky130_fd_sc_hd__buf_2
XANTENNA__21065__B2 _21063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20243_ _20864_/A _20238_/X _20239_/X _20240_/X _20242_/X VGND VGND VPWR VPWR _20244_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21566__A _21542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20174_ _20163_/Y _20164_/Y _11567_/X _20173_/X VGND VGND VPWR VPWR _20174_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15564__A _14431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21368__A2 _21341_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23933_ _23582_/CLK _23933_/D VGND VGND VPWR VPWR _13896_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23864_ _23864_/CLK _23864_/D VGND VGND VPWR VPWR _23864_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22317__B2 _22312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22397__A _22357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22815_ _22801_/X VGND VGND VPWR VPWR _22815_/X sky130_fd_sc_hd__buf_2
XFILLER_26_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16395__A _16009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23795_ _23760_/CLK _21531_/X VGND VGND VPWR VPWR _23795_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14908__A _11928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13812__A _12470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22746_ _19519_/X _22745_/Y HREADY VGND VGND VPWR VPWR _22746_/X sky130_fd_sc_hd__o21a_4
XFILLER_41_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21540__A2 _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22677_ _22468_/X _22672_/X _14387_/B _22676_/X VGND VGND VPWR VPWR _22677_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12428__A _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12430_ _13792_/A VGND VGND VPWR VPWR _14905_/A sky130_fd_sc_hd__buf_2
X_24416_ _23476_/CLK _18872_/X HRESETn VGND VGND VPWR VPWR _24416_/Q sky130_fd_sc_hd__dfrtp_4
X_21628_ _21553_/X _21627_/X _12919_/B _21624_/X VGND VGND VPWR VPWR _23753_/D sky130_fd_sc_hd__o22a_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23021__A _18272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12361_ _12407_/A _12361_/B VGND VGND VPWR VPWR _12365_/B sky130_fd_sc_hd__or2_4
XANTENNA__15739__A _11701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24347_ _24382_/CLK _24347_/D HRESETn VGND VGND VPWR VPWR _11521_/A sky130_fd_sc_hd__dfstp_4
X_21559_ _21558_/X _21554_/X _23783_/Q _21549_/X VGND VGND VPWR VPWR _23783_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18115__A _18485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14643__A _13882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20364__B _20364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14100_ _11869_/A _14100_/B _14099_/X VGND VGND VPWR VPWR _14100_/X sky130_fd_sc_hd__or3_4
XFILLER_165_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15080_ _15080_/A _23541_/Q VGND VGND VPWR VPWR _15081_/C sky130_fd_sc_hd__or2_4
XFILLER_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15458__B _15458_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12292_ _13183_/A VGND VGND VPWR VPWR _12735_/A sky130_fd_sc_hd__buf_2
X_24278_ _24292_/CLK _19318_/X HRESETn VGND VGND VPWR VPWR _24278_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14362__B _14362_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14031_ _14056_/A _23296_/Q VGND VGND VPWR VPWR _14031_/X sky130_fd_sc_hd__or2_4
XANTENNA__13259__A _11682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23229_ _23229_/CLK _22525_/X VGND VGND VPWR VPWR _13848_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15474__A _12626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18770_ _17100_/A _19963_/B _17100_/A _19963_/B VGND VGND VPWR VPWR _18770_/X sky130_fd_sc_hd__a2bb2o_4
X_15982_ _15982_/A _23982_/Q VGND VGND VPWR VPWR _15983_/C sky130_fd_sc_hd__or2_4
XANTENNA__22556__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17721_ _17721_/A VGND VGND VPWR VPWR _18533_/A sky130_fd_sc_hd__buf_2
X_14933_ _14922_/A _14871_/B VGND VGND VPWR VPWR _14933_/X sky130_fd_sc_hd__or2_4
XANTENNA__15193__B _15129_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17652_ _16932_/X VGND VGND VPWR VPWR _17652_/X sky130_fd_sc_hd__buf_2
X_14864_ _14127_/A _14864_/B VGND VGND VPWR VPWR _14864_/X sky130_fd_sc_hd__or2_4
XFILLER_75_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16603_ _16602_/X VGND VGND VPWR VPWR _16687_/A sky130_fd_sc_hd__inv_2
XFILLER_169_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13815_ _12503_/A VGND VGND VPWR VPWR _14319_/A sky130_fd_sc_hd__buf_2
XFILLER_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17583_ _17583_/A _17583_/B _18099_/A _18138_/A VGND VGND VPWR VPWR _17583_/X sky130_fd_sc_hd__or4_4
X_14795_ _14674_/A _14727_/B VGND VGND VPWR VPWR _14795_/X sky130_fd_sc_hd__or2_4
XFILLER_95_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19322_ _23086_/B _19226_/B _19321_/Y VGND VGND VPWR VPWR _24277_/D sky130_fd_sc_hd__o21a_4
XFILLER_73_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13746_ _12635_/A _13744_/X _13745_/X VGND VGND VPWR VPWR _13747_/C sky130_fd_sc_hd__and3_4
X_16534_ _11960_/A VGND VGND VPWR VPWR _16534_/X sky130_fd_sc_hd__buf_2
XFILLER_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21531__A2 _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19253_ _19253_/A _19253_/B VGND VGND VPWR VPWR _19254_/B sky130_fd_sc_hd__and2_4
X_16465_ _16465_/A _16463_/X _16464_/X VGND VGND VPWR VPWR _16470_/B sky130_fd_sc_hd__and3_4
X_13677_ _13677_/A _13677_/B _13677_/C VGND VGND VPWR VPWR _13681_/B sky130_fd_sc_hd__and3_4
XANTENNA__12338__A _12401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18204_ _18320_/A _18203_/Y VGND VGND VPWR VPWR _18204_/X sky130_fd_sc_hd__and2_4
X_12628_ _12975_/A _12624_/X _12628_/C VGND VGND VPWR VPWR _12629_/C sky130_fd_sc_hd__and3_4
X_15416_ _13628_/A _15473_/B VGND VGND VPWR VPWR _15416_/X sky130_fd_sc_hd__or2_4
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16396_ _16011_/A _16394_/X _16395_/X VGND VGND VPWR VPWR _16396_/X sky130_fd_sc_hd__and3_4
X_19184_ _24329_/Q _19185_/A _19183_/Y VGND VGND VPWR VPWR _19184_/X sky130_fd_sc_hd__o21a_4
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15347_ _11673_/A _15347_/B _15346_/X VGND VGND VPWR VPWR _15347_/X sky130_fd_sc_hd__or3_4
X_18135_ _18168_/A _18134_/X VGND VGND VPWR VPWR _18135_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15649__A _15649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12559_ _12559_/A _12671_/B VGND VGND VPWR VPWR _12559_/X sky130_fd_sc_hd__or2_4
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14553__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18066_ _17664_/Y _18014_/X _17664_/Y _18014_/X VGND VGND VPWR VPWR _18066_/X sky130_fd_sc_hd__a2bb2o_4
X_15278_ _14994_/A _23448_/Q VGND VGND VPWR VPWR _15278_/X sky130_fd_sc_hd__or2_4
XANTENNA__21047__B2 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13169__A _13301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17017_ _17017_/A _17017_/B VGND VGND VPWR VPWR _17025_/A sky130_fd_sc_hd__or2_4
X_14229_ _14229_/A VGND VGND VPWR VPWR _14623_/A sky130_fd_sc_hd__buf_2
XANTENNA__12073__A _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12801__A _12801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18968_ _19021_/A VGND VGND VPWR VPWR _18968_/X sky130_fd_sc_hd__buf_2
XFILLER_140_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22547__B2 _22541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17919_ _18168_/A VGND VGND VPWR VPWR _17919_/X sky130_fd_sc_hd__buf_2
XFILLER_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12520__B _12520_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18899_ _18928_/A VGND VGND VPWR VPWR _18900_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_72_0_HCLK clkbuf_7_72_0_HCLK/A VGND VGND VPWR VPWR _23904_/CLK sky130_fd_sc_hd__clkbuf_1
X_20930_ _20930_/A _20929_/X VGND VGND VPWR VPWR _20930_/Y sky130_fd_sc_hd__nor2_4
XFILLER_54_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20861_ _20510_/A VGND VGND VPWR VPWR _20861_/X sky130_fd_sc_hd__buf_2
XANTENNA__22010__A _22010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14728__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22600_ _22423_/X _22594_/X _16273_/B _22598_/X VGND VGND VPWR VPWR _22600_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13632__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23580_ _23515_/CLK _23580_/D VGND VGND VPWR VPWR _14360_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20792_ _20781_/X _20790_/X _24319_/Q _20791_/X VGND VGND VPWR VPWR _20792_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22945__A _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22531_ _22476_/X _22529_/X _14753_/B _22526_/X VGND VGND VPWR VPWR _22531_/X sky130_fd_sc_hd__o22a_4
XFILLER_23_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22462_ _22462_/A VGND VGND VPWR VPWR _22462_/X sky130_fd_sc_hd__buf_2
X_24201_ _23671_/CLK _19739_/X HRESETn VGND VGND VPWR VPWR _12466_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20089__A2 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21413_ _21304_/X _21412_/X _14688_/B _21409_/X VGND VGND VPWR VPWR _21413_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21286__B2 _21276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15559__A _11886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14463__A _13010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22393_ _22151_/X _22390_/X _13811_/B _22387_/X VGND VGND VPWR VPWR _23293_/D sky130_fd_sc_hd__o22a_4
XFILLER_163_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24132_ _24137_/CLK _20205_/Y HRESETn VGND VGND VPWR VPWR _18576_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21344_ _21273_/X _21341_/X _13161_/B _21338_/X VGND VGND VPWR VPWR _21344_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16162__B1 _11608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24063_ _23997_/CLK _24063_/D VGND VGND VPWR VPWR _24063_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21275_ _21560_/A VGND VGND VPWR VPWR _21275_/X sky130_fd_sc_hd__buf_2
XFILLER_150_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23014_ _22949_/A _23014_/B VGND VGND VPWR VPWR _23016_/B sky130_fd_sc_hd__or2_4
X_20226_ _16937_/X VGND VGND VPWR VPWR _20226_/X sky130_fd_sc_hd__buf_2
XFILLER_131_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20157_ _20157_/A VGND VGND VPWR VPWR _20157_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12711__A _12279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23912__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19403__A1 _19399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20088_ _20088_/A VGND VGND VPWR VPWR _20088_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21210__B2 _21209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11930_ _11930_/A VGND VGND VPWR VPWR _11931_/A sky130_fd_sc_hd__buf_2
XFILLER_85_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23916_ _23500_/CLK _23916_/D VGND VGND VPWR VPWR _12268_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23847_ _23111_/CLK _23847_/D VGND VGND VPWR VPWR _23847_/Q sky130_fd_sc_hd__dfxtp_4
X_11861_ _13586_/A VGND VGND VPWR VPWR _13689_/A sky130_fd_sc_hd__buf_2
XFILLER_166_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _14296_/A VGND VGND VPWR VPWR _13601_/A sky130_fd_sc_hd__buf_2
XPHY_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13542__A _13542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14301_/A _14580_/B _14579_/X VGND VGND VPWR VPWR _14580_/X sky130_fd_sc_hd__or3_4
XPHY_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23778_ _23650_/CLK _23778_/D VGND VGND VPWR VPWR _23778_/Q sky130_fd_sc_hd__dfxtp_4
X_11792_ _11768_/X VGND VGND VPWR VPWR _11792_/X sky130_fd_sc_hd__buf_2
XPHY_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17717__B2 _17360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _13531_/A _23909_/Q VGND VGND VPWR VPWR _13533_/B sky130_fd_sc_hd__or2_4
XANTENNA__22710__B2 _22705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22729_ _22722_/A VGND VGND VPWR VPWR _22729_/X sky130_fd_sc_hd__buf_2
X_16250_ _16096_/A VGND VGND VPWR VPWR _16282_/A sky130_fd_sc_hd__buf_2
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13462_ _13462_/A _13462_/B VGND VGND VPWR VPWR _13464_/B sky130_fd_sc_hd__or2_4
XFILLER_16_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20375__A _20358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15201_ _14783_/X _15201_/B _15200_/X VGND VGND VPWR VPWR _15201_/X sky130_fd_sc_hd__or3_4
XFILLER_51_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12413_ _15851_/A _23660_/Q VGND VGND VPWR VPWR _12413_/X sky130_fd_sc_hd__or2_4
X_16181_ _13378_/A VGND VGND VPWR VPWR _16181_/X sky130_fd_sc_hd__buf_2
XANTENNA__21277__B2 _21276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15469__A _12576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13393_ _13384_/A _13316_/B VGND VGND VPWR VPWR _13393_/X sky130_fd_sc_hd__or2_4
XANTENNA__14373__A _12616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15132_ _14897_/X VGND VGND VPWR VPWR _15269_/A sky130_fd_sc_hd__buf_2
X_12344_ _12827_/A _12344_/B VGND VGND VPWR VPWR _12346_/B sky130_fd_sc_hd__or2_4
XANTENNA__23442__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19940_ _19938_/X _24169_/Q _19939_/X _20512_/B VGND VGND VPWR VPWR _24169_/D sky130_fd_sc_hd__o22a_4
X_15063_ _15086_/A _23285_/Q VGND VGND VPWR VPWR _15063_/X sky130_fd_sc_hd__or2_4
XFILLER_154_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12275_ _12726_/A _12275_/B _12274_/X VGND VGND VPWR VPWR _12275_/X sky130_fd_sc_hd__or3_4
XFILLER_99_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14014_ _13951_/X _11625_/X _13982_/X _11603_/A _14013_/X VGND VGND VPWR VPWR _14014_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19871_ _19700_/A _19867_/X _19870_/Y _21081_/A _19552_/X VGND VGND VPWR VPWR _19871_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20252__A2 _20246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18822_ _13945_/X _18817_/X _24445_/Q _18818_/X VGND VGND VPWR VPWR _24445_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23592__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12621__A _12604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18753_ _18753_/A VGND VGND VPWR VPWR _18753_/Y sky130_fd_sc_hd__inv_2
X_15965_ _15961_/A _15965_/B _15965_/C VGND VGND VPWR VPWR _15971_/B sky130_fd_sc_hd__and3_4
XANTENNA__24443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_59_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14482__A3 _14451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17704_ _17703_/X VGND VGND VPWR VPWR _17704_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20004__A2 _19983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21201__B2 _21195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14916_ _13717_/A VGND VGND VPWR VPWR _14916_/X sky130_fd_sc_hd__buf_2
X_18684_ _18064_/X _18671_/X _18019_/X _18683_/X VGND VGND VPWR VPWR _18684_/X sky130_fd_sc_hd__o22a_4
XFILLER_64_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15896_ _15903_/A _15840_/B VGND VGND VPWR VPWR _15896_/X sky130_fd_sc_hd__or2_4
XANTENNA__13690__A1 _11969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21752__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17635_ _17635_/A _17635_/B _17617_/Y _17635_/D VGND VGND VPWR VPWR _17636_/B sky130_fd_sc_hd__or4_4
XFILLER_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14847_ _14767_/Y _14844_/X _15387_/B VGND VGND VPWR VPWR _14847_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14548__A _14547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13452__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17566_ _11611_/C _17035_/A VGND VGND VPWR VPWR _17566_/X sky130_fd_sc_hd__and2_4
X_14778_ _15112_/A _14774_/X _14778_/C VGND VGND VPWR VPWR _14778_/X sky130_fd_sc_hd__and3_4
XANTENNA__22765__A SYSTICKCLKDIV[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21504__A2 _21499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19305_ _19234_/B VGND VGND VPWR VPWR _19305_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16517_ _16163_/X _16517_/B _16517_/C VGND VGND VPWR VPWR _16518_/C sky130_fd_sc_hd__and3_4
X_13729_ _13743_/A _13729_/B _13728_/X VGND VGND VPWR VPWR _13730_/C sky130_fd_sc_hd__and3_4
XANTENNA__16763__A _16647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17497_ _13583_/X _17530_/B VGND VGND VPWR VPWR _17497_/X sky130_fd_sc_hd__and2_4
XANTENNA__12068__A _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19236_ _24287_/Q _19236_/B VGND VGND VPWR VPWR _19237_/B sky130_fd_sc_hd__and2_4
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16448_ _13468_/A _16444_/X _16448_/C VGND VGND VPWR VPWR _16448_/X sky130_fd_sc_hd__or3_4
XFILLER_108_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15379__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19167_ _19159_/B VGND VGND VPWR VPWR _19167_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22465__B1 _13702_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16379_ _13416_/A _16361_/X _16378_/X VGND VGND VPWR VPWR _16379_/X sky130_fd_sc_hd__or3_4
XANTENNA__14283__A _14448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18118_ _18378_/A _18118_/B VGND VGND VPWR VPWR _18119_/D sky130_fd_sc_hd__and2_4
X_19098_ _11521_/A VGND VGND VPWR VPWR _19098_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22217__B1 _23417_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18049_ _17849_/A _17879_/X _17227_/X _18048_/X VGND VGND VPWR VPWR _18049_/X sky130_fd_sc_hd__o22a_4
XFILLER_144_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21060_ _20659_/X _21059_/X _15756_/B _21056_/X VGND VGND VPWR VPWR _21060_/X sky130_fd_sc_hd__o22a_4
XFILLER_154_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15826__B _15826_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20011_ _20010_/X VGND VGND VPWR VPWR _20011_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21440__B2 _21438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12531__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19397__B1 _19396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21962_ _21841_/X _21960_/X _13006_/B _21957_/X VGND VGND VPWR VPWR _23560_/D sky130_fd_sc_hd__o22a_4
XFILLER_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21743__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23701_ _23456_/CLK _23701_/D VGND VGND VPWR VPWR _23701_/Q sky130_fd_sc_hd__dfxtp_4
X_20913_ _24218_/Q _20895_/X _20912_/Y VGND VGND VPWR VPWR _22158_/A sky130_fd_sc_hd__o21a_4
X_21893_ _21887_/Y _21892_/X _21811_/X _21892_/X VGND VGND VPWR VPWR _23604_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14458__A _12461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13362__A _13392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23632_ _23533_/CLK _23632_/D VGND VGND VPWR VPWR _16424_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_82_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20844_ _20844_/A _20844_/B VGND VGND VPWR VPWR _20844_/X sky130_fd_sc_hd__or2_4
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_2_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR _24382_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23563_ _24074_/CLK _21958_/X VGND VGND VPWR VPWR _12514_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20775_ HRDATA[10] _20668_/A VGND VGND VPWR VPWR _20777_/B sky130_fd_sc_hd__or2_4
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19687__C _19687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22514_ _22447_/X _22508_/X _23237_/Q _22512_/X VGND VGND VPWR VPWR _22514_/X sky130_fd_sc_hd__o22a_4
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23494_ _24102_/CLK _22065_/X VGND VGND VPWR VPWR _23494_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22445_ _22433_/A VGND VGND VPWR VPWR _22445_/X sky130_fd_sc_hd__buf_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15289__A _14277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12706__A _13145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11610__A _11609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22376_ _22376_/A VGND VGND VPWR VPWR _22376_/X sky130_fd_sc_hd__buf_2
X_24115_ _23764_/CLK _24115_/D VGND VGND VPWR VPWR _24115_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21327_ _21341_/A VGND VGND VPWR VPWR _21327_/X sky130_fd_sc_hd__buf_2
XANTENNA__20482__A2 _20468_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14921__A _15369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24046_ _23438_/CLK _21098_/X VGND VGND VPWR VPWR _24046_/Q sky130_fd_sc_hd__dfxtp_4
X_12060_ _12059_/X _24019_/Q VGND VGND VPWR VPWR _12061_/C sky130_fd_sc_hd__or2_4
X_21258_ _21256_/X _21257_/X _16038_/B _21252_/X VGND VGND VPWR VPWR _23950_/D sky130_fd_sc_hd__o22a_4
XFILLER_89_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20234__A2 _18779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20209_ _20208_/X VGND VGND VPWR VPWR _20209_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21189_ _21183_/Y _21188_/X _20299_/X _21188_/X VGND VGND VPWR VPWR _21189_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21982__A2 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15752__A _12758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12962_ _12962_/A _12962_/B _12961_/X VGND VGND VPWR VPWR _12978_/B sky130_fd_sc_hd__and3_4
X_15750_ _13092_/A _15740_/X _15750_/C VGND VGND VPWR VPWR _15750_/X sky130_fd_sc_hd__and3_4
XFILLER_18_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11913_ _11913_/A VGND VGND VPWR VPWR _11914_/A sky130_fd_sc_hd__buf_2
X_14701_ _14700_/X VGND VGND VPWR VPWR _14701_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15471__B _15471_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12893_ _12889_/A _12891_/X _12892_/X VGND VGND VPWR VPWR _12893_/X sky130_fd_sc_hd__and3_4
X_15681_ _12240_/A _15737_/B VGND VGND VPWR VPWR _15681_/X sky130_fd_sc_hd__or2_4
XANTENNA__20942__B1 HRDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17420_ _17161_/X _17421_/B VGND VGND VPWR VPWR _17423_/A sky130_fd_sc_hd__and2_4
X_11844_ _12168_/A _11844_/B _11844_/C VGND VGND VPWR VPWR _11848_/B sky130_fd_sc_hd__and3_4
XFILLER_33_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14632_ _14819_/A _14560_/B VGND VGND VPWR VPWR _14632_/X sky130_fd_sc_hd__or2_4
XFILLER_61_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18782__B _18782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17310_/X _17351_/B _17301_/A _18600_/A VGND VGND VPWR VPWR _17351_/X sky130_fd_sc_hd__and4_4
X_14563_ _14304_/A _14563_/B VGND VGND VPWR VPWR _14565_/B sky130_fd_sc_hd__or2_4
XPHY_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21498__B2 _21496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11775_ _11834_/A _11770_/X _11774_/X VGND VGND VPWR VPWR _11775_/X sky130_fd_sc_hd__and3_4
XPHY_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16006_/A _16300_/X _16301_/X VGND VGND VPWR VPWR _16302_/X sky130_fd_sc_hd__and3_4
X_13514_ _13514_/A _13514_/B _13513_/X VGND VGND VPWR VPWR _13514_/X sky130_fd_sc_hd__and3_4
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14494_ _14506_/A _24027_/Q VGND VGND VPWR VPWR _14494_/X sky130_fd_sc_hd__or2_4
X_17282_ _17302_/B VGND VGND VPWR VPWR _17303_/B sky130_fd_sc_hd__inv_2
XANTENNA__20170__B2 IRQ[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19021_ _19021_/A VGND VGND VPWR VPWR _19021_/X sky130_fd_sc_hd__buf_2
X_16233_ _16202_/A _16149_/B VGND VGND VPWR VPWR _16233_/X sky130_fd_sc_hd__or2_4
X_13445_ _13468_/A _13445_/B _13445_/C VGND VGND VPWR VPWR _13445_/X sky130_fd_sc_hd__or3_4
XFILLER_16_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12616__A _12616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23958__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13376_ _13376_/A _13376_/B _13376_/C VGND VGND VPWR VPWR _13381_/B sky130_fd_sc_hd__and3_4
X_16164_ _13408_/A VGND VGND VPWR VPWR _16164_/X sky130_fd_sc_hd__buf_2
XFILLER_154_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12327_ _12327_/A VGND VGND VPWR VPWR _12580_/A sky130_fd_sc_hd__buf_2
X_15115_ _15649_/A _15099_/X _15115_/C VGND VGND VPWR VPWR _15116_/C sky130_fd_sc_hd__or3_4
XFILLER_103_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16095_ _12559_/A VGND VGND VPWR VPWR _16096_/A sky130_fd_sc_hd__buf_2
XFILLER_127_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14831__A _14658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19923_ _22922_/A VGND VGND VPWR VPWR _19924_/A sky130_fd_sc_hd__buf_2
XFILLER_48_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15046_ _11853_/A _11625_/X _15015_/X _11603_/A _15045_/X VGND VGND VPWR VPWR _15047_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_142_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12258_ _12258_/A VGND VGND VPWR VPWR _12702_/A sky130_fd_sc_hd__buf_2
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14550__B _14549_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19854_ _19471_/X _19850_/X _19851_/X _21370_/B _19552_/X VGND VGND VPWR VPWR _19854_/X
+ sky130_fd_sc_hd__a32o_4
X_12189_ _13627_/A VGND VGND VPWR VPWR _12190_/A sky130_fd_sc_hd__buf_2
X_18805_ _17156_/A _18803_/X _24458_/Q _18804_/X VGND VGND VPWR VPWR _18805_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21973__A2 _21967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19785_ _20598_/B _19518_/X _19784_/X _19638_/X VGND VGND VPWR VPWR _19785_/X sky130_fd_sc_hd__a211o_4
X_16997_ _16997_/A _16997_/B VGND VGND VPWR VPWR _17008_/A sky130_fd_sc_hd__or2_4
XFILLER_77_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15662__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18736_ _18735_/X VGND VGND VPWR VPWR _18736_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15948_ _15978_/A VGND VGND VPWR VPWR _16003_/A sky130_fd_sc_hd__buf_2
XFILLER_48_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21725__A2 _21720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18667_ _18399_/X VGND VGND VPWR VPWR _18667_/X sky130_fd_sc_hd__buf_2
X_15879_ _13529_/A _15879_/B _15879_/C VGND VGND VPWR VPWR _15880_/C sky130_fd_sc_hd__and3_4
XFILLER_37_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14278__A _14278_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13182__A _12866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16601__A1 _11984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17618_ _17632_/A VGND VGND VPWR VPWR _17618_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18598_ _17632_/D _17620_/B VGND VGND VPWR VPWR _18599_/B sky130_fd_sc_hd__or2_4
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17549_ _17548_/X VGND VGND VPWR VPWR _17659_/B sky130_fd_sc_hd__inv_2
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22150__A2 _22147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13910__A _14335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20560_ _20533_/X _20559_/X _24105_/Q _20510_/X VGND VGND VPWR VPWR _20560_/X sky130_fd_sc_hd__o22a_4
XFILLER_165_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19219_ _19219_/A VGND VGND VPWR VPWR _19219_/Y sky130_fd_sc_hd__inv_2
X_20491_ _24427_/Q _20318_/B VGND VGND VPWR VPWR _20491_/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12526__A _12473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22230_ _22244_/A VGND VGND VPWR VPWR _22230_/X sky130_fd_sc_hd__buf_2
XANTENNA__21839__A _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15837__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22161_ _20937_/A VGND VGND VPWR VPWR _22161_/X sky130_fd_sc_hd__buf_2
XFILLER_161_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21661__B2 _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14741__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21112_ _20659_/X _21111_/X _24036_/Q _21108_/X VGND VGND VPWR VPWR _24036_/D sky130_fd_sc_hd__o22a_4
X_22092_ _22147_/A VGND VGND VPWR VPWR _22118_/A sky130_fd_sc_hd__inv_2
XANTENNA__14460__B _14460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21413__A1 _21304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13357__A _13385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21043_ _20395_/X _21038_/X _16425_/B _21042_/X VGND VGND VPWR VPWR _21043_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21413__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12261__A _12266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24386__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16668__A _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15572__A _12461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24263__CLK _24271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22994_ _22993_/X VGND VGND VPWR VPWR HADDR[15] sky130_fd_sc_hd__inv_2
XFILLER_28_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21716__A2 _21713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_42_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_42_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19979__A _19951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21945_ _21941_/A VGND VGND VPWR VPWR _21960_/A sky130_fd_sc_hd__buf_2
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13092__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19790__B1 _16675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _21874_/X _21875_/X _23610_/Q _21870_/X VGND VGND VPWR VPWR _23610_/D sky130_fd_sc_hd__o22a_4
XFILLER_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ _23518_/CLK _21864_/X VGND VGND VPWR VPWR _23615_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22677__B1 _14387_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20827_ _20827_/A _20730_/B VGND VGND VPWR VPWR _20827_/X sky130_fd_sc_hd__or2_4
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19542__B1 HRDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23546_ _23515_/CLK _21982_/X VGND VGND VPWR VPWR _23546_/Q sky130_fd_sc_hd__dfxtp_4
X_11560_ _24449_/Q IRQ[12] VGND VGND VPWR VPWR _11560_/X sky130_fd_sc_hd__and2_4
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20758_ _20349_/A VGND VGND VPWR VPWR _20758_/X sky130_fd_sc_hd__buf_2
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23477_ _23617_/CLK _22087_/X VGND VGND VPWR VPWR _23477_/Q sky130_fd_sc_hd__dfxtp_4
X_20689_ _24259_/Q _20661_/X _20688_/X VGND VGND VPWR VPWR _20690_/B sky130_fd_sc_hd__o21a_4
XFILLER_10_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13230_/A _13161_/B VGND VGND VPWR VPWR _13230_/X sky130_fd_sc_hd__or2_4
X_22428_ _22113_/A VGND VGND VPWR VPWR _22428_/X sky130_fd_sc_hd__buf_2
XFILLER_136_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13161_ _13277_/A _13161_/B VGND VGND VPWR VPWR _13161_/X sky130_fd_sc_hd__or2_4
XANTENNA__15747__A _15778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21652__B2 _21617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22359_ _22366_/A VGND VGND VPWR VPWR _22359_/X sky130_fd_sc_hd__buf_2
XANTENNA__21761__A2_N _21760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14651__A _14647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12112_ _12111_/X VGND VGND VPWR VPWR _12112_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13092_ _13092_/A _13092_/B _13092_/C VGND VGND VPWR VPWR _13093_/C sky130_fd_sc_hd__and3_4
XANTENNA__15466__B _15466_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20207__A2 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24029_ _23880_/CLK _21121_/X VGND VGND VPWR VPWR _24029_/Q sky130_fd_sc_hd__dfxtp_4
X_16920_ _16912_/Y _17096_/A _16915_/C _16919_/X VGND VGND VPWR VPWR _16920_/X sky130_fd_sc_hd__a211o_4
X_12043_ _16561_/A _12043_/B _12042_/X VGND VGND VPWR VPWR _12043_/X sky130_fd_sc_hd__or3_4
XANTENNA__13267__A _13049_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_124_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR _23880_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21955__A2 _21953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17681__B _17456_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16851_ _13269_/X _16841_/B VGND VGND VPWR VPWR _16852_/D sky130_fd_sc_hd__nand2_4
XFILLER_133_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15802_ _12866_/A _15798_/X _15802_/C VGND VGND VPWR VPWR _15802_/X sky130_fd_sc_hd__or3_4
X_19570_ _19469_/X _19569_/X _17406_/Y _19515_/X VGND VGND VPWR VPWR _19570_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__21168__B1 _24000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16782_ _16621_/A _16782_/B VGND VGND VPWR VPWR _16782_/X sky130_fd_sc_hd__or2_4
XFILLER_18_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13994_ _12502_/A _23424_/Q VGND VGND VPWR VPWR _13995_/C sky130_fd_sc_hd__or2_4
XFILLER_20_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18521_ _18461_/A VGND VGND VPWR VPWR _18565_/A sky130_fd_sc_hd__buf_2
X_15733_ _13123_/A _15733_/B _15733_/C VGND VGND VPWR VPWR _15751_/B sky130_fd_sc_hd__and3_4
X_12945_ _12945_/A _12941_/X _12945_/C VGND VGND VPWR VPWR _12946_/C sky130_fd_sc_hd__or3_4
XANTENNA__14098__A _14138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18452_ _18400_/X _18451_/X _24483_/Q _18400_/X VGND VGND VPWR VPWR _18452_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15664_ _12689_/A _15726_/B VGND VGND VPWR VPWR _15664_/X sky130_fd_sc_hd__or2_4
XFILLER_73_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12876_ _12876_/A _23593_/Q VGND VGND VPWR VPWR _12877_/C sky130_fd_sc_hd__or2_4
X_17403_ _13945_/X _17438_/B VGND VGND VPWR VPWR _18557_/A sky130_fd_sc_hd__or2_4
X_14615_ _14615_/A VGND VGND VPWR VPWR _14660_/A sky130_fd_sc_hd__buf_2
XANTENNA__22668__B1 _15493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18383_ _17187_/X VGND VGND VPWR VPWR _18383_/Y sky130_fd_sc_hd__inv_2
X_11827_ _11832_/A _11827_/B VGND VGND VPWR VPWR _11827_/X sky130_fd_sc_hd__or2_4
X_15595_ _15595_/A VGND VGND VPWR VPWR _15612_/A sky130_fd_sc_hd__buf_2
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14826__A _14682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17623_/A _17333_/X VGND VGND VPWR VPWR _18709_/A sky130_fd_sc_hd__and2_4
X_11758_ _13414_/A VGND VGND VPWR VPWR _16214_/A sky130_fd_sc_hd__buf_2
X_14546_ _11813_/A _14546_/B _14546_/C VGND VGND VPWR VPWR _14547_/C sky130_fd_sc_hd__or3_4
XFILLER_53_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17265_ _17264_/X VGND VGND VPWR VPWR _17913_/B sky130_fd_sc_hd__inv_2
X_11689_ _12630_/A VGND VGND VPWR VPWR _11689_/X sky130_fd_sc_hd__buf_2
XANTENNA__12346__A _11739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14477_ _12504_/A _14477_/B VGND VGND VPWR VPWR _14477_/X sky130_fd_sc_hd__or2_4
X_19004_ _19004_/A VGND VGND VPWR VPWR _19004_/Y sky130_fd_sc_hd__inv_2
X_16216_ _16216_/A _16140_/B VGND VGND VPWR VPWR _16216_/X sky130_fd_sc_hd__or2_4
X_13428_ _13327_/A _13426_/X _13428_/C VGND VGND VPWR VPWR _13428_/X sky130_fd_sc_hd__and3_4
XANTENNA__21659__A _21674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17196_ _17120_/Y _17192_/X _14845_/Y _17193_/X VGND VGND VPWR VPWR _17196_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24136__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16147_ _16147_/A _24109_/Q VGND VGND VPWR VPWR _16148_/C sky130_fd_sc_hd__or2_4
X_13359_ _13374_/A _13286_/B VGND VGND VPWR VPWR _13361_/B sky130_fd_sc_hd__or2_4
XANTENNA__15657__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21643__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14561__A _14270_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18033__A _18032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16078_ _16066_/A _16078_/B _16078_/C VGND VGND VPWR VPWR _16078_/X sky130_fd_sc_hd__and3_4
XANTENNA__22199__A2 _22194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19906_ _19402_/A VGND VGND VPWR VPWR _19906_/X sky130_fd_sc_hd__buf_2
XANTENNA__17872__A _18413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15029_ _15029_/A _15025_/X _15029_/C VGND VGND VPWR VPWR _15029_/X sky130_fd_sc_hd__or3_4
XANTENNA__24286__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19837_ _19467_/X _19836_/X _19516_/X _19749_/X VGND VGND VPWR VPWR _19837_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16488__A _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15392__A _12530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13905__A _14507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19768_ _19787_/B _19767_/X _19687_/C VGND VGND VPWR VPWR _19768_/Y sky130_fd_sc_hd__o21ai_4
X_18719_ _18718_/X _18630_/C _18698_/X VGND VGND VPWR VPWR _18719_/X sky130_fd_sc_hd__a21o_4
XANTENNA__13624__B _13624_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_29_0_HCLK clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19699_ _19689_/X _19695_/X _19556_/X _19698_/X VGND VGND VPWR VPWR _19699_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22371__A2 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19772__B1 _16684_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21730_ _21558_/X _21727_/X _23687_/Q _21724_/X VGND VGND VPWR VPWR _23687_/D sky130_fd_sc_hd__o22a_4
XFILLER_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19949__D _19948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21661_ _21655_/Y _21660_/X _21526_/X _21660_/X VGND VGND VPWR VPWR _23732_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14736__A _13617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23400_ _23496_/CLK _23400_/D VGND VGND VPWR VPWR _13028_/B sky130_fd_sc_hd__dfxtp_4
X_20612_ _20612_/A VGND VGND VPWR VPWR _21560_/A sky130_fd_sc_hd__buf_2
X_24380_ _24382_/CLK _24380_/D HRESETn VGND VGND VPWR VPWR _19094_/A sky130_fd_sc_hd__dfstp_4
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21592_ _20938_/A VGND VGND VPWR VPWR _21592_/X sky130_fd_sc_hd__buf_2
XFILLER_162_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22953__A _22952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23331_ _23241_/CLK _23331_/D VGND VGND VPWR VPWR _23331_/Q sky130_fd_sc_hd__dfxtp_4
X_20543_ _20543_/A _20494_/B VGND VGND VPWR VPWR _20543_/X sky130_fd_sc_hd__or2_4
XFILLER_20_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21882__B2 _21809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12256__A _15439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23262_ _23679_/CLK _22465_/X VGND VGND VPWR VPWR _13702_/B sky130_fd_sc_hd__dfxtp_4
X_20474_ _20425_/X _20473_/X _24300_/Q _20349_/X VGND VGND VPWR VPWR _20474_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22213_ _22153_/X _22208_/X _14392_/B _22212_/X VGND VGND VPWR VPWR _23420_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15567__A _14430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20437__A2 _20423_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12914__A3 _12883_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23193_ _23194_/CLK _23193_/D VGND VGND VPWR VPWR _14713_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_133_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14471__A _11880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15313__A1 _13951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22144_ _22459_/A VGND VGND VPWR VPWR _22144_/X sky130_fd_sc_hd__buf_2
XFILLER_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15313__B2 _15312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14190__B _23743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22075_ _21862_/X _22074_/X _23487_/Q _22071_/X VGND VGND VPWR VPWR _22075_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21026_ _24084_/Q VGND VGND VPWR VPWR _21026_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16398__A _16009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13815__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22898__B1 _15915_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22977_ _22908_/A VGND VGND VPWR VPWR _22977_/X sky130_fd_sc_hd__buf_2
XFILLER_76_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12730_ _13164_/A _12819_/B VGND VGND VPWR VPWR _12730_/X sky130_fd_sc_hd__or2_4
XFILLER_16_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19502__A _19823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21928_ _21869_/X _21923_/X _14360_/B _21927_/X VGND VGND VPWR VPWR _23580_/D sky130_fd_sc_hd__o22a_4
XFILLER_16_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12661_ _12646_/A _12564_/B VGND VGND VPWR VPWR _12661_/X sky130_fd_sc_hd__or2_4
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _21857_/X _21851_/X _15555_/B _21858_/X VGND VGND VPWR VPWR _21859_/X sky130_fd_sc_hd__o22a_4
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22114__A2 _22111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _12583_/A _14400_/B VGND VGND VPWR VPWR _14400_/X sky130_fd_sc_hd__or2_4
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11612_ _17062_/D VGND VGND VPWR VPWR _18888_/B sky130_fd_sc_hd__buf_2
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12592_/A VGND VGND VPWR VPWR _12971_/A sky130_fd_sc_hd__buf_2
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15380_ _15380_/A VGND VGND VPWR VPWR _15381_/A sky130_fd_sc_hd__inv_2
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24159__CLK _24271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_49_0_HCLK clkbuf_7_49_0_HCLK/A VGND VGND VPWR VPWR _23922_/CLK sky130_fd_sc_hd__clkbuf_1
X_14331_ _14331_/A _14327_/X _14330_/X VGND VGND VPWR VPWR _14332_/B sky130_fd_sc_hd__or3_4
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _24369_/Q _11543_/B VGND VGND VPWR VPWR _18964_/A sky130_fd_sc_hd__or2_4
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23529_ _23241_/CLK _22011_/X VGND VGND VPWR VPWR _12916_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21873__B2 _21870_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17050_ _17418_/A VGND VGND VPWR VPWR _17050_/X sky130_fd_sc_hd__buf_2
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _14263_/B VGND VGND VPWR VPWR _14262_/X sky130_fd_sc_hd__buf_2
XANTENNA__19818__A1 _19724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17676__B _17482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16001_ _15969_/A _23662_/Q VGND VGND VPWR VPWR _16001_/X sky130_fd_sc_hd__or2_4
X_13213_ _13200_/X _23591_/Q VGND VGND VPWR VPWR _13214_/C sky130_fd_sc_hd__or2_4
XFILLER_13_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21625__B2 _21624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14193_ _15330_/A VGND VGND VPWR VPWR _14630_/A sky130_fd_sc_hd__buf_2
XANTENNA__24216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13144_ _13164_/A _23687_/Q VGND VGND VPWR VPWR _13146_/B sky130_fd_sc_hd__or2_4
XFILLER_125_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13075_ _13085_/A _23592_/Q VGND VGND VPWR VPWR _13076_/C sky130_fd_sc_hd__or2_4
X_17952_ _17920_/X _17943_/Y _17944_/X _17951_/Y VGND VGND VPWR VPWR _17952_/X sky130_fd_sc_hd__a211o_4
XFILLER_3_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21389__B1 _12665_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21928__A2 _21923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16903_ _11644_/X VGND VGND VPWR VPWR _16915_/C sky130_fd_sc_hd__buf_2
X_12026_ _12025_/X VGND VGND VPWR VPWR _16905_/A sky130_fd_sc_hd__buf_2
X_17883_ _17882_/X VGND VGND VPWR VPWR _17883_/X sky130_fd_sc_hd__buf_2
XFILLER_78_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22103__A _20377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19622_ _19687_/A _19622_/B VGND VGND VPWR VPWR _19622_/X sky130_fd_sc_hd__or2_4
XANTENNA__13725__A _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16834_ _12683_/X _16833_/X _12682_/A VGND VGND VPWR VPWR _16834_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18006__B1 _17919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19553_ _19552_/X VGND VGND VPWR VPWR _19553_/X sky130_fd_sc_hd__buf_2
X_16765_ _16755_/X _24049_/Q VGND VGND VPWR VPWR _16767_/B sky130_fd_sc_hd__or2_4
XANTENNA__22889__B1 _14086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13977_ _12474_/A _23168_/Q VGND VGND VPWR VPWR _13979_/B sky130_fd_sc_hd__or2_4
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18504_ _18032_/X VGND VGND VPWR VPWR _18504_/X sky130_fd_sc_hd__buf_2
XFILLER_34_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15716_ _13307_/A _15693_/X _15700_/X _15707_/X _15715_/X VGND VGND VPWR VPWR _15716_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_80_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12928_ _12940_/A _23305_/Q VGND VGND VPWR VPWR _12929_/C sky130_fd_sc_hd__or2_4
X_19484_ _19442_/X VGND VGND VPWR VPWR _19484_/X sky130_fd_sc_hd__buf_2
X_16696_ _16561_/A _16692_/X _16696_/C VGND VGND VPWR VPWR _16696_/X sky130_fd_sc_hd__or3_4
XANTENNA__20558__A _20558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18435_ _18022_/X _18368_/X _18432_/Y _18027_/X _22984_/B VGND VGND VPWR VPWR _18435_/X
+ sky130_fd_sc_hd__a32o_4
X_15647_ _14348_/A _15643_/X _15647_/C VGND VGND VPWR VPWR _15647_/X sky130_fd_sc_hd__or3_4
X_12859_ _12884_/A _12922_/B VGND VGND VPWR VPWR _12861_/B sky130_fd_sc_hd__or2_4
XFILLER_22_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14556__A _14278_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13460__A _13474_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18366_ _18478_/A _18365_/X VGND VGND VPWR VPWR _18366_/X sky130_fd_sc_hd__or2_4
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15578_ _13687_/A _15578_/B _15577_/X VGND VGND VPWR VPWR _15579_/C sky130_fd_sc_hd__and3_4
XFILLER_109_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17317_ _17315_/Y _17316_/X VGND VGND VPWR VPWR _17318_/A sky130_fd_sc_hd__or2_4
X_14529_ _14513_/A _14525_/X _14528_/X VGND VGND VPWR VPWR _14530_/C sky130_fd_sc_hd__or3_4
XFILLER_174_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18297_ _17517_/Y _18296_/X VGND VGND VPWR VPWR _18297_/X sky130_fd_sc_hd__or2_4
XANTENNA__21864__B2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17248_ _17111_/X _18734_/B _17224_/X _17247_/X VGND VGND VPWR VPWR _17248_/X sky130_fd_sc_hd__a211o_4
XFILLER_174_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21616__B2 _21610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_6_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17179_ _17128_/X _17175_/X _17836_/A _17178_/X VGND VGND VPWR VPWR _17179_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12804__A _12834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21092__A2 _21090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20190_ _20125_/A _20190_/B VGND VGND VPWR VPWR _20191_/B sky130_fd_sc_hd__or2_4
XANTENNA__23676__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21919__A2 _21916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13635__A _15446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22900_ _22897_/A _22899_/X VGND VGND VPWR VPWR HWDATA[30] sky130_fd_sc_hd__nor2_4
X_23880_ _23880_/CLK _23880_/D VGND VGND VPWR VPWR _23880_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16011__A _16011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22831_ _22814_/X _22830_/X VGND VGND VPWR VPWR HWDATA[11] sky130_fd_sc_hd__nor2_4
XFILLER_38_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15850__A _12373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22762_ SYSTICKCLKDIV[6] VGND VGND VPWR VPWR _22762_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21713_ _21727_/A VGND VGND VPWR VPWR _21713_/X sky130_fd_sc_hd__buf_2
XANTENNA__17220__A1 _12077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24301__CLK _24302_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _22722_/A VGND VGND VPWR VPWR _22708_/A sky130_fd_sc_hd__buf_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21644_ _21582_/X _21641_/X _23741_/Q _21638_/X VGND VGND VPWR VPWR _21644_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20107__A1 _19906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24432_ _23379_/CLK _18848_/X HRESETn VGND VGND VPWR VPWR _24432_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24363_ _24357_/CLK _24363_/D HRESETn VGND VGND VPWR VPWR _19004_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__11602__B _11590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ _20770_/A VGND VGND VPWR VPWR _21575_/X sky130_fd_sc_hd__buf_2
XFILLER_36_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16681__A _16659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18720__B2 _18719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23314_ _23922_/CLK _22364_/X VGND VGND VPWR VPWR _16627_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_138_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20526_ _20526_/A VGND VGND VPWR VPWR _20526_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21299__A _20860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24294_ _24294_/CLK _24294_/D HRESETn VGND VGND VPWR VPWR _24294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23245_ _23533_/CLK _22503_/X VGND VGND VPWR VPWR _16149_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19992__A _18670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15297__A _14574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20457_ _18140_/X _20446_/X _20638_/A _20456_/Y VGND VGND VPWR VPWR _20457_/X sky130_fd_sc_hd__a211o_4
XFILLER_10_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17287__A1 _17284_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23176_ _23496_/CLK _23176_/D VGND VGND VPWR VPWR _13012_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_161_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20388_ _20388_/A _20387_/X VGND VGND VPWR VPWR _20388_/Y sky130_fd_sc_hd__nor2_4
XFILLER_134_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20291__B1 _20343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22127_ _20595_/A VGND VGND VPWR VPWR _22127_/X sky130_fd_sc_hd__buf_2
XFILLER_47_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22058_ _21833_/X _22053_/X _12668_/B _22057_/X VGND VGND VPWR VPWR _22058_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23019__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22032__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13545__A _12971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21009_ _20943_/A _21008_/X VGND VGND VPWR VPWR _21009_/X sky130_fd_sc_hd__and2_4
X_13900_ _14390_/A _13900_/B VGND VGND VPWR VPWR _13900_/X sky130_fd_sc_hd__or2_4
X_14880_ _14096_/A _14880_/B VGND VGND VPWR VPWR _14880_/X sky130_fd_sc_hd__or2_4
XANTENNA__21762__A _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13831_ _15395_/A _13831_/B VGND VGND VPWR VPWR _13831_/X sky130_fd_sc_hd__or2_4
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19736__B1 _19705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15760__A _12783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16550_ _11939_/X _16550_/B _16550_/C VGND VGND VPWR VPWR _16550_/X sky130_fd_sc_hd__or3_4
X_13762_ _12587_/A _13760_/X _13762_/C VGND VGND VPWR VPWR _13763_/C sky130_fd_sc_hd__and3_4
Xclkbuf_5_12_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_15501_ _15477_/A _15501_/B VGND VGND VPWR VPWR _15501_/X sky130_fd_sc_hd__or2_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12713_ _12702_/A _12797_/B VGND VGND VPWR VPWR _12713_/X sky130_fd_sc_hd__or2_4
X_16481_ _13385_/A VGND VGND VPWR VPWR _16481_/X sky130_fd_sc_hd__buf_2
X_13693_ _12367_/A VGND VGND VPWR VPWR _14372_/A sky130_fd_sc_hd__buf_2
X_18220_ _18220_/A VGND VGND VPWR VPWR _18405_/A sky130_fd_sc_hd__buf_2
X_15432_ _12191_/A _15432_/B VGND VGND VPWR VPWR _15432_/X sky130_fd_sc_hd__or2_4
X_12644_ _12644_/A _23979_/Q VGND VGND VPWR VPWR _12645_/C sky130_fd_sc_hd__or2_4
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22593__A _22622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12608__B _12608_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18151_ _18222_/A _17537_/Y VGND VGND VPWR VPWR _18155_/B sky130_fd_sc_hd__and2_4
X_12575_ _11681_/A VGND VGND VPWR VPWR _12576_/A sky130_fd_sc_hd__buf_2
X_15363_ _15326_/A _15304_/B VGND VGND VPWR VPWR _15365_/B sky130_fd_sc_hd__or2_4
XFILLER_129_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17102_ _17101_/Y VGND VGND VPWR VPWR _18440_/A sky130_fd_sc_hd__buf_2
X_14314_ _15402_/A _14391_/B VGND VGND VPWR VPWR _14316_/B sky130_fd_sc_hd__or2_4
XFILLER_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11526_ _24352_/Q _11525_/X VGND VGND VPWR VPWR _11526_/X sky130_fd_sc_hd__or2_4
X_18082_ _17229_/X _17843_/X _17823_/A _17859_/X VGND VGND VPWR VPWR _18083_/A sky130_fd_sc_hd__o22a_4
XFILLER_141_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15294_ _15294_/A _23416_/Q VGND VGND VPWR VPWR _15294_/X sky130_fd_sc_hd__or2_4
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14823__B _23417_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17033_ _17033_/A VGND VGND VPWR VPWR _17481_/B sky130_fd_sc_hd__inv_2
XFILLER_109_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14245_ _14240_/A _23807_/Q VGND VGND VPWR VPWR _14245_/X sky130_fd_sc_hd__or2_4
XFILLER_109_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15000__A _15000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14176_ _11663_/A VGND VGND VPWR VPWR _14614_/A sky130_fd_sc_hd__buf_2
XANTENNA__21074__A2 _21073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22271__B2 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20841__A _20841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15935__A _15934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13127_ _12693_/A _23271_/Q VGND VGND VPWR VPWR _13129_/B sky130_fd_sc_hd__or2_4
XANTENNA__19407__A _19406_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18984_ _18963_/X _18982_/X _18983_/Y _18968_/X VGND VGND VPWR VPWR _18984_/X sky130_fd_sc_hd__o22a_4
X_13058_ _13058_/A VGND VGND VPWR VPWR _13096_/A sky130_fd_sc_hd__buf_2
X_17935_ _17934_/X VGND VGND VPWR VPWR _17935_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22023__B2 _22021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13455__A _13455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12009_ _11951_/X _12009_/B _12009_/C VGND VGND VPWR VPWR _12010_/C sky130_fd_sc_hd__and3_4
X_17866_ _17809_/X _17846_/X _17848_/X _17865_/X VGND VGND VPWR VPWR _17867_/A sky130_fd_sc_hd__o22a_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16817_ _16683_/A _16809_/X _16816_/X VGND VGND VPWR VPWR _16818_/C sky130_fd_sc_hd__and3_4
X_19605_ _19604_/Y _19788_/A VGND VGND VPWR VPWR _19605_/X sky130_fd_sc_hd__and2_4
XANTENNA__24324__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17797_ _17797_/A VGND VGND VPWR VPWR _17798_/A sky130_fd_sc_hd__buf_2
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15670__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19536_ _19504_/B VGND VGND VPWR VPWR _19623_/A sky130_fd_sc_hd__inv_2
XFILLER_53_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16748_ _11868_/X _16748_/B VGND VGND VPWR VPWR _16748_/X sky130_fd_sc_hd__and2_4
XANTENNA__20288__A _20267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19467_ _19859_/A VGND VGND VPWR VPWR _19467_/X sky130_fd_sc_hd__buf_2
XFILLER_62_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14286__A _13823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16679_ _16672_/A _16679_/B VGND VGND VPWR VPWR _16679_/X sky130_fd_sc_hd__or2_4
XANTENNA__13190__A _11864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18418_ _18418_/A VGND VGND VPWR VPWR _18418_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24474__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19398_ _19396_/X _18149_/X _19396_/X _24236_/Q VGND VGND VPWR VPWR _19398_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12518__B _12619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18349_ _17509_/Y _18348_/B _18176_/X VGND VGND VPWR VPWR _18349_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21837__B2 _21834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24138__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_32_0_HCLK clkbuf_6_16_0_HCLK/X VGND VGND VPWR VPWR _23668_/CLK sky130_fd_sc_hd__clkbuf_1
X_21360_ _21299_/X _21355_/X _14376_/B _21359_/X VGND VGND VPWR VPWR _21360_/X sky130_fd_sc_hd__o22a_4
X_20311_ _20259_/A VGND VGND VPWR VPWR _20847_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_95_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR _23772_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_162_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21291_ _21290_/X _21281_/X _14035_/B _21288_/X VGND VGND VPWR VPWR _23936_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12534__A _12487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23030_ _23043_/A _23030_/B VGND VGND VPWR VPWR _23030_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21065__A2 _21059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20242_ _20865_/A HRDATA[7] _19908_/A VGND VGND VPWR VPWR _20242_/X sky130_fd_sc_hd__o21a_4
XANTENNA__11553__A2 IRQ[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15845__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20173_ _20165_/Y _20166_/Y _11565_/X _20172_/X VGND VGND VPWR VPWR _20173_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_3_1_0_HCLK clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23932_ _23515_/CLK _23932_/D VGND VGND VPWR VPWR _14359_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20576__A1 _20533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21773__B1 _23660_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20576__B2 _20510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21582__A _20841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23863_ _23194_/CLK _23863_/D VGND VGND VPWR VPWR _15180_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22317__A2 _22315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15580__A _13689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22814_ _22884_/A VGND VGND VPWR VPWR _22814_/X sky130_fd_sc_hd__buf_2
X_23794_ _23728_/CLK _23794_/D VGND VGND VPWR VPWR _23794_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22745_ _22745_/A _22737_/X VGND VGND VPWR VPWR _22745_/Y sky130_fd_sc_hd__nor2_4
XFILLER_38_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18941__A1 _15118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22676_ _22655_/A VGND VGND VPWR VPWR _22676_/X sky130_fd_sc_hd__buf_2
XFILLER_13_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21627_ _21620_/A VGND VGND VPWR VPWR _21627_/X sky130_fd_sc_hd__buf_2
XFILLER_139_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24415_ _24419_/CLK _18873_/X HRESETn VGND VGND VPWR VPWR _24415_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21828__B2 _21822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12360_ _13248_/A VGND VGND VPWR VPWR _12407_/A sky130_fd_sc_hd__buf_2
XANTENNA__17300__A _14844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21558_ _20596_/A VGND VGND VPWR VPWR _21558_/X sky130_fd_sc_hd__buf_2
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24346_ _24382_/CLK _24346_/D HRESETn VGND VGND VPWR VPWR _11520_/A sky130_fd_sc_hd__dfstp_4
X_20509_ _20509_/A VGND VGND VPWR VPWR _20509_/X sky130_fd_sc_hd__buf_2
XFILLER_153_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12291_ _12239_/A VGND VGND VPWR VPWR _13183_/A sky130_fd_sc_hd__buf_2
X_24277_ _24277_/CLK _24277_/D HRESETn VGND VGND VPWR VPWR _19226_/B sky130_fd_sc_hd__dfrtp_4
X_21489_ _21489_/A VGND VGND VPWR VPWR _21489_/X sky130_fd_sc_hd__buf_2
XANTENNA__12444__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14030_ _12580_/A VGND VGND VPWR VPWR _14056_/A sky130_fd_sc_hd__buf_2
X_23228_ _23587_/CLK _22527_/X VGND VGND VPWR VPWR _14406_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23991__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22253__B2 _22248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23159_ _23862_/CLK _23159_/D VGND VGND VPWR VPWR _15149_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_134_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18472__A3 _18465_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18209__B1 _18060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22005__B2 _22000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15474__B _15474_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15981_ _15944_/A _16054_/B VGND VGND VPWR VPWR _15981_/X sky130_fd_sc_hd__or2_4
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23221__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13275__A _13318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22556__A2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17720_ _17720_/A _17720_/B VGND VGND VPWR VPWR _17720_/X sky130_fd_sc_hd__or2_4
X_14932_ _15377_/A _14921_/X _14931_/X VGND VGND VPWR VPWR _14932_/X sky130_fd_sc_hd__and3_4
XANTENNA__17970__A _18407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21492__A _21492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17651_ _16943_/X _17012_/X _17014_/X _17650_/X VGND VGND VPWR VPWR _17651_/X sky130_fd_sc_hd__o22a_4
XFILLER_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14863_ _14133_/A _14863_/B _14862_/X VGND VGND VPWR VPWR _14863_/X sky130_fd_sc_hd__or3_4
XFILLER_75_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16602_ _11858_/X _11632_/X _16570_/X _11608_/X _16601_/X VGND VGND VPWR VPWR _16602_/X
+ sky130_fd_sc_hd__a32o_4
X_13814_ _12497_/A _23677_/Q VGND VGND VPWR VPWR _13814_/X sky130_fd_sc_hd__or2_4
X_17582_ _18113_/B VGND VGND VPWR VPWR _18138_/A sky130_fd_sc_hd__inv_2
X_14794_ _14841_/A _14782_/X _14793_/X VGND VGND VPWR VPWR _14794_/X sky130_fd_sc_hd__and3_4
XFILLER_169_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19321_ _19321_/A VGND VGND VPWR VPWR _19321_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16533_ _15933_/X _16528_/X _16532_/Y VGND VGND VPWR VPWR _16533_/X sky130_fd_sc_hd__o21a_4
X_13745_ _12610_/A _23550_/Q VGND VGND VPWR VPWR _13745_/X sky130_fd_sc_hd__or2_4
XANTENNA__17196__B1 _14845_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18932__A1 _13945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19252_ _19252_/A _19252_/B VGND VGND VPWR VPWR _19253_/B sky130_fd_sc_hd__and2_4
X_16464_ _16454_/A _16395_/B VGND VGND VPWR VPWR _16464_/X sky130_fd_sc_hd__or2_4
X_13676_ _13676_/A _24094_/Q VGND VGND VPWR VPWR _13677_/C sky130_fd_sc_hd__or2_4
X_18203_ _17874_/X _18086_/X _18053_/X VGND VGND VPWR VPWR _18203_/Y sky130_fd_sc_hd__o21ai_4
X_15415_ _15415_/A _15413_/X _15414_/X VGND VGND VPWR VPWR _15415_/X sky130_fd_sc_hd__and3_4
X_12627_ _12974_/A _23467_/Q VGND VGND VPWR VPWR _12628_/C sky130_fd_sc_hd__or2_4
X_19183_ _19151_/B VGND VGND VPWR VPWR _19183_/Y sky130_fd_sc_hd__inv_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16395_ _16009_/X _16395_/B VGND VGND VPWR VPWR _16395_/X sky130_fd_sc_hd__or2_4
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18134_ _18131_/X _18133_/X _18053_/X VGND VGND VPWR VPWR _18134_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18696__B1 _18691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15346_ _15362_/A _15338_/X _15346_/C VGND VGND VPWR VPWR _15346_/X sky130_fd_sc_hd__and3_4
X_12558_ _12568_/A VGND VGND VPWR VPWR _12559_/A sky130_fd_sc_hd__buf_2
Xclkbuf_6_19_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22492__B2 _22491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14553__B _14618_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18065_ _18064_/X VGND VGND VPWR VPWR _18065_/X sky130_fd_sc_hd__buf_2
XFILLER_8_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12354__A _12354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15277_ _14169_/A _23160_/Q VGND VGND VPWR VPWR _15279_/B sky130_fd_sc_hd__or2_4
X_12489_ _12869_/A _12489_/B _12488_/X VGND VGND VPWR VPWR _12490_/C sky130_fd_sc_hd__and3_4
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17016_ _17038_/A _17038_/B _17016_/C _11598_/D VGND VGND VPWR VPWR _17017_/B sky130_fd_sc_hd__or4_4
XANTENNA__21047__A2 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21667__A _21667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14228_ _14631_/A _14228_/B _14228_/C VGND VGND VPWR VPWR _14228_/X sky130_fd_sc_hd__and3_4
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15665__A _12690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14159_ _15007_/A VGND VGND VPWR VPWR _14988_/A sky130_fd_sc_hd__buf_2
XANTENNA__18041__A _18545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18967_ _18960_/X VGND VGND VPWR VPWR _19021_/A sky130_fd_sc_hd__buf_2
XFILLER_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22547__A2 _22544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17918_ _17109_/X VGND VGND VPWR VPWR _18168_/A sky130_fd_sc_hd__buf_2
X_18898_ _18896_/A VGND VGND VPWR VPWR _18928_/A sky130_fd_sc_hd__inv_2
XANTENNA__22498__A _22498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17849_ _17849_/A VGND VGND VPWR VPWR _17849_/X sky130_fd_sc_hd__buf_2
XANTENNA__16496__A _16370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13913__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20860_ _20860_/A VGND VGND VPWR VPWR _20860_/X sky130_fd_sc_hd__buf_2
XANTENNA__21507__B1 _23807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19519_ _19474_/X VGND VGND VPWR VPWR _19519_/X sky130_fd_sc_hd__buf_2
X_20791_ _20264_/X VGND VGND VPWR VPWR _20791_/X sky130_fd_sc_hd__buf_2
XANTENNA__23864__CLK _23864_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17187__B1 _18744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12529__A _14295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24319__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18923__A1 _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22530_ _22473_/X _22529_/X _14600_/B _22526_/X VGND VGND VPWR VPWR _23226_/D sky130_fd_sc_hd__o22a_4
XFILLER_90_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20746__A _20510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22461_ _22461_/A VGND VGND VPWR VPWR _22461_/X sky130_fd_sc_hd__buf_2
XFILLER_33_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14744__A _13655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24200_ _24184_/CLK _19760_/X HRESETn VGND VGND VPWR VPWR _13792_/A sky130_fd_sc_hd__dfrtp_4
X_21412_ _21405_/A VGND VGND VPWR VPWR _21412_/X sky130_fd_sc_hd__buf_2
XANTENNA__17120__A _16523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21286__A2 _21281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18687__B1 _18467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22392_ _22149_/X _22390_/X _13624_/B _22387_/X VGND VGND VPWR VPWR _23294_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22483__B2 _22421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14463__B _14463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24131_ _23126_/CLK _20209_/Y HRESETn VGND VGND VPWR VPWR _24131_/Q sky130_fd_sc_hd__dfrtp_4
X_21343_ _21271_/X _21341_/X _13018_/B _21338_/X VGND VGND VPWR VPWR _21343_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16162__A1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12264__A _11606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22228__A2_N _22227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24062_ _23997_/CLK _24062_/D VGND VGND VPWR VPWR _24062_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21577__A _20801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21274_ _21273_/X _21269_/X _23943_/Q _21264_/X VGND VGND VPWR VPWR _23943_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22235__B2 _22234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20481__A _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23013_ _23013_/A VGND VGND VPWR VPWR HADDR[18] sky130_fd_sc_hd__inv_2
X_20225_ _20396_/A VGND VGND VPWR VPWR _20225_/X sky130_fd_sc_hd__buf_2
XFILLER_2_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15575__A _12427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20156_ _20125_/B VGND VGND VPWR VPWR _20156_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13807__B _13807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18886__A _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11608__A _11608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20087_ _20087_/A VGND VGND VPWR VPWR _20087_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21210__A2 _21205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23915_ _24074_/CLK _23915_/D VGND VGND VPWR VPWR _12533_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22201__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13823__A _13823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23846_ _23397_/CLK _21446_/X VGND VGND VPWR VPWR _23846_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_150_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11860_ _14012_/A VGND VGND VPWR VPWR _13586_/A sky130_fd_sc_hd__buf_2
XFILLER_26_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _11704_/X VGND VGND VPWR VPWR _16635_/A sky130_fd_sc_hd__buf_2
XFILLER_60_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12439__A _12848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23777_ _23744_/CLK _23777_/D VGND VGND VPWR VPWR _23777_/Q sky130_fd_sc_hd__dfxtp_4
X_20989_ _20988_/Y _20493_/A VGND VGND VPWR VPWR _20989_/X sky130_fd_sc_hd__or2_4
XPHY_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22710__A2 _22708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _13530_/A _13510_/X _13530_/C VGND VGND VPWR VPWR _13566_/B sky130_fd_sc_hd__or3_4
XPHY_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22728_ _20892_/A _22722_/X _14531_/B _22726_/X VGND VGND VPWR VPWR _23099_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20656__A _20857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23032__A _18210_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13461_ _13475_/A _13457_/X _13461_/C VGND VGND VPWR VPWR _13461_/X sky130_fd_sc_hd__or3_4
XFILLER_55_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22659_ _22437_/X _22658_/X _23145_/Q _22655_/X VGND VGND VPWR VPWR _22659_/X sky130_fd_sc_hd__o22a_4
XFILLER_139_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15200_ _14616_/A _15200_/B _15199_/X VGND VGND VPWR VPWR _15200_/X sky130_fd_sc_hd__and3_4
X_12412_ _12373_/X _12303_/B VGND VGND VPWR VPWR _12412_/X sky130_fd_sc_hd__or2_4
X_16180_ _13413_/A VGND VGND VPWR VPWR _16185_/A sky130_fd_sc_hd__buf_2
XANTENNA__21277__A2 _21269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18678__B1 _17594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13392_ _13392_/A _13392_/B _13392_/C VGND VGND VPWR VPWR _13400_/B sky130_fd_sc_hd__or3_4
XFILLER_16_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22871__A _22870_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15131_ _14149_/A _15129_/X _15131_/C VGND VGND VPWR VPWR _15131_/X sky130_fd_sc_hd__and3_4
X_12343_ _11689_/X _12343_/B _12342_/X VGND VGND VPWR VPWR _12343_/X sky130_fd_sc_hd__or3_4
X_24329_ _24342_/CLK _19184_/X HRESETn VGND VGND VPWR VPWR _24329_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12274_ _12698_/A _12274_/B _12274_/C VGND VGND VPWR VPWR _12274_/X sky130_fd_sc_hd__and3_4
XFILLER_126_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15062_ _15075_/A _24021_/Q VGND VGND VPWR VPWR _15064_/B sky130_fd_sc_hd__or2_4
XANTENNA__17684__B _17511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15485__A _13229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14013_ _11967_/A _13989_/X _13996_/X _14004_/X _14012_/X VGND VGND VPWR VPWR _14013_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_122_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19870_ _19861_/X _19869_/X _19613_/X VGND VGND VPWR VPWR _19870_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_49_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18821_ _17153_/A _18817_/X _24446_/Q _18818_/X VGND VGND VPWR VPWR _18821_/X sky130_fd_sc_hd__o22a_4
XFILLER_150_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18796__A _18796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18752_ _18131_/X _18751_/X _18200_/X _18387_/X VGND VGND VPWR VPWR _18753_/A sky130_fd_sc_hd__o22a_4
X_15964_ _15960_/A _24014_/Q VGND VGND VPWR VPWR _15965_/C sky130_fd_sc_hd__or2_4
XFILLER_0_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17703_ _17703_/A _17483_/Y VGND VGND VPWR VPWR _17703_/X sky130_fd_sc_hd__or2_4
XANTENNA__21201__A2 _21198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14915_ _11697_/A _14915_/B _14914_/X VGND VGND VPWR VPWR _14921_/B sky130_fd_sc_hd__and3_4
X_18683_ _18032_/X _18681_/X _16943_/A _18682_/X VGND VGND VPWR VPWR _18683_/X sky130_fd_sc_hd__o22a_4
X_15895_ _13529_/A _15887_/X _15894_/X VGND VGND VPWR VPWR _15911_/B sky130_fd_sc_hd__and3_4
XANTENNA__22111__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17634_ _18557_/B VGND VGND VPWR VPWR _17635_/D sky130_fd_sc_hd__inv_2
X_14846_ _14766_/X _14845_/Y VGND VGND VPWR VPWR _15387_/B sky130_fd_sc_hd__or2_4
XANTENNA__20960__A1 _20894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24483__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20960__B2 _20861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21950__A _21950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17565_ _18035_/B VGND VGND VPWR VPWR _17583_/B sky130_fd_sc_hd__inv_2
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14777_ _15080_/A _23513_/Q VGND VGND VPWR VPWR _14778_/C sky130_fd_sc_hd__or2_4
XANTENNA__18905__A1 _16523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22162__B1 _14731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11989_ _12012_/A VGND VGND VPWR VPWR _11990_/A sky130_fd_sc_hd__buf_2
X_19304_ _19234_/A _19234_/B _19303_/Y VGND VGND VPWR VPWR _24285_/D sky130_fd_sc_hd__o21a_4
XANTENNA__24412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16516_ _16166_/X _16439_/B VGND VGND VPWR VPWR _16517_/C sky130_fd_sc_hd__or2_4
X_13728_ _13742_/A _13624_/B VGND VGND VPWR VPWR _13728_/X sky130_fd_sc_hd__or2_4
XANTENNA__20712__A1 _18472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17496_ _17495_/X VGND VGND VPWR VPWR _17496_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19235_ _19235_/A _19235_/B VGND VGND VPWR VPWR _19236_/B sky130_fd_sc_hd__and2_4
X_16447_ _11917_/X _16445_/X _16446_/X VGND VGND VPWR VPWR _16448_/C sky130_fd_sc_hd__and3_4
X_13659_ _13632_/A _24062_/Q VGND VGND VPWR VPWR _13659_/X sky130_fd_sc_hd__or2_4
XANTENNA__14564__A _12454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19166_ _19159_/A _19159_/B _19165_/Y VGND VGND VPWR VPWR _24338_/D sky130_fd_sc_hd__o21a_4
X_16378_ _11684_/X _16369_/X _16377_/X VGND VGND VPWR VPWR _16378_/X sky130_fd_sc_hd__and3_4
XANTENNA__22465__B2 _22457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23267__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18117_ _17101_/Y VGND VGND VPWR VPWR _18378_/A sky130_fd_sc_hd__buf_2
X_15329_ _13695_/A _15326_/X _15328_/X VGND VGND VPWR VPWR _15329_/X sky130_fd_sc_hd__and3_4
X_19097_ _19082_/X _19095_/X _19096_/X _11522_/A VGND VGND VPWR VPWR _24348_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19881__A2 _19811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18048_ _17878_/X _17217_/X _17878_/X _17202_/Y VGND VGND VPWR VPWR _18048_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22217__B2 _22212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15395__A _15395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13908__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12812__A _12800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20010_ _19992_/X _18070_/A _19998_/X _20009_/X VGND VGND VPWR VPWR _20010_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21440__A2 _21434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19999_ _19999_/A VGND VGND VPWR VPWR _19999_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21961_ _21838_/X _21960_/X _23561_/Q _21957_/X VGND VGND VPWR VPWR _21961_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14739__A _13652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22021__A _22007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23700_ _23668_/CLK _23700_/D VGND VGND VPWR VPWR _21705_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__13643__A _13652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20912_ _20977_/A _20911_/X VGND VGND VPWR VPWR _20912_/Y sky130_fd_sc_hd__nand2_4
X_21892_ _21899_/A VGND VGND VPWR VPWR _21892_/X sky130_fd_sc_hd__buf_2
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23631_ _23918_/CLK _21825_/X VGND VGND VPWR VPWR _16282_/B sky130_fd_sc_hd__dfxtp_4
X_20843_ HRDATA[7] _20843_/B VGND VGND VPWR VPWR _20843_/X sky130_fd_sc_hd__or2_4
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12259__A _12702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23562_ _23467_/CLK _21959_/X VGND VGND VPWR VPWR _12804_/B sky130_fd_sc_hd__dfxtp_4
X_20774_ _18597_/Y VGND VGND VPWR VPWR _20935_/A sky130_fd_sc_hd__buf_2
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22513_ _22444_/X _22508_/X _23238_/Q _22512_/X VGND VGND VPWR VPWR _22513_/X sky130_fd_sc_hd__o22a_4
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23493_ _23493_/CLK _23493_/D VGND VGND VPWR VPWR _13469_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_149_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14474__A _15400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24346__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22444_ _20612_/A VGND VGND VPWR VPWR _22444_/X sky130_fd_sc_hd__buf_2
XFILLER_149_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22691__A _22698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24192__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22375_ _22120_/X _22369_/X _12785_/B _22373_/X VGND VGND VPWR VPWR _23306_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24114_ _23404_/CLK _24114_/D VGND VGND VPWR VPWR _24114_/Q sky130_fd_sc_hd__dfxtp_4
X_21326_ _21322_/A VGND VGND VPWR VPWR _21341_/A sky130_fd_sc_hd__buf_2
XFILLER_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24045_ _24045_/CLK _21099_/X VGND VGND VPWR VPWR _24045_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_159_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21257_ _21269_/A VGND VGND VPWR VPWR _21257_/X sky130_fd_sc_hd__buf_2
XFILLER_85_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13818__A _13658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12722__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20208_ _19402_/A _17751_/A _20200_/A _20207_/X VGND VGND VPWR VPWR _20208_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21188_ _21195_/A VGND VGND VPWR VPWR _21188_/X sky130_fd_sc_hd__buf_2
XFILLER_89_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20139_ _11572_/X _20138_/X _20109_/Y VGND VGND VPWR VPWR _20139_/X sky130_fd_sc_hd__o21a_4
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12961_ _12659_/A _12957_/X _12961_/C VGND VGND VPWR VPWR _12961_/X sky130_fd_sc_hd__or3_4
XFILLER_38_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14649__A _14657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22392__B1 _13624_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14700_ _11668_/A _14700_/B _14699_/X VGND VGND VPWR VPWR _14700_/X sky130_fd_sc_hd__and3_4
X_11912_ _11912_/A VGND VGND VPWR VPWR _11913_/A sky130_fd_sc_hd__buf_2
X_15680_ _12279_/A _15680_/B _15679_/X VGND VGND VPWR VPWR _15680_/X sky130_fd_sc_hd__and3_4
X_12892_ _12864_/A _23849_/Q VGND VGND VPWR VPWR _12892_/X sky130_fd_sc_hd__or2_4
XFILLER_161_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21770__A _21770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14631_ _14631_/A VGND VGND VPWR VPWR _14667_/A sky130_fd_sc_hd__buf_2
X_11843_ _12167_/A _24116_/Q VGND VGND VPWR VPWR _11844_/C sky130_fd_sc_hd__or2_4
XFILLER_45_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23829_ _23456_/CLK _23829_/D VGND VGND VPWR VPWR _23829_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17350_ _17630_/A _17350_/B VGND VGND VPWR VPWR _18600_/A sky130_fd_sc_hd__nor2_4
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21498__A2 _21492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22695__A1 _21528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14562_ _14280_/A _14562_/B _14561_/X VGND VGND VPWR VPWR _14562_/X sky130_fd_sc_hd__and3_4
XPHY_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22695__B2 _22691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11774_ _11833_/A _11774_/B VGND VGND VPWR VPWR _11774_/X sky130_fd_sc_hd__or2_4
XPHY_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _11903_/X _16301_/B VGND VGND VPWR VPWR _16301_/X sky130_fd_sc_hd__or2_4
XFILLER_13_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13535_/A _13447_/B VGND VGND VPWR VPWR _13513_/X sky130_fd_sc_hd__or2_4
X_17281_ _14483_/Y _17019_/X _17026_/X _17280_/X VGND VGND VPWR VPWR _17302_/B sky130_fd_sc_hd__o22a_4
X_14493_ _12401_/A _14493_/B _14492_/X VGND VGND VPWR VPWR _14493_/X sky130_fd_sc_hd__and3_4
XANTENNA__20170__A2 IRQ[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19020_ _19020_/A VGND VGND VPWR VPWR _19020_/Y sky130_fd_sc_hd__inv_2
X_16232_ _16220_/A _16230_/X _16232_/C VGND VGND VPWR VPWR _16236_/B sky130_fd_sc_hd__and3_4
X_13444_ _13467_/A _13444_/B _13444_/C VGND VGND VPWR VPWR _13445_/C sky130_fd_sc_hd__and3_4
XFILLER_127_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16163_ _13413_/A VGND VGND VPWR VPWR _16163_/X sky130_fd_sc_hd__buf_2
X_13375_ _13375_/A _13294_/B VGND VGND VPWR VPWR _13376_/C sky130_fd_sc_hd__or2_4
XFILLER_166_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15114_ _14841_/A _15114_/B _15113_/X VGND VGND VPWR VPWR _15115_/C sky130_fd_sc_hd__and3_4
X_12326_ _11720_/A VGND VGND VPWR VPWR _12327_/A sky130_fd_sc_hd__buf_2
XFILLER_170_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16094_ _16094_/A VGND VGND VPWR VPWR _16144_/A sky130_fd_sc_hd__buf_2
XFILLER_126_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22106__A _22106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19922_ _19438_/A VGND VGND VPWR VPWR _22922_/A sky130_fd_sc_hd__inv_2
X_15045_ _11967_/A _15022_/X _15029_/X _15036_/X _15044_/X VGND VGND VPWR VPWR _15045_/X
+ sky130_fd_sc_hd__a32o_4
X_12257_ _13152_/A _12361_/B VGND VGND VPWR VPWR _12260_/B sky130_fd_sc_hd__or2_4
XANTENNA__16104__A _15971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21958__B1 _12514_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21945__A _21941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19853_ _22687_/B VGND VGND VPWR VPWR _21370_/B sky130_fd_sc_hd__buf_2
X_12188_ _12188_/A VGND VGND VPWR VPWR _13627_/A sky130_fd_sc_hd__buf_2
XFILLER_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15943__A _16011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18804_ _18790_/A VGND VGND VPWR VPWR _18804_/X sky130_fd_sc_hd__buf_2
XANTENNA__21944__A2_N _21943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16996_ _17659_/A _16996_/B VGND VGND VPWR VPWR _16997_/B sky130_fd_sc_hd__or2_4
X_19784_ _19474_/X HRDATA[1] VGND VGND VPWR VPWR _19784_/X sky130_fd_sc_hd__and2_4
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15947_ _15971_/A _15941_/X _15947_/C VGND VGND VPWR VPWR _15947_/X sky130_fd_sc_hd__or3_4
X_18735_ _17108_/X _17246_/Y _18265_/A _18734_/X VGND VGND VPWR VPWR _18735_/X sky130_fd_sc_hd__a211o_4
XFILLER_77_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14559__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13463__A _13431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18666_ _16935_/A _18663_/X _17652_/X _18665_/X VGND VGND VPWR VPWR _18666_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15878_ _13528_/A _15874_/X _15877_/X VGND VGND VPWR VPWR _15879_/C sky130_fd_sc_hd__or3_4
XFILLER_23_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14278__B _14349_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17617_ _17436_/A _17412_/X VGND VGND VPWR VPWR _17617_/Y sky130_fd_sc_hd__nand2_4
X_14829_ _14676_/A _14827_/X _14828_/X VGND VGND VPWR VPWR _14833_/B sky130_fd_sc_hd__and3_4
X_18597_ _16937_/X VGND VGND VPWR VPWR _18597_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14612__A1 _14450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17548_ _17047_/X _17547_/X _17051_/X VGND VGND VPWR VPWR _17548_/X sky130_fd_sc_hd__o21a_4
XFILLER_51_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16924__D _16898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17479_ _17600_/C VGND VGND VPWR VPWR _17490_/C sky130_fd_sc_hd__inv_2
XANTENNA__14294__A _15022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11711__A _12372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19218_ _24312_/Q _19219_/A _19217_/Y VGND VGND VPWR VPWR _24312_/D sky130_fd_sc_hd__o21a_4
X_20490_ _20490_/A VGND VGND VPWR VPWR _20490_/X sky130_fd_sc_hd__buf_2
XFILLER_118_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19149_ _19149_/A _19149_/B VGND VGND VPWR VPWR _19185_/A sky130_fd_sc_hd__and2_4
XFILLER_30_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21110__B2 _21108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22160_ _22158_/X _22159_/X _23450_/Q _22154_/X VGND VGND VPWR VPWR _22160_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15837__B _15837_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21111_ _21104_/A VGND VGND VPWR VPWR _21111_/X sky130_fd_sc_hd__buf_2
XANTENNA__13638__A _15447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22091_ _22090_/X VGND VGND VPWR VPWR _22147_/A sky130_fd_sc_hd__buf_2
XFILLER_114_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21042_ _21042_/A VGND VGND VPWR VPWR _21042_/X sky130_fd_sc_hd__buf_2
XFILLER_119_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21413__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22610__B2 _22605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19325__A _19428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22993_ _22977_/X _18402_/A _22989_/X _22992_/X VGND VGND VPWR VPWR _22993_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22374__B1 _12611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24334__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21177__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13373__A _13392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21944_ _21937_/Y _21943_/X _21811_/X _21943_/X VGND VGND VPWR VPWR _21944_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21590__A _21523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16684__A _16684_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21875_ _21808_/A VGND VGND VPWR VPWR _21875_/X sky130_fd_sc_hd__buf_2
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20918__B _20364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23323_/CLK _21866_/X VGND VGND VPWR VPWR _23614_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _24445_/Q VGND VGND VPWR VPWR _20827_/A sky130_fd_sc_hd__inv_2
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22677__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20688__B1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23545_ _23391_/CLK _23545_/D VGND VGND VPWR VPWR _14724_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20757_ _20703_/X _20756_/X _24384_/Q _20647_/X VGND VGND VPWR VPWR _20757_/X sky130_fd_sc_hd__o22a_4
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11621__A _12473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22429__B2 _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20688_ _20662_/X _20674_/X _20537_/X _20687_/Y VGND VGND VPWR VPWR _20688_/X sky130_fd_sc_hd__a211o_4
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23476_ _23476_/CLK _22096_/X VGND VGND VPWR VPWR _11795_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22427_ _22425_/X _22426_/X _23278_/Q _22421_/X VGND VGND VPWR VPWR _23278_/D sky130_fd_sc_hd__o22a_4
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14932__A _15377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13160_ _13339_/A _13133_/X _13141_/X _13151_/X _13159_/X VGND VGND VPWR VPWR _13160_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_164_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22358_ _22358_/A VGND VGND VPWR VPWR _22366_/A sky130_fd_sc_hd__buf_2
XANTENNA__21652__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12111_ _12027_/X _11633_/X _12076_/X _11609_/X _12110_/X VGND VGND VPWR VPWR _12111_/X
+ sky130_fd_sc_hd__a32o_4
X_13091_ _13091_/A _13091_/B _13090_/X VGND VGND VPWR VPWR _13092_/C sky130_fd_sc_hd__or3_4
X_21309_ _20959_/A VGND VGND VPWR VPWR _21309_/X sky130_fd_sc_hd__buf_2
X_22289_ _22113_/X _22287_/X _23373_/Q _22284_/X VGND VGND VPWR VPWR _23373_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12452__A _15017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12042_ _16695_/A _12039_/X _12042_/C VGND VGND VPWR VPWR _12042_/X sky130_fd_sc_hd__and3_4
X_24028_ _23592_/CLK _21123_/X VGND VGND VPWR VPWR _24028_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18805__B1 _24458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21404__A2 _21398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13267__B _13266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16850_ _14266_/A _16849_/X _14266_/A _16849_/X VGND VGND VPWR VPWR _16850_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22044__A2_N _22043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15801_ _12440_/A _15799_/X _15800_/X VGND VGND VPWR VPWR _15802_/C sky130_fd_sc_hd__and3_4
XFILLER_133_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16781_ _16767_/A _16781_/B _16781_/C VGND VGND VPWR VPWR _16785_/B sky130_fd_sc_hd__and3_4
X_13993_ _12495_/A _14062_/B VGND VGND VPWR VPWR _13993_/X sky130_fd_sc_hd__or2_4
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21168__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13283__A _12559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18520_ _18518_/X _17615_/A _18519_/X VGND VGND VPWR VPWR _18520_/X sky130_fd_sc_hd__a21o_4
X_15732_ _13100_/A _15728_/X _15731_/X VGND VGND VPWR VPWR _15733_/C sky130_fd_sc_hd__or3_4
X_12944_ _12944_/A _12944_/B _12944_/C VGND VGND VPWR VPWR _12945_/C sky130_fd_sc_hd__and3_4
XFILLER_19_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14098__B _23743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18451_ _18356_/X _18449_/X _18396_/X _18450_/X VGND VGND VPWR VPWR _18451_/X sky130_fd_sc_hd__o22a_4
XFILLER_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15663_ _12571_/A _15659_/X _15662_/X VGND VGND VPWR VPWR _15663_/X sky130_fd_sc_hd__or3_4
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12875_ _12875_/A _23945_/Q VGND VGND VPWR VPWR _12877_/B sky130_fd_sc_hd__or2_4
XFILLER_60_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20391__A2 _20381_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17402_ _17402_/A VGND VGND VPWR VPWR _17438_/B sky130_fd_sc_hd__inv_2
XFILLER_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14614_ _14614_/A VGND VGND VPWR VPWR _14841_/A sky130_fd_sc_hd__buf_2
XFILLER_92_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18382_ _17849_/X _18127_/X VGND VGND VPWR VPWR _18382_/X sky130_fd_sc_hd__or2_4
X_11826_ _11705_/X _11824_/X _11825_/X VGND VGND VPWR VPWR _11826_/X sky130_fd_sc_hd__and3_4
XANTENNA__22668__B2 _22662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23925__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15594_ _12337_/A _15594_/B _15594_/C VGND VGND VPWR VPWR _15599_/B sky130_fd_sc_hd__and3_4
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _15251_/A _17333_/B VGND VGND VPWR VPWR _17333_/X sky130_fd_sc_hd__or2_4
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _11681_/A _14537_/X _14544_/X VGND VGND VPWR VPWR _14546_/C sky130_fd_sc_hd__and3_4
XFILLER_14_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11757_ _13392_/A VGND VGND VPWR VPWR _13414_/A sky130_fd_sc_hd__buf_2
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21340__B2 _21338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15003__A _13990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17264_ _17261_/Y _17024_/X _17031_/X _17263_/Y VGND VGND VPWR VPWR _17264_/X sky130_fd_sc_hd__o22a_4
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14476_ _15402_/A _14534_/B VGND VGND VPWR VPWR _14476_/X sky130_fd_sc_hd__or2_4
X_11688_ _12367_/A VGND VGND VPWR VPWR _12630_/A sky130_fd_sc_hd__buf_2
XANTENNA__20844__A _20844_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19003_ _18993_/X _19002_/X _18993_/X _11538_/A VGND VGND VPWR VPWR _24364_/D sky130_fd_sc_hd__a2bb2o_4
X_16215_ _16215_/A _16139_/B VGND VGND VPWR VPWR _16215_/X sky130_fd_sc_hd__or2_4
X_13427_ _13427_/A _23781_/Q VGND VGND VPWR VPWR _13428_/C sky130_fd_sc_hd__or2_4
XFILLER_174_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17195_ _17160_/A _17191_/X _17164_/A _17194_/X VGND VGND VPWR VPWR _17195_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24392__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14842__A _15649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16146_ _16142_/A _23501_/Q VGND VGND VPWR VPWR _16148_/B sky130_fd_sc_hd__or2_4
X_13358_ _13410_/A _13358_/B _13358_/C VGND VGND VPWR VPWR _13358_/X sky130_fd_sc_hd__and3_4
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21643__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14561__B _14633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13458__A _13462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12309_ _12300_/A VGND VGND VPWR VPWR _12745_/A sky130_fd_sc_hd__buf_2
X_16077_ _16049_/A _24110_/Q VGND VGND VPWR VPWR _16078_/C sky130_fd_sc_hd__or2_4
XANTENNA__23305__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13289_ _12904_/A _13285_/X _13289_/C VGND VGND VPWR VPWR _13289_/X sky130_fd_sc_hd__or3_4
XFILLER_143_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12362__A _12362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15376__C _15375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19905_ _19469_/X _19904_/X _17087_/A _19515_/X VGND VGND VPWR VPWR _19905_/Y sky130_fd_sc_hd__a22oi_4
X_15028_ _13985_/A _15028_/B _15027_/X VGND VGND VPWR VPWR _15029_/C sky130_fd_sc_hd__and3_4
XFILLER_29_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16769__A _16683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19836_ _19839_/A _19687_/D _19890_/A _19835_/X VGND VGND VPWR VPWR _19836_/X sky130_fd_sc_hd__o22a_4
XFILLER_96_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15392__B _15454_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23455__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19767_ _19767_/A _19742_/A VGND VGND VPWR VPWR _19767_/X sky130_fd_sc_hd__and2_4
X_16979_ _17721_/A _16978_/X VGND VGND VPWR VPWR _16979_/X sky130_fd_sc_hd__or2_4
XFILLER_83_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13193__A _11668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18718_ _17749_/A VGND VGND VPWR VPWR _18718_/X sky130_fd_sc_hd__buf_2
X_19698_ _17005_/X _19696_/X _21007_/B _19703_/A HRDATA[8] VGND VGND VPWR VPWR _19698_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_64_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19772__A1 _19469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18649_ _17301_/A _18648_/X VGND VGND VPWR VPWR _18649_/Y sky130_fd_sc_hd__nand2_4
XFILLER_52_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13921__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22659__A1 _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22659__B2 _22655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21660_ _21667_/A VGND VGND VPWR VPWR _21660_/X sky130_fd_sc_hd__buf_2
X_20611_ _24230_/Q _20534_/X _20610_/Y VGND VGND VPWR VPWR _20612_/A sky130_fd_sc_hd__o21a_4
X_21591_ _21589_/X _21590_/X _14633_/B _21585_/X VGND VGND VPWR VPWR _21591_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12537__A _12537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16009__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23330_ _23656_/CLK _22340_/X VGND VGND VPWR VPWR _23330_/Q sky130_fd_sc_hd__dfxtp_4
X_20542_ _11556_/A VGND VGND VPWR VPWR _20543_/A sky130_fd_sc_hd__inv_2
XANTENNA__21882__A2 _21875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20473_ _20470_/X _20472_/X _24396_/Q _20429_/X VGND VGND VPWR VPWR _20473_/X sky130_fd_sc_hd__o22a_4
X_23261_ _23229_/CLK _23261_/D VGND VGND VPWR VPWR _13796_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14752__A _12251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22212_ _22176_/A VGND VGND VPWR VPWR _22212_/X sky130_fd_sc_hd__buf_2
X_23192_ _23192_/CLK _23192_/D VGND VGND VPWR VPWR _15260_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_146_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20842__B1 _24093_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22143_ _22141_/X _22135_/X _15607_/B _22142_/X VGND VGND VPWR VPWR _23457_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12272__A _12727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24230__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21585__A _21549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22074_ _22041_/A VGND VGND VPWR VPWR _22074_/X sky130_fd_sc_hd__buf_2
XFILLER_133_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16679__A _16672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21025_ _20533_/A _21024_/X _24085_/Q _20396_/A VGND VGND VPWR VPWR _21025_/X sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_3_1_0_HCLK_A clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18894__A _18837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11616__A _13662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17006__C _17005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22898__B2 _20665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22976_ _22975_/X VGND VGND VPWR VPWR HADDR[12] sky130_fd_sc_hd__inv_2
XFILLER_142_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21927_ _21906_/A VGND VGND VPWR VPWR _21927_/X sky130_fd_sc_hd__buf_2
XFILLER_16_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13831__A _15395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17303__A _14548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12660_ _12962_/A _12649_/X _12660_/C VGND VGND VPWR VPWR _12676_/B sky130_fd_sc_hd__and3_4
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21858_ _21834_/A VGND VGND VPWR VPWR _21858_/X sky130_fd_sc_hd__buf_2
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _17274_/A _11611_/B _11611_/C VGND VGND VPWR VPWR _17062_/D sky130_fd_sc_hd__or3_4
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20644_/X _20808_/X _19235_/A _20758_/X VGND VGND VPWR VPWR _20809_/X sky130_fd_sc_hd__o22a_4
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12625_/A VGND VGND VPWR VPWR _12592_/A sky130_fd_sc_hd__buf_2
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12447__A _12877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21789_ _21572_/X _21784_/X _23649_/Q _21788_/X VGND VGND VPWR VPWR _23649_/D sky130_fd_sc_hd__o22a_4
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _11913_/A _14330_/B _14330_/C VGND VGND VPWR VPWR _14330_/X sky130_fd_sc_hd__and3_4
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23528_ _23656_/CLK _23528_/D VGND VGND VPWR VPWR _23528_/Q sky130_fd_sc_hd__dfxtp_4
X_11542_ _24368_/Q _11542_/B VGND VGND VPWR VPWR _11543_/B sky130_fd_sc_hd__or2_4
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21873__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15758__A _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _14261_/A VGND VGND VPWR VPWR _14263_/B sky130_fd_sc_hd__inv_2
X_23459_ _23908_/CLK _22138_/X VGND VGND VPWR VPWR _15869_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24402__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14662__A _11675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23328__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16000_ _15967_/A _16000_/B VGND VGND VPWR VPWR _16000_/X sky130_fd_sc_hd__or2_4
X_13212_ _13220_/A _23943_/Q VGND VGND VPWR VPWR _13212_/X sky130_fd_sc_hd__or2_4
XANTENNA__21625__A2 _21620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14192_ _14615_/A _14192_/B _14191_/X VGND VGND VPWR VPWR _14192_/X sky130_fd_sc_hd__or3_4
XFILLER_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13143_ _12301_/A VGND VGND VPWR VPWR _13290_/A sky130_fd_sc_hd__buf_2
XFILLER_139_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12182__A _12111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13074_ _13097_/A _23944_/Q VGND VGND VPWR VPWR _13076_/B sky130_fd_sc_hd__or2_4
XANTENNA__23478__CLK _23864_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17951_ _17807_/A _17950_/X VGND VGND VPWR VPWR _17951_/Y sky130_fd_sc_hd__nor2_4
XFILLER_140_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21389__B2 _21388_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16902_ _16902_/A VGND VGND VPWR VPWR _17060_/B sky130_fd_sc_hd__buf_2
X_12025_ _12025_/A _12025_/B VGND VGND VPWR VPWR _12025_/X sky130_fd_sc_hd__or2_4
XFILLER_39_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17882_ _17245_/X VGND VGND VPWR VPWR _17882_/X sky130_fd_sc_hd__buf_2
XANTENNA__12910__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19621_ _19504_/B _19624_/B VGND VGND VPWR VPWR _19622_/B sky130_fd_sc_hd__or2_4
XFILLER_4_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16833_ _12986_/X _16832_/X _13578_/B VGND VGND VPWR VPWR _16833_/X sky130_fd_sc_hd__o21a_4
XFILLER_76_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18006__A1 _17974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16764_ _11704_/X VGND VGND VPWR VPWR _16767_/A sky130_fd_sc_hd__buf_2
X_19552_ _19719_/A VGND VGND VPWR VPWR _19552_/X sky130_fd_sc_hd__buf_2
XFILLER_150_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13976_ _12233_/A _13976_/B _13976_/C VGND VGND VPWR VPWR _13976_/X sky130_fd_sc_hd__and3_4
XFILLER_111_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21010__B1 _22737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15715_ _11864_/A _15714_/X VGND VGND VPWR VPWR _15715_/X sky130_fd_sc_hd__and2_4
X_18503_ _18502_/X VGND VGND VPWR VPWR _18503_/Y sky130_fd_sc_hd__inv_2
X_12927_ _12927_/A VGND VGND VPWR VPWR _12940_/A sky130_fd_sc_hd__buf_2
XFILLER_20_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19483_ _24176_/Q _19481_/X HRDATA[28] _19482_/X VGND VGND VPWR VPWR _19483_/X sky130_fd_sc_hd__o22a_4
X_16695_ _16695_/A _16695_/B _16695_/C VGND VGND VPWR VPWR _16696_/C sky130_fd_sc_hd__and3_4
XFILLER_111_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14837__A _14657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18434_ _24145_/Q _18433_/Y _18403_/B VGND VGND VPWR VPWR _22984_/B sky130_fd_sc_hd__o21a_4
X_15646_ _13923_/A _15646_/B _15646_/C VGND VGND VPWR VPWR _15647_/C sky130_fd_sc_hd__and3_4
X_12858_ _12858_/A VGND VGND VPWR VPWR _12866_/A sky130_fd_sc_hd__buf_2
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11809_ _16053_/A _11777_/X _11809_/C VGND VGND VPWR VPWR _11809_/X sky130_fd_sc_hd__or3_4
X_18365_ _18500_/A _18364_/X VGND VGND VPWR VPWR _18365_/X sky130_fd_sc_hd__or2_4
X_15577_ _14270_/A _15638_/B VGND VGND VPWR VPWR _15577_/X sky130_fd_sc_hd__or2_4
X_12789_ _12800_/A _12789_/B VGND VGND VPWR VPWR _12789_/X sky130_fd_sc_hd__or2_4
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _14845_/Y _17300_/B VGND VGND VPWR VPWR _17316_/X sky130_fd_sc_hd__and2_4
X_14528_ _14540_/A _14526_/X _14527_/X VGND VGND VPWR VPWR _14528_/X sky130_fd_sc_hd__and3_4
XFILLER_109_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18296_ _18095_/X _17522_/X _18292_/X _18168_/X _18295_/Y VGND VGND VPWR VPWR _18296_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21864__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20574__A _22440_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15668__A _12273_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17247_ _18320_/A _17246_/Y VGND VGND VPWR VPWR _17247_/X sky130_fd_sc_hd__and2_4
X_14459_ _12531_/A _14523_/B VGND VGND VPWR VPWR _14459_/X sky130_fd_sc_hd__or2_4
XANTENNA__14572__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24253__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21616__A2 _21613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17178_ _17160_/X _17176_/X _17838_/A _17177_/X VGND VGND VPWR VPWR _17178_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16129_ _16129_/A _16123_/X _16129_/C VGND VGND VPWR VPWR _16129_/X sky130_fd_sc_hd__or3_4
XANTENNA__13188__A _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22577__B1 _14349_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13916__A _13916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12820__A _12834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19819_ _19819_/A _19818_/X VGND VGND VPWR VPWR _19819_/Y sky130_fd_sc_hd__nand2_4
XFILLER_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22830_ _14086_/A _22816_/X _22818_/X _22829_/X VGND VGND VPWR VPWR _22830_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_55_0_HCLK clkbuf_6_27_0_HCLK/X VGND VGND VPWR VPWR _23588_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20749__A HRDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15850__B _15789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22761_ _22760_/Y _22784_/A _22760_/Y _22784_/A VGND VGND VPWR VPWR _22761_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21552__B2 _21549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18219__A _18032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14747__A _14329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24500_ _24471_/CLK _23087_/X HRESETn VGND VGND VPWR VPWR _24500_/Q sky130_fd_sc_hd__dfrtp_4
X_21712_ _21741_/A VGND VGND VPWR VPWR _21727_/A sky130_fd_sc_hd__buf_2
XFILLER_25_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22692_ _22686_/Y _22691_/X _21526_/A _22691_/X VGND VGND VPWR VPWR _23124_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ _24428_/CLK _24431_/D HRESETn VGND VGND VPWR VPWR _24431_/Q sky130_fd_sc_hd__dfrtp_4
X_21643_ _21580_/X _21641_/X _13713_/B _21638_/X VGND VGND VPWR VPWR _21643_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12267__A _13042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24362_ _24357_/CLK _24362_/D HRESETn VGND VGND VPWR VPWR _11536_/A sky130_fd_sc_hd__dfstp_4
X_21574_ _21572_/X _21566_/X _23777_/Q _21573_/X VGND VGND VPWR VPWR _23777_/D sky130_fd_sc_hd__o22a_4
XFILLER_138_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18720__A2 _18717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23313_ _23761_/CLK _22365_/X VGND VGND VPWR VPWR _16766_/B sky130_fd_sc_hd__dfxtp_4
X_20525_ _18238_/X _20469_/X _20514_/X _20524_/Y VGND VGND VPWR VPWR _20525_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15578__A _13687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24293_ _24294_/CLK _24293_/D HRESETn VGND VGND VPWR VPWR _19242_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23244_ _23500_/CLK _23244_/D VGND VGND VPWR VPWR _12303_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_107_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20456_ _20313_/X _20455_/X VGND VGND VPWR VPWR _20456_/Y sky130_fd_sc_hd__nor2_4
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18889__A _17817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17793__A _17792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23175_ _24039_/CLK _22611_/X VGND VGND VPWR VPWR _13216_/B sky130_fd_sc_hd__dfxtp_4
X_20387_ _20343_/X _20386_/X _24336_/Q _20352_/X VGND VGND VPWR VPWR _20387_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22126_ _22125_/X _22123_/X _13013_/B _22118_/X VGND VGND VPWR VPWR _22126_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22568__B1 _15399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13826__A _14329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22057_ _22057_/A VGND VGND VPWR VPWR _22057_/X sky130_fd_sc_hd__buf_2
XFILLER_121_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22032__A2 _22031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12730__A _13164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21008_ _20864_/X _21006_/X _21007_/X HRDATA[8] _20869_/X VGND VGND VPWR VPWR _21008_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17017__B _17017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13830_ _14480_/A _13806_/X _13813_/X _13821_/X _13829_/X VGND VGND VPWR VPWR _13830_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24126__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13761_ _12927_/A _13761_/B VGND VGND VPWR VPWR _13762_/C sky130_fd_sc_hd__or2_4
XFILLER_56_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22959_ _23048_/A VGND VGND VPWR VPWR _22959_/X sky130_fd_sc_hd__buf_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14657__A _14657_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21543__B2 _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15500_ _12616_/A _15492_/X _15499_/X VGND VGND VPWR VPWR _15500_/X sky130_fd_sc_hd__and3_4
X_12712_ _13152_/A _12794_/B VGND VGND VPWR VPWR _12714_/B sky130_fd_sc_hd__or2_4
X_16480_ _16479_/X _16403_/B VGND VGND VPWR VPWR _16480_/X sky130_fd_sc_hd__or2_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13692_ _13692_/A VGND VGND VPWR VPWR _13692_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22874__A _22874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15431_ _15408_/A _15431_/B _15431_/C VGND VGND VPWR VPWR _15435_/B sky130_fd_sc_hd__and3_4
XFILLER_62_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12643_ _12651_/A _12533_/B VGND VGND VPWR VPWR _12643_/X sky130_fd_sc_hd__or2_4
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12177__A _11686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24276__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ _18150_/A _17600_/C VGND VGND VPWR VPWR _18150_/X sky130_fd_sc_hd__or2_4
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15362_ _15362_/A _15362_/B _15361_/X VGND VGND VPWR VPWR _15378_/B sky130_fd_sc_hd__and3_4
X_12574_ _11857_/A _11631_/A _12525_/X _11607_/A _12573_/X VGND VGND VPWR VPWR _12574_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_141_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20394__A _22420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17101_ _17101_/A VGND VGND VPWR VPWR _17101_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14313_ _14448_/A _14313_/B _14313_/C VGND VGND VPWR VPWR _14317_/B sky130_fd_sc_hd__and3_4
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ _19075_/A _19076_/A VGND VGND VPWR VPWR _11525_/X sky130_fd_sc_hd__or2_4
X_18081_ _17850_/X _17828_/X _17986_/X _17840_/X VGND VGND VPWR VPWR _18081_/Y sky130_fd_sc_hd__a22oi_4
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15293_ _14267_/A _23384_/Q VGND VGND VPWR VPWR _15293_/X sky130_fd_sc_hd__or2_4
XANTENNA__12905__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17032_ _17016_/C _11598_/D _17038_/A _17087_/A VGND VGND VPWR VPWR _17033_/A sky130_fd_sc_hd__or4_4
X_14244_ _14623_/A _23103_/Q VGND VGND VPWR VPWR _14244_/X sky130_fd_sc_hd__or2_4
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12624__B _12520_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14175_ _13951_/X _11627_/A _14135_/X _11604_/A _14174_/X VGND VGND VPWR VPWR _14263_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22271__A2 _22244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19672__B1 _20422_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13126_ _13049_/Y _13125_/X VGND VGND VPWR VPWR _13126_/X sky130_fd_sc_hd__or2_4
X_18983_ _18983_/A VGND VGND VPWR VPWR _18983_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18311__B _17522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13057_ _13103_/A _13054_/X _13057_/C VGND VGND VPWR VPWR _13057_/X sky130_fd_sc_hd__and3_4
XFILLER_112_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17934_ _17825_/X _17200_/X _17814_/X _17185_/X VGND VGND VPWR VPWR _17934_/X sky130_fd_sc_hd__o22a_4
XFILLER_87_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22023__A2 _22017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12640__A _12962_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12008_ _12106_/A _23668_/Q VGND VGND VPWR VPWR _12009_/C sky130_fd_sc_hd__or2_4
XANTENNA__21231__B1 _23958_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17419__A2_N _17020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21953__A _21960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17865_ _17849_/X _17855_/X _17856_/X _17864_/Y VGND VGND VPWR VPWR _17865_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20585__A2 _20583_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21782__B2 _21781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19604_ _19563_/X VGND VGND VPWR VPWR _19604_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16816_ _16682_/A _16812_/X _16815_/X VGND VGND VPWR VPWR _16816_/X sky130_fd_sc_hd__or3_4
XFILLER_4_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17796_ _18485_/A VGND VGND VPWR VPWR _17797_/A sky130_fd_sc_hd__inv_2
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19727__B2 _19797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19535_ _19545_/B VGND VGND VPWR VPWR _19848_/A sky130_fd_sc_hd__buf_2
X_13959_ _15029_/A _13954_/X _13959_/C VGND VGND VPWR VPWR _13959_/X sky130_fd_sc_hd__or3_4
X_16747_ _12108_/A _16747_/B _16746_/X VGND VGND VPWR VPWR _16748_/B sky130_fd_sc_hd__or3_4
XANTENNA__14567__A _12530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22731__B1 _14827_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13471__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16678_ _16678_/A _16676_/X _16678_/C VGND VGND VPWR VPWR _16682_/B sky130_fd_sc_hd__and3_4
X_19466_ _19612_/A VGND VGND VPWR VPWR _19859_/A sky130_fd_sc_hd__buf_2
XFILLER_35_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18417_ _17609_/D _18417_/B VGND VGND VPWR VPWR _18417_/X sky130_fd_sc_hd__or2_4
XFILLER_107_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15629_ _15641_/A _15562_/B VGND VGND VPWR VPWR _15629_/X sky130_fd_sc_hd__or2_4
X_19397_ _19396_/X _18112_/X _19396_/X _24237_/Q VGND VGND VPWR VPWR _24237_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21837__A2 _21827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18348_ _17509_/Y _18348_/B VGND VGND VPWR VPWR _18348_/X sky130_fd_sc_hd__or2_4
XANTENNA__23643__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15398__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18279_ _18405_/A _17517_/A VGND VGND VPWR VPWR _18279_/X sky130_fd_sc_hd__or2_4
XANTENNA__12815__A _13563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20310_ _20253_/Y VGND VGND VPWR VPWR _20714_/A sky130_fd_sc_hd__buf_2
XFILLER_163_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21290_ _20770_/A VGND VGND VPWR VPWR _21290_/X sky130_fd_sc_hd__buf_2
XFILLER_162_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20241_ _20241_/A VGND VGND VPWR VPWR _20865_/A sky130_fd_sc_hd__buf_2
XFILLER_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20172_ _20167_/Y _20168_/Y _11547_/X _20171_/Y VGND VGND VPWR VPWR _20172_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22024__A _21991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17118__A _12064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12550__A _12869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22959__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24149__CLK _24306_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23931_ _23515_/CLK _21303_/X VGND VGND VPWR VPWR _14499_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21863__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21773__B2 _21767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23862_ _23862_/CLK _23862_/D VGND VGND VPWR VPWR _23862_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15452__A1 _11854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22813_ _22799_/X VGND VGND VPWR VPWR _22884_/A sky130_fd_sc_hd__buf_2
XFILLER_26_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23793_ _23728_/CLK _21535_/X VGND VGND VPWR VPWR _23793_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14477__A _12504_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13381__A _13399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24299__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22744_ _23086_/A _19325_/X _23086_/B _22743_/Y VGND VGND VPWR VPWR _24129_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22694__A _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14196__B _23775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11613__B _18888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22675_ _22466_/X _22672_/X _13838_/B _22669_/X VGND VGND VPWR VPWR _22675_/X sky130_fd_sc_hd__o22a_4
XFILLER_13_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16692__A _16702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24414_ _23476_/CLK _18874_/X HRESETn VGND VGND VPWR VPWR _24414_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21828__A2 _21827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21626_ _21551_/X _21620_/X _23754_/Q _21624_/X VGND VGND VPWR VPWR _21626_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24345_ _24382_/CLK _24345_/D HRESETn VGND VGND VPWR VPWR _11519_/A sky130_fd_sc_hd__dfstp_4
X_21557_ _21556_/X _21554_/X _23784_/Q _21549_/X VGND VGND VPWR VPWR _23784_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12725__A _12704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20508_ _22117_/A VGND VGND VPWR VPWR _20509_/A sky130_fd_sc_hd__buf_2
X_12290_ _12858_/A VGND VGND VPWR VPWR _13306_/A sky130_fd_sc_hd__buf_2
XFILLER_119_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24276_ _24134_/CLK _24276_/D HRESETn VGND VGND VPWR VPWR _24276_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21488_ _21261_/X _21485_/X _12399_/B _21482_/X VGND VGND VPWR VPWR _23820_/D sky130_fd_sc_hd__o22a_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23227_ _24096_/CLK _23227_/D VGND VGND VPWR VPWR _14469_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22253__A2 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19654__B1 _19888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20439_ _24238_/Q _20420_/X _20438_/Y VGND VGND VPWR VPWR _22110_/A sky130_fd_sc_hd__o21a_4
XFILLER_106_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21461__B1 _14460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23158_ _23862_/CLK _23158_/D VGND VGND VPWR VPWR _23158_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13556__A _13556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22109_ _22108_/X _22099_/X _16274_/B _22106_/X VGND VGND VPWR VPWR _22109_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22005__A2 _22003_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15980_ _16160_/A _15947_/X _15962_/X _15971_/X _15979_/X VGND VGND VPWR VPWR _15980_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12460__A _12288_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23089_ VGND VGND VPWR VPWR _23089_/HI HSIZE[2] sky130_fd_sc_hd__conb_1
X_14931_ _11752_/A _14924_/X _14930_/X VGND VGND VPWR VPWR _14931_/X sky130_fd_sc_hd__or3_4
XANTENNA__21764__B2 _21760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15771__A _15778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14862_ _11618_/A _14862_/B _14862_/C VGND VGND VPWR VPWR _14862_/X sky130_fd_sc_hd__and3_4
X_17650_ _17085_/X _17105_/Y _17248_/X _17647_/Y _17649_/X VGND VGND VPWR VPWR _17650_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_57_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13813_ _15405_/A _13813_/B _13812_/X VGND VGND VPWR VPWR _13813_/X sky130_fd_sc_hd__or3_4
X_16601_ _11984_/X _16577_/X _16584_/X _16592_/X _16600_/X VGND VGND VPWR VPWR _16601_/X
+ sky130_fd_sc_hd__a32o_4
X_17581_ _18118_/B _18116_/B VGND VGND VPWR VPWR _18113_/B sky130_fd_sc_hd__or2_4
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14793_ _15091_/A _14789_/X _14793_/C VGND VGND VPWR VPWR _14793_/X sky130_fd_sc_hd__or3_4
XFILLER_75_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21516__B2 _21510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13291__A _13303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11804__A _11792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19320_ _19319_/X VGND VGND VPWR VPWR _23086_/B sky130_fd_sc_hd__buf_2
XFILLER_73_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16532_ _16531_/X VGND VGND VPWR VPWR _16532_/Y sky130_fd_sc_hd__inv_2
X_13744_ _13744_/A _23326_/Q VGND VGND VPWR VPWR _13744_/X sky130_fd_sc_hd__or2_4
XFILLER_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17196__A1 _17120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12619__B _12619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18393__B1 _17648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16463_ _11715_/A _16394_/B VGND VGND VPWR VPWR _16463_/X sky130_fd_sc_hd__or2_4
X_19251_ _24302_/Q _19251_/B VGND VGND VPWR VPWR _19252_/B sky130_fd_sc_hd__and2_4
XFILLER_32_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13675_ _13675_/A _13772_/B VGND VGND VPWR VPWR _13677_/B sky130_fd_sc_hd__or2_4
XFILLER_143_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18202_ _18202_/A VGND VGND VPWR VPWR _18202_/Y sky130_fd_sc_hd__inv_2
X_15414_ _13655_/A _15471_/B VGND VGND VPWR VPWR _15414_/X sky130_fd_sc_hd__or2_4
X_12626_ _12626_/A VGND VGND VPWR VPWR _12974_/A sky130_fd_sc_hd__buf_2
X_19182_ _19151_/A _19151_/B _19181_/Y VGND VGND VPWR VPWR _19182_/X sky130_fd_sc_hd__o21a_4
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16394_ _16007_/X _16394_/B VGND VGND VPWR VPWR _16394_/X sky130_fd_sc_hd__or2_4
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18133_ _17977_/X _18132_/X _17880_/X VGND VGND VPWR VPWR _18133_/X sky130_fd_sc_hd__o21a_4
X_15345_ _15369_/A _15345_/B _15344_/X VGND VGND VPWR VPWR _15346_/C sky130_fd_sc_hd__or3_4
X_12557_ _12515_/A _12555_/X _12557_/C VGND VGND VPWR VPWR _12563_/B sky130_fd_sc_hd__and3_4
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_4_0_HCLK_A clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18064_ _16932_/X VGND VGND VPWR VPWR _18064_/X sky130_fd_sc_hd__buf_2
X_15276_ _14114_/A _15276_/B _15275_/X VGND VGND VPWR VPWR _15276_/X sky130_fd_sc_hd__and3_4
X_12488_ _12868_/A _12611_/B VGND VGND VPWR VPWR _12488_/X sky130_fd_sc_hd__or2_4
XFILLER_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17015_ _12182_/B VGND VGND VPWR VPWR _17015_/X sky130_fd_sc_hd__buf_2
X_14227_ _14665_/A _23967_/Q VGND VGND VPWR VPWR _14228_/C sky130_fd_sc_hd__or2_4
XFILLER_144_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19418__A _19406_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14850__A _12218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24200__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15665__B _23780_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14158_ _14272_/A _14154_/X _14158_/C VGND VGND VPWR VPWR _14164_/B sky130_fd_sc_hd__and3_4
XANTENNA__13466__A _13443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13109_ _13097_/A _13109_/B VGND VGND VPWR VPWR _13109_/X sky130_fd_sc_hd__or2_4
X_18966_ _24402_/Q VGND VGND VPWR VPWR _18966_/Y sky130_fd_sc_hd__inv_2
X_14089_ _11623_/A _23263_/Q VGND VGND VPWR VPWR _14092_/B sky130_fd_sc_hd__or2_4
XFILLER_86_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17917_ _17917_/A VGND VGND VPWR VPWR _17917_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18897_ _18897_/A VGND VGND VPWR VPWR _18897_/X sky130_fd_sc_hd__buf_2
XFILLER_152_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17848_ _17848_/A VGND VGND VPWR VPWR _17848_/X sky130_fd_sc_hd__buf_2
XFILLER_67_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17779_ _17663_/A _17779_/B _17779_/C _17779_/D VGND VGND VPWR VPWR _17779_/X sky130_fd_sc_hd__or4_4
XANTENNA__14297__A _14297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21507__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11714__A _11714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19518_ _19518_/A VGND VGND VPWR VPWR _19518_/X sky130_fd_sc_hd__buf_2
X_20790_ _20782_/X _20788_/X _19075_/A _20789_/X VGND VGND VPWR VPWR _20790_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17187__A1 _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19449_ HRDATA[0] _19518_/A _19448_/X VGND VGND VPWR VPWR _19450_/A sky130_fd_sc_hd__a21o_4
XFILLER_22_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17401__A _13947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22460_ _22459_/X _22450_/X _23264_/Q _22457_/X VGND VGND VPWR VPWR _23264_/D sky130_fd_sc_hd__o22a_4
XFILLER_33_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21411_ _21302_/X _21405_/X _14477_/B _21409_/X VGND VGND VPWR VPWR _23867_/D sky130_fd_sc_hd__o22a_4
XFILLER_33_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18687__A1 _18413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12545__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22391_ _22146_/X _22390_/X _23295_/Q _22387_/X VGND VGND VPWR VPWR _23295_/D sky130_fd_sc_hd__o22a_4
XFILLER_148_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24130_ _24342_/CLK _24130_/D HRESETn VGND VGND VPWR VPWR _19223_/A sky130_fd_sc_hd__dfrtp_4
X_21342_ _21268_/X _21341_/X _23913_/Q _21338_/X VGND VGND VPWR VPWR _23913_/D sky130_fd_sc_hd__o22a_4
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16162__A2 _11632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15856__A _15894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24061_ _23880_/CLK _24061_/D VGND VGND VPWR VPWR _24061_/Q sky130_fd_sc_hd__dfxtp_4
X_21273_ _20596_/A VGND VGND VPWR VPWR _21273_/X sky130_fd_sc_hd__buf_2
XANTENNA__22235__A2 _22230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23012_ _23007_/X _17688_/A _22989_/X _23011_/X VGND VGND VPWR VPWR _23013_/A sky130_fd_sc_hd__a211o_4
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20224_ _20510_/A VGND VGND VPWR VPWR _20396_/A sky130_fd_sc_hd__buf_2
XANTENNA__21994__B2 _21993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20155_ _20155_/A VGND VGND VPWR VPWR _20155_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22689__A _22722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18886__B _17398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20086_ _20064_/X _18553_/A _20070_/X _20085_/X VGND VGND VPWR VPWR _20087_/A sky130_fd_sc_hd__o22a_4
XFILLER_134_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21746__A1 _21584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16687__A _16687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21746__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23914_ _23467_/CLK _21340_/X VGND VGND VPWR VPWR _12809_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24369__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15591__A _15616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_HCLK_A clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23845_ _23557_/CLK _23845_/D VGND VGND VPWR VPWR _23845_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19998__A _19956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_25_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23776_ _23649_/CLK _21576_/X VGND VGND VPWR VPWR _23776_/Q sky130_fd_sc_hd__dfxtp_4
X_11790_ _12122_/A _11788_/X _11790_/C VGND VGND VPWR VPWR _11790_/X sky130_fd_sc_hd__and3_4
XANTENNA__14000__A _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20937__A _20937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20988_ _24438_/Q VGND VGND VPWR VPWR _20988_/Y sky130_fd_sc_hd__inv_2
XPHY_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12439__B _12584_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22727_ _20860_/A _22722_/X _14396_/B _22726_/X VGND VGND VPWR VPWR _22727_/X sky130_fd_sc_hd__o22a_4
XPHY_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19432__A2_N _18719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18407__A _18407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13460_ _13474_/A _13458_/X _13460_/C VGND VGND VPWR VPWR _13461_/C sky130_fd_sc_hd__and3_4
X_22658_ _22658_/A VGND VGND VPWR VPWR _22658_/X sky130_fd_sc_hd__buf_2
XFILLER_9_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12411_ _12957_/A VGND VGND VPWR VPWR _13542_/A sky130_fd_sc_hd__buf_2
XFILLER_139_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21609_ _21624_/A VGND VGND VPWR VPWR _21617_/A sky130_fd_sc_hd__buf_2
X_13391_ _13413_/A _13391_/B _13390_/X VGND VGND VPWR VPWR _13392_/C sky130_fd_sc_hd__and3_4
XANTENNA__12455__A _12455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22589_ _22622_/A VGND VGND VPWR VPWR _22605_/A sky130_fd_sc_hd__inv_2
XFILLER_51_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15130_ _15257_/A _15130_/B VGND VGND VPWR VPWR _15131_/C sky130_fd_sc_hd__or2_4
XANTENNA__21682__B1 _23718_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12342_ _12339_/X _12340_/X _12341_/X VGND VGND VPWR VPWR _12342_/X sky130_fd_sc_hd__and3_4
X_24328_ _24342_/CLK _24328_/D HRESETn VGND VGND VPWR VPWR _19149_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20672__A _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24314__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15766__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15061_ _14073_/A _15059_/X _15060_/X VGND VGND VPWR VPWR _15065_/B sky130_fd_sc_hd__and3_4
X_12273_ _12273_/A _24076_/Q VGND VGND VPWR VPWR _12274_/C sky130_fd_sc_hd__or2_4
X_24259_ _24137_/CLK _24259_/D HRESETn VGND VGND VPWR VPWR _24259_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14012_ _14012_/A _14011_/X VGND VGND VPWR VPWR _14012_/X sky130_fd_sc_hd__and2_4
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21985__B2 _21950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17981__A _17980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18820_ _14261_/A _18817_/X _11567_/A _18818_/X VGND VGND VPWR VPWR _18820_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12190__A _12190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18751_ _17856_/X _18749_/X _17849_/X _18750_/Y VGND VGND VPWR VPWR _18751_/X sky130_fd_sc_hd__o22a_4
X_15963_ _15957_/A _23694_/Q VGND VGND VPWR VPWR _15965_/B sky130_fd_sc_hd__or2_4
Xclkbuf_7_107_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR _23397_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21737__B2 _21731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17702_ _17702_/A _17473_/A VGND VGND VPWR VPWR _17702_/X sky130_fd_sc_hd__and2_4
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14914_ _14919_/A _14850_/B VGND VGND VPWR VPWR _14914_/X sky130_fd_sc_hd__or2_4
X_15894_ _15894_/A _15894_/B _15894_/C VGND VGND VPWR VPWR _15894_/X sky130_fd_sc_hd__or3_4
XFILLER_23_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18682_ _18627_/X _18630_/X _18627_/X _18630_/X VGND VGND VPWR VPWR _18682_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17633_ _17307_/X _17621_/X _17632_/X VGND VGND VPWR VPWR _18557_/B sky130_fd_sc_hd__or3_4
XFILLER_5_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14845_ _14843_/X VGND VGND VPWR VPWR _14845_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17564_ _18041_/B _18039_/B VGND VGND VPWR VPWR _18035_/B sky130_fd_sc_hd__or2_4
X_14776_ _15076_/A VGND VGND VPWR VPWR _15080_/A sky130_fd_sc_hd__buf_2
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11988_ _12102_/A _21805_/A VGND VGND VPWR VPWR _11991_/B sky130_fd_sc_hd__or2_4
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12349__B _24044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20847__A _20847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19303_ _19235_/B VGND VGND VPWR VPWR _19303_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22162__B2 _22154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16515_ _16164_/X _16438_/B VGND VGND VPWR VPWR _16517_/B sky130_fd_sc_hd__or2_4
X_13727_ _12600_/A VGND VGND VPWR VPWR _13742_/A sky130_fd_sc_hd__buf_2
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14845__A _14843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17495_ _13583_/X _17530_/B VGND VGND VPWR VPWR _17495_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19234_ _19234_/A _19234_/B VGND VGND VPWR VPWR _19235_/B sky130_fd_sc_hd__and2_4
XFILLER_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16446_ _16413_/A _16446_/B VGND VGND VPWR VPWR _16446_/X sky130_fd_sc_hd__or2_4
X_13658_ _13658_/A _23614_/Q VGND VGND VPWR VPWR _13658_/X sky130_fd_sc_hd__or2_4
XANTENNA__24452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12609_ _12625_/A VGND VGND VPWR VPWR _12610_/A sky130_fd_sc_hd__buf_2
XFILLER_157_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16377_ _16370_/X _16373_/X _16377_/C VGND VGND VPWR VPWR _16377_/X sky130_fd_sc_hd__or3_4
X_19165_ _19160_/B VGND VGND VPWR VPWR _19165_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13589_ _13589_/A VGND VGND VPWR VPWR _14292_/A sky130_fd_sc_hd__buf_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21673__B1 _23724_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15328_ _15328_/A _15264_/B VGND VGND VPWR VPWR _15328_/X sky130_fd_sc_hd__or2_4
X_18116_ _18377_/A _18116_/B VGND VGND VPWR VPWR _18119_/C sky130_fd_sc_hd__nor2_4
XFILLER_172_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19096_ _18957_/X VGND VGND VPWR VPWR _19096_/X sky130_fd_sc_hd__buf_2
XANTENNA__15676__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19618__B1 HRDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15259_ _11869_/A _15259_/B _15259_/C VGND VGND VPWR VPWR _15259_/X sky130_fd_sc_hd__or3_4
X_18047_ _17227_/X _18044_/Y _17849_/A _18046_/Y VGND VGND VPWR VPWR _18047_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22217__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14580__A _14301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15395__B _15458_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21976__A1 _21865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13196__A _13205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21976__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11709__A _13866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19998_ _19956_/A VGND VGND VPWR VPWR _19998_/X sky130_fd_sc_hd__buf_2
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18949_ _18949_/A _18949_/B VGND VGND VPWR VPWR _18950_/A sky130_fd_sc_hd__and2_4
XFILLER_101_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21728__B2 _21724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13924__A _14390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21960_ _21960_/A VGND VGND VPWR VPWR _21960_/X sky130_fd_sc_hd__buf_2
XFILLER_67_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20911_ _20695_/X _20902_/Y _20909_/X _20910_/Y _20714_/X VGND VGND VPWR VPWR _20911_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_67_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21891_ _21906_/A VGND VGND VPWR VPWR _21899_/A sky130_fd_sc_hd__buf_2
X_23630_ _24078_/CLK _21828_/X VGND VGND VPWR VPWR _16057_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20842_ _20772_/X _20841_/X _24093_/Q _20746_/X VGND VGND VPWR VPWR _20842_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23561_ _23561_/CLK _21961_/X VGND VGND VPWR VPWR _23561_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20773_ _20895_/A VGND VGND VPWR VPWR _20773_/X sky130_fd_sc_hd__buf_2
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14755__A _12299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21900__B2 _21899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22512_ _22505_/A VGND VGND VPWR VPWR _22512_/X sky130_fd_sc_hd__buf_2
XFILLER_50_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23492_ _23303_/CLK _23492_/D VGND VGND VPWR VPWR _15701_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22972__A _22910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22443_ _22442_/X _22438_/X _23271_/Q _22433_/X VGND VGND VPWR VPWR _23271_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12275__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24122__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22374_ _22117_/X _22369_/X _12611_/B _22373_/X VGND VGND VPWR VPWR _23307_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24113_ _23889_/CLK _24113_/D VGND VGND VPWR VPWR _24113_/Q sky130_fd_sc_hd__dfxtp_4
X_21325_ _21317_/Y _21324_/X _21241_/X _21324_/X VGND VGND VPWR VPWR _21325_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15586__A _13866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24487__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24044_ _24012_/CLK _24044_/D VGND VGND VPWR VPWR _24044_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21256_ _20441_/A VGND VGND VPWR VPWR _21256_/X sky130_fd_sc_hd__buf_2
XFILLER_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20207_ _18777_/X _20079_/X _20206_/Y _19951_/X VGND VGND VPWR VPWR _20207_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18832__A1 _16866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21187_ _21202_/A VGND VGND VPWR VPWR _21195_/A sky130_fd_sc_hd__buf_2
XFILLER_133_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20138_ _11561_/X _20136_/X _20137_/Y VGND VGND VPWR VPWR _20138_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22212__A _22176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21719__B2 _21717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12960_ _12670_/A _12960_/B _12960_/C VGND VGND VPWR VPWR _12961_/C sky130_fd_sc_hd__and3_4
X_20069_ _20069_/A VGND VGND VPWR VPWR _20069_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14649__B _14649_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11911_ _12233_/A VGND VGND VPWR VPWR _11912_/A sky130_fd_sc_hd__buf_2
XFILLER_85_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22392__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12891_ _12891_/A _23145_/Q VGND VGND VPWR VPWR _12891_/X sky130_fd_sc_hd__or2_4
X_14630_ _14630_/A VGND VGND VPWR VPWR _14840_/A sky130_fd_sc_hd__buf_2
X_23828_ _23668_/CLK _23828_/D VGND VGND VPWR VPWR _23828_/Q sky130_fd_sc_hd__dfxtp_4
X_11842_ _11772_/X VGND VGND VPWR VPWR _12167_/A sky130_fd_sc_hd__buf_2
XPHY_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23043__A _23043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14561_ _14270_/A _14633_/B VGND VGND VPWR VPWR _14561_/X sky130_fd_sc_hd__or2_4
XPHY_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23759_ _23662_/CLK _23759_/D VGND VGND VPWR VPWR _16253_/B sky130_fd_sc_hd__dfxtp_4
X_11773_ _11772_/X VGND VGND VPWR VPWR _11833_/A sky130_fd_sc_hd__buf_2
XFILLER_26_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22695__A2 _22694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _13534_/A _13512_/B VGND VGND VPWR VPWR _13514_/B sky130_fd_sc_hd__or2_4
X_16300_ _11889_/X _16300_/B VGND VGND VPWR VPWR _16300_/X sky130_fd_sc_hd__or2_4
XPHY_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17280_ _17280_/A _17280_/B VGND VGND VPWR VPWR _17280_/X sky130_fd_sc_hd__or2_4
XPHY_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14517_/A _23771_/Q VGND VGND VPWR VPWR _14492_/X sky130_fd_sc_hd__or2_4
X_16231_ _16231_/A _24109_/Q VGND VGND VPWR VPWR _16232_/C sky130_fd_sc_hd__or2_4
X_13443_ _13443_/A _23557_/Q VGND VGND VPWR VPWR _13444_/C sky130_fd_sc_hd__or2_4
XANTENNA__15582__B1 _11606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12185__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16162_ _11858_/X _11632_/X _16131_/X _11608_/X _16161_/X VGND VGND VPWR VPWR _16162_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_142_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13374_ _13374_/A _23686_/Q VGND VGND VPWR VPWR _13376_/B sky130_fd_sc_hd__or2_4
XANTENNA__17695__B _17501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15113_ _15091_/A _15113_/B _15113_/C VGND VGND VPWR VPWR _15113_/X sky130_fd_sc_hd__or3_4
XFILLER_155_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12325_ _12827_/A _12193_/B VGND VGND VPWR VPWR _12333_/B sky130_fd_sc_hd__or2_4
X_16093_ _13467_/A VGND VGND VPWR VPWR _16094_/A sky130_fd_sc_hd__buf_2
XFILLER_5_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19921_ _19920_/X VGND VGND VPWR VPWR _19921_/X sky130_fd_sc_hd__buf_2
X_15044_ _11625_/A _15044_/B VGND VGND VPWR VPWR _15044_/X sky130_fd_sc_hd__and2_4
XFILLER_141_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12256_ _15439_/A VGND VGND VPWR VPWR _13152_/A sky130_fd_sc_hd__buf_2
XANTENNA__13728__B _13624_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12632__B _12632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21958__B2 _21957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19852_ _19852_/A VGND VGND VPWR VPWR _22687_/B sky130_fd_sc_hd__buf_2
XANTENNA__18823__A1 _17272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12187_ _13045_/A VGND VGND VPWR VPWR _12571_/A sky130_fd_sc_hd__buf_2
XFILLER_110_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18803_ _18796_/A VGND VGND VPWR VPWR _18803_/X sky130_fd_sc_hd__buf_2
XFILLER_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19783_ HRDATA[17] VGND VGND VPWR VPWR _20598_/B sky130_fd_sc_hd__buf_2
XANTENNA__22122__A _20558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16995_ _17660_/A _16995_/B VGND VGND VPWR VPWR _16996_/B sky130_fd_sc_hd__or2_4
XFILLER_62_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18734_ _17075_/X _18734_/B VGND VGND VPWR VPWR _18734_/X sky130_fd_sc_hd__and2_4
X_15946_ _15993_/A _15946_/B _15946_/C VGND VGND VPWR VPWR _15947_/C sky130_fd_sc_hd__and3_4
XFILLER_110_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16120__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24352__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18665_ _17746_/X _18664_/X _17746_/X _18664_/X VGND VGND VPWR VPWR _18665_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15877_ _13547_/A _15877_/B _15876_/X VGND VGND VPWR VPWR _15877_/X sky130_fd_sc_hd__and3_4
XFILLER_64_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17616_ _17636_/A _17616_/B VGND VGND VPWR VPWR _17637_/C sky130_fd_sc_hd__nor2_4
XFILLER_91_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14828_ _14823_/A _14758_/B VGND VGND VPWR VPWR _14828_/X sky130_fd_sc_hd__or2_4
X_18596_ _17737_/X _18595_/X _17737_/X _18595_/X VGND VGND VPWR VPWR _18596_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17547_ _17274_/A _17035_/A VGND VGND VPWR VPWR _17547_/X sky130_fd_sc_hd__and2_4
XANTENNA__14575__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14759_ _11877_/A _14757_/X _14758_/X VGND VGND VPWR VPWR _14759_/X sky130_fd_sc_hd__and3_4
XFILLER_20_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17478_ _18154_/B _17478_/B VGND VGND VPWR VPWR _17600_/C sky130_fd_sc_hd__or2_4
XFILLER_165_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19217_ _19133_/X VGND VGND VPWR VPWR _19217_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16429_ _16409_/A _16429_/B VGND VGND VPWR VPWR _16429_/X sky130_fd_sc_hd__or2_4
XANTENNA__12095__A _12064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16790__A _16647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19148_ _19148_/A _19148_/B VGND VGND VPWR VPWR _19149_/B sky130_fd_sc_hd__and2_4
XFILLER_30_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21110__A2 _21104_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13919__A _14385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19079_ _18960_/X VGND VGND VPWR VPWR _19079_/X sky130_fd_sc_hd__buf_2
X_21110_ _20633_/X _21104_/X _24037_/Q _21108_/X VGND VGND VPWR VPWR _21110_/X sky130_fd_sc_hd__o22a_4
XFILLER_172_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22090_ _22090_/A _22173_/B _21320_/C _21030_/A VGND VGND VPWR VPWR _22090_/X sky130_fd_sc_hd__or4_4
XANTENNA__12542__B _12647_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21949__B2 _21943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21041_ _20378_/X _21038_/X _24081_/Q _21035_/X VGND VGND VPWR VPWR _21041_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18814__A1 _15916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22610__A2 _22608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16030__A _16047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20909__C1 _20908_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22992_ _22978_/X _22990_/X _22992_/C VGND VGND VPWR VPWR _22992_/X sky130_fd_sc_hd__and3_4
XANTENNA__22967__A _18525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21177__A2 _21176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22374__B2 _22373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14469__B _14469_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21943_ _21950_/A VGND VGND VPWR VPWR _21943_/X sky130_fd_sc_hd__buf_2
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21874_ _21304_/A VGND VGND VPWR VPWR _21874_/X sky130_fd_sc_hd__buf_2
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22126__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23678_/CLK _23613_/D VGND VGND VPWR VPWR _23613_/Q sky130_fd_sc_hd__dfxtp_4
X_20825_ _20825_/A _20316_/X VGND VGND VPWR VPWR _20825_/Y sky130_fd_sc_hd__nand2_4
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14485__A _12362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20688__A1 _20662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23727__CLK _23246_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23544_ _23544_/CLK _23544_/D VGND VGND VPWR VPWR _15343_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20756_ _24416_/Q _20645_/X _24448_/Q _20704_/X VGND VGND VPWR VPWR _20756_/X sky130_fd_sc_hd__o22a_4
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17796__A _18485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22429__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23475_ _23475_/CLK _23475_/D VGND VGND VPWR VPWR _12136_/B sky130_fd_sc_hd__dfxtp_4
X_20687_ _20686_/X VGND VGND VPWR VPWR _20687_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22426_ _22438_/A VGND VGND VPWR VPWR _22426_/X sky130_fd_sc_hd__buf_2
XANTENNA__21637__B1 _23746_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23877__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21111__A _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13829__A _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22357_ _22357_/A VGND VGND VPWR VPWR _22358_/A sky130_fd_sc_hd__inv_2
XFILLER_163_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12110_ _12077_/X _12085_/X _12092_/X _12101_/X _12109_/X VGND VGND VPWR VPWR _12110_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_152_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21308_ _21307_/X _21305_/X _14727_/B _21300_/X VGND VGND VPWR VPWR _21308_/X sky130_fd_sc_hd__o22a_4
XFILLER_163_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13090_ _13090_/A _13090_/B _13089_/X VGND VGND VPWR VPWR _13090_/X sky130_fd_sc_hd__and3_4
XFILLER_124_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22288_ _22110_/X _22287_/X _23374_/Q _22284_/X VGND VGND VPWR VPWR _23374_/D sky130_fd_sc_hd__o22a_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24027_ _23592_/CLK _24027_/D VGND VGND VPWR VPWR _24027_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_46_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12041_ _12041_/A _23763_/Q VGND VGND VPWR VPWR _12042_/C sky130_fd_sc_hd__or2_4
X_21239_ _21264_/A VGND VGND VPWR VPWR _21239_/X sky130_fd_sc_hd__buf_2
XFILLER_78_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18805__A1 _17156_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23038__A _23043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13564__A _13564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15800_ _12860_/A _15800_/B VGND VGND VPWR VPWR _15800_/X sky130_fd_sc_hd__or2_4
XFILLER_59_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17036__A _18782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16780_ _16757_/X _24017_/Q VGND VGND VPWR VPWR _16781_/C sky130_fd_sc_hd__or2_4
X_13992_ _12468_/A _13990_/X _13991_/X VGND VGND VPWR VPWR _13996_/B sky130_fd_sc_hd__and3_4
XANTENNA__21168__A2 _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22877__A _20665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22365__B2 _22359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12943_ _12943_/A _23561_/Q VGND VGND VPWR VPWR _12944_/C sky130_fd_sc_hd__or2_4
X_15731_ _12778_/X _15729_/X _15730_/X VGND VGND VPWR VPWR _15731_/X sky130_fd_sc_hd__and3_4
XFILLER_19_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18450_ _17767_/C _17714_/X _17767_/C _17714_/X VGND VGND VPWR VPWR _18450_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12874_ _12874_/A _12874_/B _12874_/C VGND VGND VPWR VPWR _12874_/X sky130_fd_sc_hd__or3_4
X_15662_ _12722_/A _15660_/X _15662_/C VGND VGND VPWR VPWR _15662_/X sky130_fd_sc_hd__and3_4
X_17401_ _13947_/X _17402_/A VGND VGND VPWR VPWR _17401_/X sky130_fd_sc_hd__or2_4
XFILLER_57_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14613_ _11854_/A _11628_/A _14582_/X _11605_/A _14612_/X VGND VGND VPWR VPWR _14613_/X
+ sky130_fd_sc_hd__a32o_4
X_11825_ _12156_/A _23860_/Q VGND VGND VPWR VPWR _11825_/X sky130_fd_sc_hd__or2_4
X_18381_ _17810_/X _18122_/Y VGND VGND VPWR VPWR _18381_/X sky130_fd_sc_hd__or2_4
X_15593_ _15620_/A _23777_/Q VGND VGND VPWR VPWR _15594_/C sky130_fd_sc_hd__or2_4
XANTENNA__14395__A _11781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12908__A _12510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11812__A _11812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _13756_/A _14544_/B _14543_/X VGND VGND VPWR VPWR _14544_/X sky130_fd_sc_hd__or3_4
XFILLER_109_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17332_ _15252_/X _17332_/B VGND VGND VPWR VPWR _17623_/A sky130_fd_sc_hd__or2_4
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11755_/X VGND VGND VPWR VPWR _13392_/A sky130_fd_sc_hd__buf_2
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21340__A2 _21334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12627__B _23467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _12470_/A _14473_/X _14475_/C VGND VGND VPWR VPWR _14475_/X sky130_fd_sc_hd__and3_4
X_17263_ _17047_/X _17262_/X _17051_/X VGND VGND VPWR VPWR _17263_/Y sky130_fd_sc_hd__o21ai_4
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _13865_/A VGND VGND VPWR VPWR _12367_/A sky130_fd_sc_hd__buf_2
X_19002_ _18987_/X _19000_/Y _19001_/Y _18990_/X VGND VGND VPWR VPWR _19002_/X sky130_fd_sc_hd__o22a_4
X_16214_ _16214_/A _16210_/X _16214_/C VGND VGND VPWR VPWR _16222_/B sky130_fd_sc_hd__or3_4
X_13426_ _13455_/A _13500_/B VGND VGND VPWR VPWR _13426_/X sky130_fd_sc_hd__or2_4
X_17194_ _16383_/X _17192_/X _14701_/Y _17193_/X VGND VGND VPWR VPWR _17194_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22117__A _22117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16145_ _16145_/A _16145_/B _16145_/C VGND VGND VPWR VPWR _16145_/X sky130_fd_sc_hd__or3_4
XANTENNA__21021__A _20977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13357_ _13385_/A _23782_/Q VGND VGND VPWR VPWR _13358_/C sky130_fd_sc_hd__or2_4
XFILLER_170_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20300__B1 _20225_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12308_ _13306_/A _12308_/B _12307_/X VGND VGND VPWR VPWR _12308_/X sky130_fd_sc_hd__or3_4
X_16076_ _16048_/A _16076_/B VGND VGND VPWR VPWR _16078_/B sky130_fd_sc_hd__or2_4
X_13288_ _13318_/A _13288_/B _13288_/C VGND VGND VPWR VPWR _13289_/C sky130_fd_sc_hd__and3_4
XANTENNA__20860__A _20860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19904_ _19576_/X _19902_/X _19903_/X _19603_/X _19642_/Y VGND VGND VPWR VPWR _19904_/X
+ sky130_fd_sc_hd__a32o_4
X_15027_ _13964_/A _23413_/Q VGND VGND VPWR VPWR _15027_/X sky130_fd_sc_hd__or2_4
X_12239_ _12239_/A VGND VGND VPWR VPWR _12240_/A sky130_fd_sc_hd__buf_2
XFILLER_64_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18330__A _16941_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19835_ _19809_/A _19830_/X _19834_/X VGND VGND VPWR VPWR _19835_/X sky130_fd_sc_hd__and3_4
XANTENNA__13474__A _13474_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19766_ _19528_/A _19663_/Y _19815_/B _19765_/X VGND VGND VPWR VPWR _19787_/B sky130_fd_sc_hd__and4_4
X_16978_ _17726_/A _16977_/X VGND VGND VPWR VPWR _16978_/X sky130_fd_sc_hd__or2_4
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21691__A _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18717_ _18506_/X _18709_/X _18710_/Y _18712_/X _18716_/Y VGND VGND VPWR VPWR _18717_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24182__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15929_ _15929_/A VGND VGND VPWR VPWR _15929_/Y sky130_fd_sc_hd__inv_2
X_19697_ HRDATA[24] VGND VGND VPWR VPWR _21007_/B sky130_fd_sc_hd__buf_2
XFILLER_65_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18648_ _17980_/X _18673_/B _17631_/B _17805_/X _18600_/X VGND VGND VPWR VPWR _18648_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_52_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13921__B _13838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22659__A2 _22658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18579_ _18578_/X VGND VGND VPWR VPWR _18579_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12818__A _13562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20610_ _20438_/A _20610_/B VGND VGND VPWR VPWR _20610_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__11722__A _15606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21590_ _21523_/A VGND VGND VPWR VPWR _21590_/X sky130_fd_sc_hd__buf_2
X_20541_ _20541_/A _20318_/B VGND VGND VPWR VPWR _20541_/Y sky130_fd_sc_hd__nand2_4
XFILLER_119_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18505__A _17648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23260_ _24096_/CLK _23260_/D VGND VGND VPWR VPWR _14337_/B sky130_fd_sc_hd__dfxtp_4
X_20472_ _24428_/Q _20427_/X _24460_/Q _20471_/X VGND VGND VPWR VPWR _20472_/X sky130_fd_sc_hd__o22a_4
XFILLER_158_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_15_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR _23379_/CLK sky130_fd_sc_hd__clkbuf_1
X_22211_ _22151_/X _22208_/X _13842_/B _22205_/X VGND VGND VPWR VPWR _22211_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22292__B1 _23371_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21095__B2 _21094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13649__A _12288_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23191_ _23192_/CLK _22583_/X VGND VGND VPWR VPWR _15129_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12553__A _12515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_78_0_HCLK clkbuf_7_79_0_HCLK/A VGND VGND VPWR VPWR _23641_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15849__A1 _11857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11583__A1 _24466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22142_ _22118_/A VGND VGND VPWR VPWR _22142_/X sky130_fd_sc_hd__buf_2
XANTENNA__20842__B2 _20746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15864__A _13564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22073_ _21860_/X _22067_/X _23488_/Q _22071_/X VGND VGND VPWR VPWR _22073_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18240__A _18064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18799__B1 _24462_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22595__B2 _22591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21024_ _21024_/A VGND VGND VPWR VPWR _21024_/X sky130_fd_sc_hd__buf_2
XFILLER_59_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13384__A _13384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21375__A2_N _21374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14199__B _24031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22975_ _22946_/X _18478_/A _22959_/X _22974_/X VGND VGND VPWR VPWR _22975_/X sky130_fd_sc_hd__a211o_4
XFILLER_167_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21926_ _21867_/X _21923_/X _13897_/B _21920_/X VGND VGND VPWR VPWR _23581_/D sky130_fd_sc_hd__o22a_4
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14927__B _14859_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21857_ _20745_/A VGND VGND VPWR VPWR _21857_/X sky130_fd_sc_hd__buf_2
XANTENNA__12728__A _13279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11632__A _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11609_/X VGND VGND VPWR VPWR _11610_/X sky130_fd_sc_hd__buf_2
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _20703_/X _20807_/X _24382_/Q _20647_/X VGND VGND VPWR VPWR _20808_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15104__A _15080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12590_ _12970_/A _23371_/Q VGND VGND VPWR VPWR _12590_/X sky130_fd_sc_hd__or2_4
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21788_ _21774_/A VGND VGND VPWR VPWR _21788_/X sky130_fd_sc_hd__buf_2
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23527_ _23723_/CLK _22013_/X VGND VGND VPWR VPWR _23527_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _24367_/Q _11541_/B VGND VGND VPWR VPWR _11542_/B sky130_fd_sc_hd__or2_4
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20739_ _20738_/X VGND VGND VPWR VPWR _20739_/Y sky130_fd_sc_hd__inv_2
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _11666_/X _14223_/X _14259_/X VGND VGND VPWR VPWR _14261_/A sky130_fd_sc_hd__and3_4
X_23458_ _23908_/CLK _23458_/D VGND VGND VPWR VPWR _15474_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13211_ _11682_/A _13211_/B _13210_/X VGND VGND VPWR VPWR _13229_/B sky130_fd_sc_hd__and3_4
XANTENNA__13559__A _13547_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22409_ _22421_/A VGND VGND VPWR VPWR _22409_/X sky130_fd_sc_hd__buf_2
XFILLER_125_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14191_ _14191_/A _14188_/X _14190_/X VGND VGND VPWR VPWR _14191_/X sky130_fd_sc_hd__and3_4
XFILLER_164_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12463__A _12863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24055__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23389_ _23582_/CLK _23389_/D VGND VGND VPWR VPWR _13841_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_13_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11574__A1 _24456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13142_ _13045_/A VGND VGND VPWR VPWR _13338_/A sky130_fd_sc_hd__buf_2
XFILLER_13_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13073_ _12977_/A _13062_/X _13073_/C VGND VGND VPWR VPWR _13093_/B sky130_fd_sc_hd__and3_4
XFILLER_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17950_ _17875_/X _17949_/X _17883_/X VGND VGND VPWR VPWR _17950_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18150__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21389__A2 _21384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16901_ _16901_/A VGND VGND VPWR VPWR _16902_/A sky130_fd_sc_hd__inv_2
X_12024_ _12024_/A _12020_/X VGND VGND VPWR VPWR _12025_/B sky130_fd_sc_hd__and2_4
XANTENNA__15493__B _15493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17881_ _17877_/X _17879_/X _17880_/X VGND VGND VPWR VPWR _17881_/X sky130_fd_sc_hd__o21a_4
X_19620_ _19624_/A VGND VGND VPWR VPWR _19687_/A sky130_fd_sc_hd__buf_2
XFILLER_116_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16832_ _16832_/A _16831_/X VGND VGND VPWR VPWR _16832_/X sky130_fd_sc_hd__and2_4
XFILLER_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19551_ _19516_/X _19520_/Y _19521_/Y _19550_/X VGND VGND VPWR VPWR _19551_/X sky130_fd_sc_hd__o22a_4
XFILLER_93_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16763_ _16647_/A _16761_/X _16763_/C VGND VGND VPWR VPWR _16768_/B sky130_fd_sc_hd__and3_4
X_13975_ _13606_/A _23584_/Q VGND VGND VPWR VPWR _13976_/C sky130_fd_sc_hd__or2_4
XANTENNA__24225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18502_ _18111_/A _18365_/X _18500_/Y _18026_/X _22966_/B VGND VGND VPWR VPWR _18502_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17214__B1 _13947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15714_ _11872_/A _15710_/X _15714_/C VGND VGND VPWR VPWR _15714_/X sky130_fd_sc_hd__or3_4
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12926_ _12951_/A _24041_/Q VGND VGND VPWR VPWR _12929_/B sky130_fd_sc_hd__or2_4
X_19482_ _19452_/X VGND VGND VPWR VPWR _19482_/X sky130_fd_sc_hd__buf_2
X_16694_ _16691_/A _23761_/Q VGND VGND VPWR VPWR _16695_/C sky130_fd_sc_hd__or2_4
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18433_ _18433_/A VGND VGND VPWR VPWR _18433_/Y sky130_fd_sc_hd__inv_2
X_15645_ _13885_/A _23649_/Q VGND VGND VPWR VPWR _15646_/C sky130_fd_sc_hd__or2_4
X_12857_ _12857_/A _12849_/X _12857_/C VGND VGND VPWR VPWR _12857_/X sky130_fd_sc_hd__or3_4
XANTENNA__12638__A _12944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15014__A _13981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11808_ _11786_/X _11797_/X _11807_/X VGND VGND VPWR VPWR _11809_/C sky130_fd_sc_hd__and3_4
X_18364_ _18533_/A _18533_/B VGND VGND VPWR VPWR _18364_/X sky130_fd_sc_hd__or2_4
X_12788_ _13415_/A _12771_/X _12787_/X VGND VGND VPWR VPWR _12788_/X sky130_fd_sc_hd__and3_4
X_15576_ _12434_/A _23713_/Q VGND VGND VPWR VPWR _15578_/B sky130_fd_sc_hd__or2_4
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22510__B2 _22505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17315_ _18673_/B VGND VGND VPWR VPWR _17315_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15949__A _11917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11739_ _11739_/A VGND VGND VPWR VPWR _13377_/A sky130_fd_sc_hd__buf_2
X_14527_ _14520_/A _14463_/B VGND VGND VPWR VPWR _14527_/X sky130_fd_sc_hd__or2_4
X_18295_ _17527_/D _18294_/X _17533_/Y VGND VGND VPWR VPWR _18295_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__14853__A _12218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17246_ _11610_/X _17243_/X _17245_/X VGND VGND VPWR VPWR _17246_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_174_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14458_ _12461_/A _14454_/X _14458_/C VGND VGND VPWR VPWR _14458_/X sky130_fd_sc_hd__or3_4
XFILLER_128_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13469__A _13441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13409_ _13397_/A _24102_/Q VGND VGND VPWR VPWR _13410_/C sky130_fd_sc_hd__or2_4
XANTENNA__21077__B2 _21042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12373__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14389_ _14509_/A _14387_/X _14388_/X VGND VGND VPWR VPWR _14389_/X sky130_fd_sc_hd__and3_4
X_17177_ _13583_/X _17107_/X _15786_/Y _17074_/X VGND VGND VPWR VPWR _17177_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16128_ _16155_/A _16125_/X _16128_/C VGND VGND VPWR VPWR _16129_/C sky130_fd_sc_hd__and3_4
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23422__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15684__A _12858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16059_ _16035_/A _16059_/B _16059_/C VGND VGND VPWR VPWR _16060_/C sky130_fd_sc_hd__and3_4
XFILLER_142_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22577__B2 _22576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11717__A _16079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20052__A2 _20031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19818_ _19724_/A _19808_/Y _19809_/Y _19817_/X VGND VGND VPWR VPWR _19818_/X sky130_fd_sc_hd__a211o_4
XFILLER_97_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19749_ _19682_/A VGND VGND VPWR VPWR _19749_/X sky130_fd_sc_hd__buf_2
XANTENNA__17205__B1 _17170_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22760_ SYSTICKCLKDIV[4] VGND VGND VPWR VPWR _22760_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21552__A2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14747__B _23417_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21711_ _21705_/Y _21710_/X _21526_/X _21710_/X VGND VGND VPWR VPWR _23700_/D sky130_fd_sc_hd__a2bb2o_4
X_22691_ _22698_/A VGND VGND VPWR VPWR _22691_/X sky130_fd_sc_hd__buf_2
XFILLER_13_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24430_ _24428_/CLK _24430_/D HRESETn VGND VGND VPWR VPWR _24430_/Q sky130_fd_sc_hd__dfrtp_4
X_21642_ _21577_/X _21641_/X _23743_/Q _21638_/X VGND VGND VPWR VPWR _21642_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15859__A _12402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24361_ _24360_/CLK _24361_/D HRESETn VGND VGND VPWR VPWR _11535_/A sky130_fd_sc_hd__dfstp_4
X_21573_ _21549_/A VGND VGND VPWR VPWR _21573_/X sky130_fd_sc_hd__buf_2
XFILLER_36_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23312_ _24080_/CLK _22367_/X VGND VGND VPWR VPWR _16398_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_123_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20524_ _20388_/A _20523_/X VGND VGND VPWR VPWR _20524_/Y sky130_fd_sc_hd__nor2_4
X_24292_ _24292_/CLK _24292_/D HRESETn VGND VGND VPWR VPWR _24292_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22980__A _18472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13379__A _13379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23243_ _24012_/CLK _22506_/X VGND VGND VPWR VPWR _12671_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21068__B2 _21063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20455_ _20754_/A _20454_/X _19154_/A _20761_/A VGND VGND VPWR VPWR _20455_/X sky130_fd_sc_hd__o22a_4
XFILLER_4_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21596__A _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18889__B _18889_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23174_ _24102_/CLK _23174_/D VGND VGND VPWR VPWR _23174_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20386_ _20344_/X _20385_/X _24368_/Q _20269_/X VGND VGND VPWR VPWR _20386_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22125_ _22440_/A VGND VGND VPWR VPWR _22125_/X sky130_fd_sc_hd__buf_2
XFILLER_161_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22568__B2 _22562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22056_ _21831_/X _22053_/X _12293_/B _22050_/X VGND VGND VPWR VPWR _23500_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_7_8_0_HCLK clkbuf_6_4_0_HCLK/X VGND VGND VPWR VPWR _24445_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21007_ _21007_/A _21007_/B VGND VGND VPWR VPWR _21007_/X sky130_fd_sc_hd__or2_4
XANTENNA__20043__A2 _20031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14003__A _14003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13842__A _12198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13760_ _12925_/A _13760_/B VGND VGND VPWR VPWR _13760_/X sky130_fd_sc_hd__or2_4
XFILLER_16_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17314__A _14845_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22958_ _22957_/X VGND VGND VPWR VPWR HADDR[9] sky130_fd_sc_hd__inv_2
XFILLER_56_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21543__A2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21909_ _21909_/A VGND VGND VPWR VPWR _21909_/X sky130_fd_sc_hd__buf_2
X_12711_ _12279_/A _12709_/X _12710_/X VGND VGND VPWR VPWR _12715_/B sky130_fd_sc_hd__and3_4
XFILLER_44_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13691_ _11855_/A _11629_/A _13651_/X _11606_/A _13690_/X VGND VGND VPWR VPWR _13692_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22889_ _22876_/X _22829_/X _14086_/A _22877_/X VGND VGND VPWR VPWR _22889_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12642_ _12587_/A VGND VGND VPWR VPWR _12972_/A sky130_fd_sc_hd__buf_2
X_15430_ _14319_/A _15494_/B VGND VGND VPWR VPWR _15431_/C sky130_fd_sc_hd__or2_4
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ _15321_/A _15361_/B _15360_/X VGND VGND VPWR VPWR _15361_/X sky130_fd_sc_hd__or3_4
X_12573_ _13453_/A _12544_/X _12554_/X _12563_/X _12572_/X VGND VGND VPWR VPWR _12573_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_141_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15769__A _12778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18145__A _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17100_ _17100_/A _17083_/B VGND VGND VPWR VPWR _17101_/A sky130_fd_sc_hd__or2_4
X_14312_ _12485_/A _14388_/B VGND VGND VPWR VPWR _14313_/C sky130_fd_sc_hd__or2_4
XFILLER_12_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11524_ _11524_/A _11524_/B VGND VGND VPWR VPWR _19076_/A sky130_fd_sc_hd__or2_4
XFILLER_54_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15292_ _15269_/A _15290_/X _15291_/X VGND VGND VPWR VPWR _15292_/X sky130_fd_sc_hd__and3_4
X_18080_ _18080_/A VGND VGND VPWR VPWR _18080_/Y sky130_fd_sc_hd__inv_2
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23445__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13289__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17031_ _17031_/A VGND VGND VPWR VPWR _17031_/X sky130_fd_sc_hd__buf_2
X_14243_ _14663_/A _14243_/B _14242_/X VGND VGND VPWR VPWR _14259_/B sky130_fd_sc_hd__and3_4
XANTENNA__12193__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14174_ _14302_/A _14143_/X _14150_/X _14164_/X _14173_/X VGND VGND VPWR VPWR _14174_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19672__A1 _19519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_61_0_HCLK clkbuf_6_30_0_HCLK/X VGND VGND VPWR VPWR _23723_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22008__B1 _12584_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13125_ _12979_/A _13125_/B _13124_/X VGND VGND VPWR VPWR _13125_/X sky130_fd_sc_hd__and3_4
XFILLER_98_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18982_ _18980_/Y _18981_/Y _11542_/B VGND VGND VPWR VPWR _18982_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12921__A _12659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22559__A1 _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22559__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13056_ _13095_/A _23528_/Q VGND VGND VPWR VPWR _13057_/C sky130_fd_sc_hd__or2_4
X_17933_ _17878_/X VGND VGND VPWR VPWR _17933_/X sky130_fd_sc_hd__buf_2
XANTENNA__24406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12007_ _12105_/A _11845_/B VGND VGND VPWR VPWR _12009_/B sky130_fd_sc_hd__or2_4
XANTENNA__21231__B2 _21195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15009__A _13955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17864_ _17864_/A VGND VGND VPWR VPWR _17864_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21782__A2 _21777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19603_ _19895_/A VGND VGND VPWR VPWR _19603_/X sky130_fd_sc_hd__buf_2
XFILLER_94_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16815_ _16646_/A _16813_/X _16814_/X VGND VGND VPWR VPWR _16815_/X sky130_fd_sc_hd__and3_4
XFILLER_66_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22130__A _22118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17795_ _18222_/A _17256_/B VGND VGND VPWR VPWR _17795_/X sky130_fd_sc_hd__and2_4
X_19534_ _19705_/B VGND VGND VPWR VPWR _19545_/B sky130_fd_sc_hd__inv_2
XANTENNA__17224__A _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16746_ _11963_/A _16746_/B _16746_/C VGND VGND VPWR VPWR _16746_/X sky130_fd_sc_hd__and3_4
X_13958_ _13985_/A _13956_/X _13958_/C VGND VGND VPWR VPWR _13959_/C sky130_fd_sc_hd__and3_4
XFILLER_19_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22731__B2 _22726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12909_ _12513_/A _23881_/Q VGND VGND VPWR VPWR _12909_/X sky130_fd_sc_hd__or2_4
X_19465_ _19465_/A VGND VGND VPWR VPWR _19612_/A sky130_fd_sc_hd__inv_2
X_16677_ _16677_/A _24114_/Q VGND VGND VPWR VPWR _16678_/C sky130_fd_sc_hd__or2_4
XANTENNA__12368__A _13251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13889_ _13916_/A _24029_/Q VGND VGND VPWR VPWR _13889_/X sky130_fd_sc_hd__or2_4
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18416_ _17606_/X _18416_/B VGND VGND VPWR VPWR _18417_/B sky130_fd_sc_hd__and2_4
XANTENNA__24220__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15628_ _15612_/A _15628_/B _15627_/X VGND VGND VPWR VPWR _15628_/X sky130_fd_sc_hd__and3_4
X_19396_ _19377_/A VGND VGND VPWR VPWR _19396_/X sky130_fd_sc_hd__buf_2
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15679__A _12702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18347_ _18095_/X _17495_/X _18345_/X _18168_/X _18346_/Y VGND VGND VPWR VPWR _18348_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21298__B2 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15559_ _11886_/A _15559_/B VGND VGND VPWR VPWR _15559_/X sky130_fd_sc_hd__or2_4
XANTENNA__18055__A _18320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14583__A _14278_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19360__B1 _19358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18278_ _18251_/A _23014_/B _18253_/A VGND VGND VPWR VPWR _18278_/X sky130_fd_sc_hd__o21a_4
X_17229_ _17878_/A VGND VGND VPWR VPWR _17229_/X sky130_fd_sc_hd__buf_2
XFILLER_174_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20240_ _19913_/A HRDATA[15] VGND VGND VPWR VPWR _20240_/X sky130_fd_sc_hd__or2_4
XFILLER_66_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22305__A _22291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13927__A _14335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20171_ _24442_/Q IRQ[5] _20169_/Y _20170_/X VGND VGND VPWR VPWR _20171_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__12831__A _13377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21222__B2 _21216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23930_ _24090_/CLK _21306_/X VGND VGND VPWR VPWR _14644_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_96_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21773__A2 _21770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23861_ _23392_/CLK _23861_/D VGND VGND VPWR VPWR _15104_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20981__B1 _15170_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22812_ _17273_/Y _22803_/X VGND VGND VPWR VPWR HWDATA[7] sky130_fd_sc_hd__nor2_4
XANTENNA__13662__A _13662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23792_ _23760_/CLK _23792_/D VGND VGND VPWR VPWR _16395_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22743_ _22736_/X VGND VGND VPWR VPWR _22743_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22674_ _22464_/X _22672_/X _13757_/B _22669_/X VGND VGND VPWR VPWR _22674_/X sky130_fd_sc_hd__o22a_4
XFILLER_41_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24413_ _24445_/CLK _24413_/D HRESETn VGND VGND VPWR VPWR _20825_/A sky130_fd_sc_hd__dfrtp_4
X_21625_ _21548_/X _21620_/X _23755_/Q _21624_/X VGND VGND VPWR VPWR _23755_/D sky130_fd_sc_hd__o22a_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21289__B2 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14493__A _12401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24344_ _24342_/CLK _24344_/D HRESETn VGND VGND VPWR VPWR _11518_/A sky130_fd_sc_hd__dfstp_4
X_21556_ _20575_/A VGND VGND VPWR VPWR _21556_/X sky130_fd_sc_hd__buf_2
XFILLER_126_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20507_ _24235_/Q _20420_/X _20506_/X VGND VGND VPWR VPWR _22117_/A sky130_fd_sc_hd__o21a_4
XFILLER_107_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24275_ _24471_/CLK _24275_/D HRESETn VGND VGND VPWR VPWR _24275_/Q sky130_fd_sc_hd__dfrtp_4
X_21487_ _21259_/X _21485_/X _16224_/B _21482_/X VGND VGND VPWR VPWR _23821_/D sky130_fd_sc_hd__o22a_4
XFILLER_10_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23226_ _23641_/CLK _23226_/D VGND VGND VPWR VPWR _14600_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_107_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20438_ _20438_/A _20438_/B VGND VGND VPWR VPWR _20438_/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22215__A _22208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_48_0_HCLK clkbuf_6_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_48_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13837__A _15405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23157_ _23392_/CLK _23157_/D VGND VGND VPWR VPWR _23157_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21461__B2 _21459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12741__A _12741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20369_ _20344_/X _20368_/X _24369_/Q _20269_/X VGND VGND VPWR VPWR _20369_/X sky130_fd_sc_hd__o22a_4
XFILLER_164_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22108_ _20415_/A VGND VGND VPWR VPWR _22108_/X sky130_fd_sc_hd__buf_2
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23088_ VGND VGND VPWR VPWR _24130_/D _23088_/LO sky130_fd_sc_hd__conb_1
XFILLER_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21213__B2 _21209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14930_ _14925_/X _14927_/X _14929_/X VGND VGND VPWR VPWR _14930_/X sky130_fd_sc_hd__and3_4
X_22039_ _22039_/A _22039_/B _22487_/A _21234_/B VGND VGND VPWR VPWR _22039_/X sky130_fd_sc_hd__or4_4
XANTENNA__21764__A2 _21763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14861_ _14881_/A _14929_/B VGND VGND VPWR VPWR _14862_/C sky130_fd_sc_hd__or2_4
X_16600_ _11867_/X _16600_/B VGND VGND VPWR VPWR _16600_/X sky130_fd_sc_hd__and2_4
XFILLER_29_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13812_ _12470_/A _13812_/B _13812_/C VGND VGND VPWR VPWR _13812_/X sky130_fd_sc_hd__and3_4
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24243__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17580_ _16242_/X _18114_/B VGND VGND VPWR VPWR _18116_/B sky130_fd_sc_hd__and2_4
XANTENNA__13454__A1 _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14792_ _14676_/A _14790_/X _14792_/C VGND VGND VPWR VPWR _14793_/C sky130_fd_sc_hd__and3_4
XANTENNA__14387__B _14387_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21516__A2 _21513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22713__B2 _22712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16531_ _16385_/Y _16525_/A _16526_/A _16530_/Y VGND VGND VPWR VPWR _16531_/X sky130_fd_sc_hd__a211o_4
XFILLER_95_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13743_ _13743_/A _13741_/X _13743_/C VGND VGND VPWR VPWR _13747_/B sky130_fd_sc_hd__and3_4
XFILLER_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12188__A _12188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19590__B1 HRDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19250_ _19250_/A _19250_/B VGND VGND VPWR VPWR _19251_/B sky130_fd_sc_hd__and2_4
X_16462_ _16362_/X _16455_/X _16462_/C VGND VGND VPWR VPWR _16462_/X sky130_fd_sc_hd__or3_4
XFILLER_71_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13674_ _15412_/A _13669_/X _13673_/X VGND VGND VPWR VPWR _13674_/X sky130_fd_sc_hd__or3_4
XFILLER_32_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18201_ _17874_/X _18199_/Y _18200_/X _18090_/X VGND VGND VPWR VPWR _18202_/A sky130_fd_sc_hd__o22a_4
X_15413_ _14325_/A _15470_/B VGND VGND VPWR VPWR _15413_/X sky130_fd_sc_hd__or2_4
X_12625_ _12625_/A VGND VGND VPWR VPWR _12626_/A sky130_fd_sc_hd__buf_2
X_19181_ _19151_/X VGND VGND VPWR VPWR _19181_/Y sky130_fd_sc_hd__inv_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16393_ _15934_/X _16389_/X _16392_/X VGND VGND VPWR VPWR _16393_/X sky130_fd_sc_hd__or3_4
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__A _12923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18132_ _17933_/X _17994_/X _17933_/X _17947_/Y VGND VGND VPWR VPWR _18132_/X sky130_fd_sc_hd__a2bb2o_4
X_12556_ _12514_/A _12669_/B VGND VGND VPWR VPWR _12557_/C sky130_fd_sc_hd__or2_4
X_15344_ _11735_/A _15342_/X _15343_/X VGND VGND VPWR VPWR _15344_/X sky130_fd_sc_hd__and3_4
XFILLER_156_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18063_ _17963_/X _18031_/Y _18033_/X _18062_/X VGND VGND VPWR VPWR _18063_/X sky130_fd_sc_hd__o22a_4
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15011__B _23445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12487_ _12487_/A VGND VGND VPWR VPWR _12868_/A sky130_fd_sc_hd__buf_2
X_15275_ _14131_/A _15333_/B VGND VGND VPWR VPWR _15275_/X sky130_fd_sc_hd__or2_4
XFILLER_172_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18603__A _17594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17014_ _17013_/X VGND VGND VPWR VPWR _17014_/X sky130_fd_sc_hd__buf_2
X_14226_ _14226_/A VGND VGND VPWR VPWR _14665_/A sky130_fd_sc_hd__buf_2
XANTENNA__22125__A _22440_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14850__B _14850_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14157_ _14269_/A _24095_/Q VGND VGND VPWR VPWR _14158_/C sky130_fd_sc_hd__or2_4
X_13108_ _12962_/A _13108_/B _13107_/X VGND VGND VPWR VPWR _13124_/B sky130_fd_sc_hd__and3_4
X_18965_ _24370_/Q _18964_/A _18948_/C _18964_/Y VGND VGND VPWR VPWR _18965_/X sky130_fd_sc_hd__o22a_4
X_14088_ _14085_/X _14088_/B VGND VGND VPWR VPWR _14266_/A sky130_fd_sc_hd__or2_4
XANTENNA__12370__B _24012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21204__B2 _21202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13039_ _12498_/A _13109_/B VGND VGND VPWR VPWR _13041_/B sky130_fd_sc_hd__or2_4
X_17916_ _18409_/A _17913_/X _17916_/C _17916_/D VGND VGND VPWR VPWR _17917_/A sky130_fd_sc_hd__or4_4
XFILLER_65_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18896_ _18896_/A VGND VGND VPWR VPWR _18897_/A sky130_fd_sc_hd__buf_2
XFILLER_26_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17847_ _17847_/A VGND VGND VPWR VPWR _17848_/A sky130_fd_sc_hd__buf_2
XANTENNA__20963__B1 HRDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14578__A _14296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13482__A _12874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17778_ _17777_/X VGND VGND VPWR VPWR _17779_/D sky130_fd_sc_hd__inv_2
XFILLER_54_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22704__A1 _20486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21507__A2 _21506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22704__B2 _22698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19517_ HRDATA[30] VGND VGND VPWR VPWR _20672_/A sky130_fd_sc_hd__buf_2
XFILLER_81_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16729_ _16702_/A _16727_/X _16729_/C VGND VGND VPWR VPWR _16733_/B sky130_fd_sc_hd__and3_4
XANTENNA__12098__A _12097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18384__A1 _11633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19448_ HRDATA[16] _18576_/B _19447_/Y _24164_/Q _19438_/B VGND VGND VPWR VPWR _19448_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19379_ _19377_/X _19378_/Y _19377_/X _24247_/Q VGND VGND VPWR VPWR _19379_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12826__A _13343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21410_ _21299_/X _21405_/X _14400_/B _21409_/X VGND VGND VPWR VPWR _21410_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11730__A _16080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22390_ _22357_/A VGND VGND VPWR VPWR _22390_/X sky130_fd_sc_hd__buf_2
XFILLER_124_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21341_ _21341_/A VGND VGND VPWR VPWR _21341_/X sky130_fd_sc_hd__buf_2
XANTENNA__19609__A HRDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16828__A1_N _16905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24060_ _23592_/CLK _21071_/X VGND VGND VPWR VPWR _24060_/Q sky130_fd_sc_hd__dfxtp_4
X_21272_ _21271_/X _21269_/X _23944_/Q _21264_/X VGND VGND VPWR VPWR _21272_/X sky130_fd_sc_hd__o22a_4
XFILLER_162_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12184__A1 _12112_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23011_ _23008_/X _23009_/X _23010_/X VGND VGND VPWR VPWR _23011_/X sky130_fd_sc_hd__and3_4
XFILLER_144_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20223_ _20772_/A VGND VGND VPWR VPWR _20510_/A sky130_fd_sc_hd__inv_2
XFILLER_116_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24328__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21443__B2 _21438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17129__A _12097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12561__A _12561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20154_ _20154_/A VGND VGND VPWR VPWR _20154_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23140__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18886__C _17037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24266__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20085_ _18572_/X _20079_/X _20084_/Y _20066_/X VGND VGND VPWR VPWR _20085_/X sky130_fd_sc_hd__o22a_4
XFILLER_112_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21746__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23913_ _24073_/CLK _23913_/D VGND VGND VPWR VPWR _23913_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18072__B1 _18027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13392__A _13392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23844_ _23908_/CLK _21449_/X VGND VGND VPWR VPWR _15760_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23775_ _23679_/CLK _23775_/D VGND VGND VPWR VPWR _23775_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17799__A _18335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20987_ _11513_/Y _18835_/X VGND VGND VPWR VPWR _20987_/X sky130_fd_sc_hd__or2_4
XPHY_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22726_ _22705_/A VGND VGND VPWR VPWR _22726_/X sky130_fd_sc_hd__buf_2
XPHY_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22657_ _22435_/X _22651_/X _12816_/B _22655_/X VGND VGND VPWR VPWR _23146_/D sky130_fd_sc_hd__o22a_4
XFILLER_129_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12736__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12410_ _12410_/A VGND VGND VPWR VPWR _12957_/A sky130_fd_sc_hd__buf_2
XFILLER_22_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15112__A _15112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21608_ _21608_/A VGND VGND VPWR VPWR _21624_/A sky130_fd_sc_hd__inv_2
X_13390_ _13397_/A _24070_/Q VGND VGND VPWR VPWR _13390_/X sky130_fd_sc_hd__or2_4
Xclkbuf_4_11_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22588_ _22587_/X VGND VGND VPWR VPWR _22622_/A sky130_fd_sc_hd__buf_2
XANTENNA__21131__B1 _24021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19875__B2 _19811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12341_ _12370_/A _23756_/Q VGND VGND VPWR VPWR _12341_/X sky130_fd_sc_hd__or2_4
XFILLER_103_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21539_ _21824_/A VGND VGND VPWR VPWR _21539_/X sky130_fd_sc_hd__buf_2
X_24327_ _24292_/CLK _24327_/D HRESETn VGND VGND VPWR VPWR _19148_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21682__B2 _21681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15060_ _12329_/A _23765_/Q VGND VGND VPWR VPWR _15060_/X sky130_fd_sc_hd__or2_4
XFILLER_153_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12272_ _12727_/A _23628_/Q VGND VGND VPWR VPWR _12274_/B sky130_fd_sc_hd__or2_4
X_24258_ _24137_/CLK _24258_/D HRESETn VGND VGND VPWR VPWR _20713_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_49_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14011_ _13662_/A _14007_/X _14011_/C VGND VGND VPWR VPWR _14011_/X sky130_fd_sc_hd__or3_4
X_23209_ _23561_/CLK _23209_/D VGND VGND VPWR VPWR _12922_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_141_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13567__A _13566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12471__A _12492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24189_ _23671_/CLK _19866_/Y HRESETn VGND VGND VPWR VPWR _21133_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21985__A2 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21784__A _21770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15782__A _12676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18750_ _18158_/X VGND VGND VPWR VPWR _18750_/Y sky130_fd_sc_hd__inv_2
X_15962_ _16003_/A _15952_/X _15962_/C VGND VGND VPWR VPWR _15962_/X sky130_fd_sc_hd__or3_4
XFILLER_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21737__A2 _21734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17701_ _17775_/C _17698_/X _17700_/X VGND VGND VPWR VPWR _17701_/Y sky130_fd_sc_hd__o21ai_4
X_14913_ _12327_/A VGND VGND VPWR VPWR _14919_/A sky130_fd_sc_hd__buf_2
XFILLER_49_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18681_ _18176_/A _18675_/X _18677_/X _18679_/Y _18680_/X VGND VGND VPWR VPWR _18681_/X
+ sky130_fd_sc_hd__a32o_4
X_15893_ _13514_/A _15893_/B _15893_/C VGND VGND VPWR VPWR _15894_/C sky130_fd_sc_hd__and3_4
XANTENNA__23633__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20945__B1 _20561_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11815__A _13416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17632_ _17632_/A _17621_/B _17311_/Y _17632_/D VGND VGND VPWR VPWR _17632_/X sky130_fd_sc_hd__and4_4
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14844_ _14843_/X VGND VGND VPWR VPWR _14844_/X sky130_fd_sc_hd__buf_2
XFILLER_17_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17563_ _16383_/X _17561_/B VGND VGND VPWR VPWR _18039_/B sky130_fd_sc_hd__and2_4
XFILLER_91_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14775_ _14226_/A VGND VGND VPWR VPWR _15076_/A sky130_fd_sc_hd__buf_2
XFILLER_44_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11987_ _16713_/A _11985_/X _11987_/C VGND VGND VPWR VPWR _11987_/X sky130_fd_sc_hd__and3_4
X_19302_ _19235_/A _19235_/B _19301_/Y VGND VGND VPWR VPWR _19302_/X sky130_fd_sc_hd__o21a_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22162__A2 _22159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16514_ _16474_/A _16512_/X _16514_/C VGND VGND VPWR VPWR _16514_/X sky130_fd_sc_hd__and3_4
XFILLER_17_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23783__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13726_ _13753_/A _24030_/Q VGND VGND VPWR VPWR _13729_/B sky130_fd_sc_hd__or2_4
X_17494_ _17491_/Y _17021_/X _17029_/X _17493_/X VGND VGND VPWR VPWR _17530_/B sky130_fd_sc_hd__o22a_4
XFILLER_147_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19233_ _24284_/Q _19233_/B VGND VGND VPWR VPWR _19234_/B sky130_fd_sc_hd__and2_4
XFILLER_56_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16445_ _16401_/X _16445_/B VGND VGND VPWR VPWR _16445_/X sky130_fd_sc_hd__or2_4
X_13657_ _13657_/A _13653_/X _13657_/C VGND VGND VPWR VPWR _13661_/B sky130_fd_sc_hd__and3_4
XFILLER_108_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15022__A _15022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12608_ _12646_/A _12608_/B VGND VGND VPWR VPWR _12612_/B sky130_fd_sc_hd__or2_4
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19164_ _24339_/Q _19160_/B _19162_/Y VGND VGND VPWR VPWR _19164_/X sky130_fd_sc_hd__o21a_4
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16376_ _11702_/X _16374_/X _16375_/X VGND VGND VPWR VPWR _16377_/C sky130_fd_sc_hd__and3_4
XANTENNA__19554__A2_N _19551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13588_ _15029_/A VGND VGND VPWR VPWR _13589_/A sky130_fd_sc_hd__buf_2
XFILLER_157_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24139__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18115_ _18485_/A VGND VGND VPWR VPWR _18377_/A sky130_fd_sc_hd__buf_2
X_15327_ _11720_/A VGND VGND VPWR VPWR _15328_/A sky130_fd_sc_hd__buf_2
X_12539_ _12894_/A _12646_/B VGND VGND VPWR VPWR _12543_/B sky130_fd_sc_hd__or2_4
XANTENNA__21673__B2 _21667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22870__B1 _22799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19095_ _19074_/X _19093_/Y _19094_/Y _19079_/X VGND VGND VPWR VPWR _19095_/X sky130_fd_sc_hd__o22a_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24492__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18046_ _18046_/A VGND VGND VPWR VPWR _18046_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24375__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15258_ _14103_/A _15256_/X _15258_/C VGND VGND VPWR VPWR _15259_/C sky130_fd_sc_hd__and3_4
XFILLER_173_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14209_ _14254_/A _23167_/Q VGND VGND VPWR VPWR _14209_/X sky130_fd_sc_hd__or2_4
XANTENNA__21425__B2 _21424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12381__A _12978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24289__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15189_ _14235_/A _15125_/B VGND VGND VPWR VPWR _15191_/B sky130_fd_sc_hd__or2_4
XFILLER_153_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21976__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_31_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19997_ _19997_/A VGND VGND VPWR VPWR _24159_/D sky130_fd_sc_hd__inv_2
XFILLER_154_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18948_ _18948_/A _18948_/B _18948_/C _18948_/D VGND VGND VPWR VPWR _18949_/B sky130_fd_sc_hd__and4_4
XANTENNA__21728__A2 _21727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18879_ _14548_/X _18877_/X _24411_/Q _18878_/X VGND VGND VPWR VPWR _24411_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11725__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20910_ _24250_/Q VGND VGND VPWR VPWR _20910_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14101__A _11623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21890_ _21923_/A VGND VGND VPWR VPWR _21906_/A sky130_fd_sc_hd__inv_2
X_20841_ _20841_/A VGND VGND VPWR VPWR _20841_/X sky130_fd_sc_hd__buf_2
XFILLER_70_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19554__B1 _18782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13940__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23560_ _23337_/CLK _23560_/D VGND VGND VPWR VPWR _13006_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20772_ _20772_/A VGND VGND VPWR VPWR _20772_/X sky130_fd_sc_hd__buf_2
XANTENNA__21361__B1 _14452_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22511_ _22442_/X _22508_/X _13179_/B _22505_/X VGND VGND VPWR VPWR _22511_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21900__A2 _21895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23491_ _23587_/CLK _22069_/X VGND VGND VPWR VPWR _15833_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22442_ _20595_/A VGND VGND VPWR VPWR _22442_/X sky130_fd_sc_hd__buf_2
XANTENNA__21869__A _20860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20773__A _20895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21664__B2 _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22373_ _22358_/A VGND VGND VPWR VPWR _22373_/X sky130_fd_sc_hd__buf_2
XANTENNA__19339__A _19324_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21036__A2_N _21035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14771__A _14771_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23506__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_113_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR _23679_/CLK sky130_fd_sc_hd__clkbuf_1
X_24112_ _24080_/CLK _24112_/D VGND VGND VPWR VPWR _16436_/B sky130_fd_sc_hd__dfxtp_4
X_21324_ _21331_/A VGND VGND VPWR VPWR _21324_/X sky130_fd_sc_hd__buf_2
XFILLER_89_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14490__B _14490_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24043_ _24074_/CLK _24043_/D VGND VGND VPWR VPWR _12608_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21255_ _21254_/X _21245_/X _16270_/B _21252_/X VGND VGND VPWR VPWR _21255_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21416__B2 _21381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20206_ _24469_/Q VGND VGND VPWR VPWR _20206_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21186_ _21219_/A VGND VGND VPWR VPWR _21202_/A sky130_fd_sc_hd__inv_2
XANTENNA__18832__A2 _18796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20137_ _11563_/X VGND VGND VPWR VPWR _20137_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21719__A2 _21713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20068_ _20064_/X _18367_/A _20046_/X _20067_/X VGND VGND VPWR VPWR _20069_/A sky130_fd_sc_hd__o22a_4
XFILLER_38_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19793__B1 _22737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11635__A _11635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22392__A2 _22390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11910_ _11910_/A VGND VGND VPWR VPWR _12233_/A sky130_fd_sc_hd__buf_2
X_12890_ _12890_/A _12886_/X _12890_/C VGND VGND VPWR VPWR _12890_/X sky130_fd_sc_hd__or3_4
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14011__A _13662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23827_ _23764_/CLK _23827_/D VGND VGND VPWR VPWR _23827_/Q sky130_fd_sc_hd__dfxtp_4
X_11841_ _12166_/A _11841_/B VGND VGND VPWR VPWR _11844_/B sky130_fd_sc_hd__or2_4
XPHY_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _16049_/A VGND VGND VPWR VPWR _11772_/X sky130_fd_sc_hd__buf_2
X_14560_ _14278_/A _14560_/B VGND VGND VPWR VPWR _14562_/B sky130_fd_sc_hd__or2_4
XPHY_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23758_ _23501_/CLK _21621_/X VGND VGND VPWR VPWR _23758_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _12950_/A VGND VGND VPWR VPWR _13514_/A sky130_fd_sc_hd__buf_2
XPHY_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22709_ _21268_/A _22708_/X _12963_/B _22705_/X VGND VGND VPWR VPWR _23113_/D sky130_fd_sc_hd__o22a_4
X_14491_ _12372_/A _14491_/B VGND VGND VPWR VPWR _14493_/B sky130_fd_sc_hd__or2_4
XFILLER_14_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12466__A _12466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23689_ _23337_/CLK _21728_/X VGND VGND VPWR VPWR _23689_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16230_ _16181_/X _23501_/Q VGND VGND VPWR VPWR _16230_/X sky130_fd_sc_hd__or2_4
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13442_ _12872_/A VGND VGND VPWR VPWR _13443_/A sky130_fd_sc_hd__buf_2
XANTENNA__15582__A1 _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16161_ _11973_/X _16138_/X _16145_/X _16152_/X _16160_/X VGND VGND VPWR VPWR _16161_/X
+ sky130_fd_sc_hd__a32o_4
X_13373_ _13392_/A _13366_/X _13373_/C VGND VGND VPWR VPWR _13373_/X sky130_fd_sc_hd__or3_4
XFILLER_6_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23186__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18153__A _18545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15112_ _15112_/A _15110_/X _15112_/C VGND VGND VPWR VPWR _15113_/C sky130_fd_sc_hd__and3_4
X_12324_ _13230_/A VGND VGND VPWR VPWR _12827_/A sky130_fd_sc_hd__buf_2
X_16092_ _16110_/A _16092_/B _16091_/X VGND VGND VPWR VPWR _16092_/X sky130_fd_sc_hd__and3_4
X_12255_ _12279_/A _12253_/X _12255_/C VGND VGND VPWR VPWR _12261_/B sky130_fd_sc_hd__and3_4
X_19920_ _22738_/A VGND VGND VPWR VPWR _19920_/X sky130_fd_sc_hd__buf_2
X_15043_ _13662_/A _15043_/B _15043_/C VGND VGND VPWR VPWR _15044_/B sky130_fd_sc_hd__or3_4
XANTENNA__21958__A2 _21953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19851_ _19848_/A _19843_/X VGND VGND VPWR VPWR _19851_/X sky130_fd_sc_hd__or2_4
XFILLER_69_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12186_ _12186_/A VGND VGND VPWR VPWR _13045_/A sky130_fd_sc_hd__buf_2
XFILLER_134_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22080__B2 _22078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_18_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_96_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18802_ _12678_/X _18796_/X _11554_/A _18797_/X VGND VGND VPWR VPWR _18802_/X sky130_fd_sc_hd__o22a_4
X_19782_ _19732_/X _19775_/X _19781_/X _16683_/A _19719_/X VGND VGND VPWR VPWR _19782_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16401__A _12559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16994_ _16950_/Y _16994_/B VGND VGND VPWR VPWR _16995_/B sky130_fd_sc_hd__or2_4
XFILLER_7_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18733_ _17797_/A _18732_/X _17341_/B VGND VGND VPWR VPWR _18733_/X sky130_fd_sc_hd__o21a_4
XFILLER_62_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15945_ _15982_/A _23758_/Q VGND VGND VPWR VPWR _15946_/C sky130_fd_sc_hd__or2_4
XFILLER_114_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15017__A _15017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18664_ _17756_/X _17747_/X _17743_/X VGND VGND VPWR VPWR _18664_/X sky130_fd_sc_hd__o21a_4
X_15876_ _13546_/A _15807_/B VGND VGND VPWR VPWR _15876_/X sky130_fd_sc_hd__or2_4
XFILLER_64_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21591__B1 _14633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17615_ _17615_/A _17614_/X VGND VGND VPWR VPWR _17616_/B sky130_fd_sc_hd__and2_4
X_14827_ _14834_/A _14827_/B VGND VGND VPWR VPWR _14827_/X sky130_fd_sc_hd__or2_4
X_18595_ _17758_/X _17739_/X _17734_/X VGND VGND VPWR VPWR _18595_/X sky130_fd_sc_hd__o21a_4
XFILLER_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13760__A _12925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17546_ _17545_/X VGND VGND VPWR VPWR _17546_/Y sky130_fd_sc_hd__inv_2
X_14758_ _13630_/A _14758_/B VGND VGND VPWR VPWR _14758_/X sky130_fd_sc_hd__or2_4
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13709_ _12634_/A VGND VGND VPWR VPWR _13774_/A sky130_fd_sc_hd__buf_2
X_17477_ _17145_/Y _17475_/B VGND VGND VPWR VPWR _17478_/B sky130_fd_sc_hd__and2_4
XANTENNA__12376__A _15851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14689_ _14680_/A _14689_/B _14689_/C VGND VGND VPWR VPWR _14690_/C sky130_fd_sc_hd__and3_4
XANTENNA__23529__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19216_ _19134_/A _19133_/X _19215_/Y VGND VGND VPWR VPWR _19216_/X sky130_fd_sc_hd__o21a_4
X_16428_ _16402_/X _16428_/B VGND VGND VPWR VPWR _16428_/X sky130_fd_sc_hd__or2_4
XANTENNA__20593__A _20535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15687__A _12696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19147_ _19147_/A _19146_/X VGND VGND VPWR VPWR _19148_/B sky130_fd_sc_hd__and2_4
XANTENNA__21646__A1 _21584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16359_ _16465_/A _16359_/B _16358_/X VGND VGND VPWR VPWR _16359_/X sky130_fd_sc_hd__and3_4
XANTENNA__21646__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14591__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20854__C1 _20853_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19078_ _19078_/A VGND VGND VPWR VPWR _19078_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18029_ _16949_/A _18028_/Y _16996_/B VGND VGND VPWR VPWR _23054_/B sky130_fd_sc_hd__o21a_4
XFILLER_160_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21949__A2 _21946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21040_ _20361_/X _21038_/X _24082_/Q _21035_/X VGND VGND VPWR VPWR _21040_/X sky130_fd_sc_hd__o22a_4
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13935__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22991_ _18426_/X _22973_/B VGND VGND VPWR VPWR _22992_/C sky130_fd_sc_hd__or2_4
XFILLER_95_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22374__A2 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21942_ _21957_/A VGND VGND VPWR VPWR _21950_/A sky130_fd_sc_hd__buf_2
XFILLER_41_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_38_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR _23760_/CLK sky130_fd_sc_hd__clkbuf_1
X_21873_ _21872_/X _21863_/X _14455_/B _21870_/X VGND VGND VPWR VPWR _23611_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24304__CLK _24306_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22126__A2 _22123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13670__A _12251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _23675_/CLK _21871_/X VGND VGND VPWR VPWR _14380_/B sky130_fd_sc_hd__dfxtp_4
X_20824_ _20778_/A _20824_/B VGND VGND VPWR VPWR _20824_/X sky130_fd_sc_hd__or2_4
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14485__B _14485_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22983__A _22982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20755_ _20315_/X VGND VGND VPWR VPWR _20755_/X sky130_fd_sc_hd__buf_2
X_23543_ _23991_/CLK _23543_/D VGND VGND VPWR VPWR _15143_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12286__A _11930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23474_ _23922_/CLK _22102_/X VGND VGND VPWR VPWR _16640_/B sky130_fd_sc_hd__dfxtp_4
X_20686_ _18448_/X _20675_/X _20538_/X _20685_/Y VGND VGND VPWR VPWR _20686_/X sky130_fd_sc_hd__a211o_4
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22425_ _22110_/A VGND VGND VPWR VPWR _22425_/X sky130_fd_sc_hd__buf_2
XANTENNA__21637__B2 _21631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18502__A1 _18111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22356_ _22355_/X VGND VGND VPWR VPWR _22357_/A sky130_fd_sc_hd__buf_2
XFILLER_109_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21307_ _20938_/A VGND VGND VPWR VPWR _21307_/X sky130_fd_sc_hd__buf_2
X_22287_ _22294_/A VGND VGND VPWR VPWR _22287_/X sky130_fd_sc_hd__buf_2
XFILLER_3_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17069__A1 _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24026_ _24057_/CLK _24026_/D VGND VGND VPWR VPWR _14563_/B sky130_fd_sc_hd__dfxtp_4
X_12040_ _11941_/A VGND VGND VPWR VPWR _12041_/A sky130_fd_sc_hd__buf_2
XANTENNA__22062__A1 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21238_ _21238_/A VGND VGND VPWR VPWR _21264_/A sky130_fd_sc_hd__inv_2
XANTENNA__22062__B2 _22057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21169_ _21136_/A VGND VGND VPWR VPWR _21169_/X sky130_fd_sc_hd__buf_2
XFILLER_172_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17036__B _17251_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13991_ _13607_/A _23840_/Q VGND VGND VPWR VPWR _13991_/X sky130_fd_sc_hd__or2_4
XANTENNA__18569__B2 _18568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22365__A2 _22362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15730_ _12783_/X _15668_/B VGND VGND VPWR VPWR _15730_/X sky130_fd_sc_hd__or2_4
X_12942_ _12942_/A _23337_/Q VGND VGND VPWR VPWR _12944_/B sky130_fd_sc_hd__or2_4
XFILLER_58_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23054__A _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15661_ _12690_/A _23748_/Q VGND VGND VPWR VPWR _15662_/C sky130_fd_sc_hd__or2_4
X_12873_ _12873_/A _12871_/X _12872_/X VGND VGND VPWR VPWR _12874_/C sky130_fd_sc_hd__and3_4
XFILLER_2_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18148__A _18148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17400_ _17397_/Y _17019_/X _17027_/X _17399_/X VGND VGND VPWR VPWR _17402_/A sky130_fd_sc_hd__o22a_4
X_14612_ _14450_/A _14589_/X _14596_/X _14603_/X _14611_/X VGND VGND VPWR VPWR _14612_/X
+ sky130_fd_sc_hd__a32o_4
X_18380_ _18379_/X VGND VGND VPWR VPWR _18380_/Y sky130_fd_sc_hd__inv_2
X_11824_ _11717_/X _11824_/B VGND VGND VPWR VPWR _11824_/X sky130_fd_sc_hd__or2_4
X_15592_ _11710_/A _23201_/Q VGND VGND VPWR VPWR _15594_/B sky130_fd_sc_hd__or2_4
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17332_/B VGND VGND VPWR VPWR _17333_/B sky130_fd_sc_hd__inv_2
XFILLER_159_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14543_/A _14541_/X _14543_/C VGND VGND VPWR VPWR _14543_/X sky130_fd_sc_hd__and3_4
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _13063_/A VGND VGND VPWR VPWR _11755_/X sky130_fd_sc_hd__buf_2
XANTENNA__21876__B2 _21870_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _17398_/A _17251_/B VGND VGND VPWR VPWR _17262_/X sky130_fd_sc_hd__and2_4
XFILLER_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14474_ _15400_/A _14474_/B VGND VGND VPWR VPWR _14475_/C sky130_fd_sc_hd__or2_4
X_11686_ _16187_/A VGND VGND VPWR VPWR _11686_/X sky130_fd_sc_hd__buf_2
XFILLER_128_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19001_ _24396_/Q VGND VGND VPWR VPWR _19001_/Y sky130_fd_sc_hd__inv_2
X_16213_ _16185_/A _16211_/X _16213_/C VGND VGND VPWR VPWR _16214_/C sky130_fd_sc_hd__and3_4
XFILLER_174_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13425_ _13468_/A _13421_/X _13424_/X VGND VGND VPWR VPWR _13425_/X sky130_fd_sc_hd__or3_4
XFILLER_127_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21302__A _20892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21628__B2 _21624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17193_ _17198_/A VGND VGND VPWR VPWR _17193_/X sky130_fd_sc_hd__buf_2
XANTENNA__12924__A _12950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15300__A _14295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16144_ _16144_/A _16142_/X _16143_/X VGND VGND VPWR VPWR _16145_/C sky130_fd_sc_hd__and3_4
X_13356_ _13384_/A _13283_/B VGND VGND VPWR VPWR _13358_/B sky130_fd_sc_hd__or2_4
XANTENNA__12643__B _12533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12307_ _12741_/A _12303_/X _12307_/C VGND VGND VPWR VPWR _12307_/X sky130_fd_sc_hd__and3_4
X_16075_ _11693_/X _16075_/B _16074_/X VGND VGND VPWR VPWR _16083_/B sky130_fd_sc_hd__or3_4
X_13287_ _13313_/A _23302_/Q VGND VGND VPWR VPWR _13288_/C sky130_fd_sc_hd__or2_4
XANTENNA__18611__A _18610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19903_ _19903_/A _19903_/B VGND VGND VPWR VPWR _19903_/X sky130_fd_sc_hd__or2_4
X_15026_ _13983_/A _23381_/Q VGND VGND VPWR VPWR _15028_/B sky130_fd_sc_hd__or2_4
X_12238_ _12213_/A VGND VGND VPWR VPWR _12239_/A sky130_fd_sc_hd__buf_2
XFILLER_170_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13755__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12169_ _12169_/A _12169_/B _12169_/C VGND VGND VPWR VPWR _12177_/B sky130_fd_sc_hd__or3_4
X_19834_ _19834_/A _19665_/B _19833_/X VGND VGND VPWR VPWR _19834_/X sky130_fd_sc_hd__or3_4
XANTENNA__21800__B2 _21795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23201__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19765_ _19834_/A _19765_/B VGND VGND VPWR VPWR _19765_/X sky130_fd_sc_hd__or2_4
X_16977_ _17727_/A _16976_/X VGND VGND VPWR VPWR _16977_/X sky130_fd_sc_hd__or2_4
XANTENNA__24327__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19442__A _18576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18716_ _18716_/A VGND VGND VPWR VPWR _18716_/Y sky130_fd_sc_hd__inv_2
X_15928_ _15917_/X _15926_/Y _15788_/A _15927_/Y VGND VGND VPWR VPWR _15929_/A sky130_fd_sc_hd__a211o_4
X_19696_ _19447_/Y VGND VGND VPWR VPWR _19696_/X sky130_fd_sc_hd__buf_2
X_18647_ _18646_/X VGND VGND VPWR VPWR _24475_/D sky130_fd_sc_hd__inv_2
X_15859_ _12402_/X _15857_/X _15858_/X VGND VGND VPWR VPWR _15859_/X sky130_fd_sc_hd__and3_4
XFILLER_92_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14586__A _12530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24477__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18578_ _17732_/A _18577_/X VGND VGND VPWR VPWR _18578_/X sky130_fd_sc_hd__or2_4
XANTENNA__21316__B1 _23925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17529_ _17515_/B VGND VGND VPWR VPWR _18280_/B sky130_fd_sc_hd__inv_2
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20540_ _20315_/A VGND VGND VPWR VPWR _20540_/X sky130_fd_sc_hd__buf_2
XANTENNA__22308__A _22275_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21212__A _21198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21619__B2 _21617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20471_ _20282_/A VGND VGND VPWR VPWR _20471_/X sky130_fd_sc_hd__buf_2
XANTENNA__12834__A _12834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16306__A _15934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22210_ _22149_/X _22208_/X _13761_/B _22205_/X VGND VGND VPWR VPWR _23422_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17299__A1 _14767_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21095__A2 _21090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23190_ _23862_/CLK _23190_/D VGND VGND VPWR VPWR _23190_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_173_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22292__B2 _22291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11583__A2 IRQ[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22141_ _20744_/A VGND VGND VPWR VPWR _22141_/X sky130_fd_sc_hd__buf_2
XFILLER_134_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22044__B2 _22043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22072_ _21857_/X _22067_/X _15566_/B _22071_/X VGND VGND VPWR VPWR _22072_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22043__A _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18799__A1 _17139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21023_ _22169_/A VGND VGND VPWR VPWR _21024_/A sky130_fd_sc_hd__buf_2
XANTENNA__22595__A2 _22594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13665__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16041__A _16048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22978__A _22912_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15880__A _13530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22974_ _22947_/X _22974_/B _22974_/C VGND VGND VPWR VPWR _22974_/X sky130_fd_sc_hd__and3_4
X_21925_ _21865_/X _21923_/X _13733_/B _21920_/X VGND VGND VPWR VPWR _23582_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11913__A _11913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21856_ _21855_/X _21851_/X _15489_/B _21846_/X VGND VGND VPWR VPWR _23618_/D sky130_fd_sc_hd__o22a_4
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _24414_/Q _20645_/X _24446_/Q _20704_/X VGND VGND VPWR VPWR _20807_/X sky130_fd_sc_hd__o22a_4
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21787_ _21570_/X _21784_/X _15512_/B _21781_/X VGND VGND VPWR VPWR _23650_/D sky130_fd_sc_hd__o22a_4
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23526_ _23723_/CLK _22015_/X VGND VGND VPWR VPWR _13274_/B sky130_fd_sc_hd__dfxtp_4
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _24366_/Q _11540_/B VGND VGND VPWR VPWR _11541_/B sky130_fd_sc_hd__or2_4
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20738_ _18494_/X _20675_/X _20538_/X _20737_/Y VGND VGND VPWR VPWR _20738_/X sky130_fd_sc_hd__a211o_4
XFILLER_11_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14943__B _23990_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21122__A _21101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20669_ HRDATA[14] _20697_/A VGND VGND VPWR VPWR _20669_/X sky130_fd_sc_hd__or2_4
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23457_ _23617_/CLK _23457_/D VGND VGND VPWR VPWR _15607_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ _13258_/A _13210_/B _13210_/C VGND VGND VPWR VPWR _13210_/X sky130_fd_sc_hd__or3_4
X_22408_ _22433_/A VGND VGND VPWR VPWR _22421_/A sky130_fd_sc_hd__buf_2
X_14190_ _14200_/A _23743_/Q VGND VGND VPWR VPWR _14190_/X sky130_fd_sc_hd__or2_4
XFILLER_87_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22283__B2 _22277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23388_ _23772_/CLK _22263_/X VGND VGND VPWR VPWR _14391_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_104_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12463__B _12599_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11574__A2 IRQ[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13141_ _12726_/A _13136_/X _13141_/C VGND VGND VPWR VPWR _13141_/X sky130_fd_sc_hd__or3_4
X_22339_ _23331_/Q VGND VGND VPWR VPWR _23331_/D sky130_fd_sc_hd__buf_2
XFILLER_125_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19527__A _19624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13072_ _13100_/A _13072_/B _13072_/C VGND VGND VPWR VPWR _13073_/C sky130_fd_sc_hd__or3_4
XFILLER_152_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23049__A _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22035__B2 _22000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16900_ _17060_/A VGND VGND VPWR VPWR _16915_/A sky130_fd_sc_hd__buf_2
X_12023_ _11851_/X VGND VGND VPWR VPWR _12024_/A sky130_fd_sc_hd__inv_2
X_24009_ _23337_/CLK _21156_/X VGND VGND VPWR VPWR _24009_/Q sky130_fd_sc_hd__dfxtp_4
X_17880_ _17880_/A VGND VGND VPWR VPWR _17880_/X sky130_fd_sc_hd__buf_2
XANTENNA__20597__A1 _20533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20597__B2 _20510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16831_ _16831_/A _16831_/B _13272_/X _16830_/X VGND VGND VPWR VPWR _16831_/X sky130_fd_sc_hd__or4_4
XANTENNA__19739__B1 _17820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19550_ _19687_/D _19550_/B _19550_/C _19550_/D VGND VGND VPWR VPWR _19550_/X sky130_fd_sc_hd__and4_4
X_16762_ _16639_/A _23793_/Q VGND VGND VPWR VPWR _16763_/C sky130_fd_sc_hd__or2_4
X_13974_ _13974_/A _14035_/B VGND VGND VPWR VPWR _13976_/B sky130_fd_sc_hd__or2_4
XFILLER_24_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18501_ _18500_/A _16979_/X _18479_/Y VGND VGND VPWR VPWR _22966_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__17214__A1 _17145_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15713_ _12851_/A _15713_/B _15712_/X VGND VGND VPWR VPWR _15714_/C sky130_fd_sc_hd__and3_4
X_12925_ _12925_/A VGND VGND VPWR VPWR _12951_/A sky130_fd_sc_hd__buf_2
X_19481_ _19455_/Y VGND VGND VPWR VPWR _19481_/X sky130_fd_sc_hd__buf_2
XFILLER_46_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16693_ _16586_/A _16756_/B VGND VGND VPWR VPWR _16695_/B sky130_fd_sc_hd__or2_4
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17765__A2 _17360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18432_ _18368_/A _18368_/B VGND VGND VPWR VPWR _18432_/Y sky130_fd_sc_hd__nand2_4
XFILLER_146_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_21_0_HCLK clkbuf_6_10_0_HCLK/X VGND VGND VPWR VPWR _24134_/CLK sky130_fd_sc_hd__clkbuf_1
X_15644_ _13884_/A _15569_/B VGND VGND VPWR VPWR _15646_/B sky130_fd_sc_hd__or2_4
X_12856_ _12886_/A _12856_/B _12855_/X VGND VGND VPWR VPWR _12857_/C sky130_fd_sc_hd__and3_4
XFILLER_18_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_84_0_HCLK clkbuf_6_42_0_HCLK/X VGND VGND VPWR VPWR _23544_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21849__A1 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11807_ _12169_/A _11807_/B _11807_/C VGND VGND VPWR VPWR _11807_/X sky130_fd_sc_hd__or3_4
X_18363_ _18553_/A _17906_/C VGND VGND VPWR VPWR _18533_/B sky130_fd_sc_hd__or2_4
XANTENNA__21849__B2 _21846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15575_ _12427_/A _15573_/X _15574_/X VGND VGND VPWR VPWR _15575_/X sky130_fd_sc_hd__and3_4
X_12787_ _13563_/A _12776_/X _12786_/X VGND VGND VPWR VPWR _12787_/X sky130_fd_sc_hd__or3_4
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22510__A2 _22508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19911__B1 _19910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17314_ _14845_/Y _17300_/B VGND VGND VPWR VPWR _18673_/B sky130_fd_sc_hd__or2_4
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14519_/A _14462_/B VGND VGND VPWR VPWR _14526_/X sky130_fd_sc_hd__or2_4
X_11738_ _13232_/A VGND VGND VPWR VPWR _11739_/A sky130_fd_sc_hd__buf_2
X_18294_ _17509_/Y _18293_/X _17531_/X VGND VGND VPWR VPWR _18294_/X sky130_fd_sc_hd__o21a_4
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ _17245_/A VGND VGND VPWR VPWR _17245_/X sky130_fd_sc_hd__buf_2
X_14457_ _12428_/A _14455_/X _14457_/C VGND VGND VPWR VPWR _14458_/C sky130_fd_sc_hd__and3_4
XANTENNA__12654__A _12623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11669_ _12979_/A VGND VGND VPWR VPWR _13566_/A sky130_fd_sc_hd__buf_2
XANTENNA__16126__A _16099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _13408_/A _23494_/Q VGND VGND VPWR VPWR _13410_/B sky130_fd_sc_hd__or2_4
XANTENNA__21077__A2 _21073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17176_ _15786_/Y _17107_/X _13583_/X _17074_/X VGND VGND VPWR VPWR _17176_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21967__A _21960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14388_ _14378_/A _14388_/B VGND VGND VPWR VPWR _14388_/X sky130_fd_sc_hd__or2_4
X_16127_ _16157_/A _16196_/B VGND VGND VPWR VPWR _16128_/C sky130_fd_sc_hd__or2_4
X_13339_ _13339_/A _13339_/B VGND VGND VPWR VPWR _13339_/X sky130_fd_sc_hd__and2_4
XFILLER_127_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22026__A1 _21865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16058_ _16046_/A _24078_/Q VGND VGND VPWR VPWR _16059_/C sky130_fd_sc_hd__or2_4
XANTENNA__22026__B2 _22021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15009_ _13955_/A _15009_/B _15009_/C VGND VGND VPWR VPWR _15009_/X sky130_fd_sc_hd__and3_4
XFILLER_142_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23717__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19817_ _19831_/A _19816_/X _19894_/C VGND VGND VPWR VPWR _19817_/X sky130_fd_sc_hd__o21a_4
XFILLER_96_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19748_ _19683_/A _19677_/A _19748_/C VGND VGND VPWR VPWR _19748_/X sky130_fd_sc_hd__or3_4
XFILLER_42_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17205__A1 _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19679_ _19831_/A _19894_/C _19744_/A _19678_/X VGND VGND VPWR VPWR _19679_/X sky130_fd_sc_hd__a211o_4
X_21710_ _21717_/A VGND VGND VPWR VPWR _21710_/X sky130_fd_sc_hd__buf_2
X_22690_ _22705_/A VGND VGND VPWR VPWR _22698_/A sky130_fd_sc_hd__buf_2
XANTENNA__12548__B _12548_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21641_ _21608_/A VGND VGND VPWR VPWR _21641_/X sky130_fd_sc_hd__buf_2
XFILLER_40_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17420__A _17161_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21572_ _20745_/A VGND VGND VPWR VPWR _21572_/X sky130_fd_sc_hd__buf_2
X_24360_ _24360_/CLK _24360_/D HRESETn VGND VGND VPWR VPWR _24360_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_166_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23311_ _23119_/CLK _22368_/X VGND VGND VPWR VPWR _16260_/B sky130_fd_sc_hd__dfxtp_4
X_20523_ _20515_/X _20521_/X _19151_/A _20522_/X VGND VGND VPWR VPWR _20523_/X sky130_fd_sc_hd__o22a_4
X_24291_ _24292_/CLK _24291_/D HRESETn VGND VGND VPWR VPWR _19240_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12564__A _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16036__A _11759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23242_ _23531_/CLK _23242_/D VGND VGND VPWR VPWR _12836_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21068__A2 _21066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20454_ _20315_/X _20453_/X _18994_/A _20325_/X VGND VGND VPWR VPWR _20454_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18469__B1 _18467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23173_ _23397_/CLK _22614_/X VGND VGND VPWR VPWR _13449_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15875__A _13543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19347__A _19340_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20385_ _20273_/X _20384_/X _19253_/A _20349_/X VGND VGND VPWR VPWR _20385_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17141__B1 _17140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22124_ _22122_/X _22123_/X _23465_/Q _22118_/X VGND VGND VPWR VPWR _22124_/X sky130_fd_sc_hd__o22a_4
X_22055_ _21829_/X _22053_/X _23501_/Q _22050_/X VGND VGND VPWR VPWR _22055_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11908__A _16595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21006_ _20940_/A HRDATA[16] VGND VGND VPWR VPWR _21006_/X sky130_fd_sc_hd__or2_4
XFILLER_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18641__B1 _17792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22501__A _22508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22957_ _22946_/X _18553_/A _22909_/X _22956_/X VGND VGND VPWR VPWR _22957_/X sky130_fd_sc_hd__a211o_4
XFILLER_16_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12710_ _12269_/A _12790_/B VGND VGND VPWR VPWR _12710_/X sky130_fd_sc_hd__or2_4
XANTENNA__11643__A _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15115__A _15649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21908_ _21836_/X _21902_/X _12790_/B _21906_/X VGND VGND VPWR VPWR _21908_/X sky130_fd_sc_hd__o22a_4
X_13690_ _11969_/A _13661_/X _13674_/X _13681_/X _13689_/X VGND VGND VPWR VPWR _13690_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_44_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22888_ _22897_/A _22887_/X VGND VGND VPWR VPWR HWDATA[26] sky130_fd_sc_hd__nor2_4
XANTENNA__20956__A _20977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12641_ _12641_/A _12614_/X _12641_/C VGND VGND VPWR VPWR _12677_/B sky130_fd_sc_hd__or3_4
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21839_ _21839_/A VGND VGND VPWR VPWR _21839_/X sky130_fd_sc_hd__buf_2
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24022__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ _11735_/A _15360_/B _15359_/X VGND VGND VPWR VPWR _15360_/X sky130_fd_sc_hd__and3_4
X_12572_ _12912_/A _12571_/X VGND VGND VPWR VPWR _12572_/X sky130_fd_sc_hd__and2_4
XFILLER_19_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ _14311_/A _14387_/B VGND VGND VPWR VPWR _14313_/B sky130_fd_sc_hd__or2_4
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _11523_/A _11523_/B VGND VGND VPWR VPWR _11524_/B sky130_fd_sc_hd__or2_4
X_23509_ _23509_/CLK _22037_/X VGND VGND VPWR VPWR _23509_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15291_ _14269_/A _23832_/Q VGND VGND VPWR VPWR _15291_/X sky130_fd_sc_hd__or2_4
X_24489_ _24294_/CLK _24489_/D HRESETn VGND VGND VPWR VPWR _24489_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17030_ _17029_/X VGND VGND VPWR VPWR _17031_/A sky130_fd_sc_hd__buf_2
XFILLER_109_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14242_ _14615_/A _14242_/B _14241_/X VGND VGND VPWR VPWR _14242_/X sky130_fd_sc_hd__or3_4
XANTENNA__22256__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24172__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15785__A _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14173_ _14012_/A _14172_/X VGND VGND VPWR VPWR _14173_/X sky130_fd_sc_hd__and2_4
XANTENNA__19672__A2 HRDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13124_ _12676_/A _13124_/B _13124_/C VGND VGND VPWR VPWR _13124_/X sky130_fd_sc_hd__or3_4
XFILLER_98_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22008__B2 _22007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18981_ _11541_/B VGND VGND VPWR VPWR _18981_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22559__A2 _22558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13055_ _13055_/A VGND VGND VPWR VPWR _13095_/A sky130_fd_sc_hd__buf_2
X_17932_ _17236_/X _17189_/X VGND VGND VPWR VPWR _17932_/Y sky130_fd_sc_hd__nor2_4
XFILLER_65_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12006_ _12001_/X _12006_/B _12006_/C VGND VGND VPWR VPWR _12010_/B sky130_fd_sc_hd__and3_4
XFILLER_39_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21231__A2 _21226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17863_ _17229_/X _17859_/X _17823_/X _17862_/X VGND VGND VPWR VPWR _17864_/A sky130_fd_sc_hd__o22a_4
XANTENNA__19975__A3 _19969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19602_ _19612_/A VGND VGND VPWR VPWR _19895_/A sky130_fd_sc_hd__buf_2
XFILLER_66_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16814_ _16611_/A _23665_/Q VGND VGND VPWR VPWR _16814_/X sky130_fd_sc_hd__or2_4
X_17794_ _17912_/A VGND VGND VPWR VPWR _18222_/A sky130_fd_sc_hd__buf_2
X_19533_ _19899_/B _19533_/B VGND VGND VPWR VPWR _19550_/C sky130_fd_sc_hd__or2_4
XFILLER_47_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16745_ _11990_/A _23889_/Q VGND VGND VPWR VPWR _16746_/C sky130_fd_sc_hd__or2_4
X_13957_ _13957_/A _23744_/Q VGND VGND VPWR VPWR _13958_/C sky130_fd_sc_hd__or2_4
XANTENNA__17199__B1 _15382_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12649__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22192__B1 _12657_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22731__A2 _22729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12908_ _12510_/A _23721_/Q VGND VGND VPWR VPWR _12908_/X sky130_fd_sc_hd__or2_4
X_19464_ _19507_/A _19839_/A VGND VGND VPWR VPWR _19465_/A sky130_fd_sc_hd__or2_4
XANTENNA__15025__A _13965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16676_ _16676_/A _23506_/Q VGND VGND VPWR VPWR _16676_/X sky130_fd_sc_hd__or2_4
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13888_ _13888_/A VGND VGND VPWR VPWR _13916_/A sky130_fd_sc_hd__buf_2
X_18415_ _18415_/A _18415_/B _18415_/C VGND VGND VPWR VPWR _18416_/B sky130_fd_sc_hd__or3_4
X_15627_ _15611_/A _15560_/B VGND VGND VPWR VPWR _15627_/X sky130_fd_sc_hd__or2_4
X_12839_ _13563_/A _12839_/B _12839_/C VGND VGND VPWR VPWR _12840_/C sky130_fd_sc_hd__or3_4
X_19395_ _19392_/X _18073_/Y _19392_/X _24238_/Q VGND VGND VPWR VPWR _24238_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18346_ _18293_/X VGND VGND VPWR VPWR _18346_/Y sky130_fd_sc_hd__inv_2
X_15558_ _15442_/A _15558_/B _15557_/X VGND VGND VPWR VPWR _15558_/X sky130_fd_sc_hd__or3_4
XANTENNA__21298__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22495__B2 _22491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14509_ _14509_/A _14506_/X _14509_/C VGND VGND VPWR VPWR _14513_/B sky130_fd_sc_hd__and3_4
X_18277_ _17686_/A _16988_/B _16989_/B VGND VGND VPWR VPWR _23014_/B sky130_fd_sc_hd__a21bo_4
XANTENNA__12384__A _11739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15489_ _13744_/A _15489_/B VGND VGND VPWR VPWR _15491_/B sky130_fd_sc_hd__or2_4
X_17228_ _17137_/X VGND VGND VPWR VPWR _17878_/A sky130_fd_sc_hd__buf_2
XANTENNA__13199__B _13199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22247__B2 _22241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17159_ _12093_/X VGND VGND VPWR VPWR _17836_/A sky130_fd_sc_hd__buf_2
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17674__A1 _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20170_ _24438_/Q IRQ[1] _11552_/Y _24440_/Q IRQ[3] VGND VGND VPWR VPWR _20170_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_66_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13160__A1 _13339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17415__A _22039_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13943__A _13894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23860_ _23668_/CLK _23860_/D VGND VGND VPWR VPWR _23860_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20981__A1 _20894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20981__B2 _20396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22811_ _14483_/Y _22803_/X VGND VGND VPWR VPWR HWDATA[6] sky130_fd_sc_hd__nor2_4
XFILLER_38_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23791_ _23662_/CLK _23791_/D VGND VGND VPWR VPWR _16257_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12559__A _12559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18926__A1 _15651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22742_ _22742_/A VGND VGND VPWR VPWR _23086_/A sky130_fd_sc_hd__buf_2
XFILLER_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20776__A _20776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22673_ _22461_/X _22672_/X _23135_/Q _22669_/X VGND VGND VPWR VPWR _22673_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14774__A _15103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24412_ _24445_/CLK _18876_/X HRESETn VGND VGND VPWR VPWR _24412_/Q sky130_fd_sc_hd__dfrtp_4
X_21624_ _21624_/A VGND VGND VPWR VPWR _21624_/X sky130_fd_sc_hd__buf_2
XANTENNA__21289__A2 _21281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22991__A _18426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14493__B _14493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24343_ _24342_/CLK _24343_/D HRESETn VGND VGND VPWR VPWR _11514_/A sky130_fd_sc_hd__dfstp_4
X_21555_ _21553_/X _21554_/X _23785_/Q _21549_/X VGND VGND VPWR VPWR _23785_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12294__A _12294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20506_ _20334_/A _20505_/X VGND VGND VPWR VPWR _20506_/X sky130_fd_sc_hd__or2_4
XANTENNA__22238__B2 _22234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21486_ _21256_/X _21485_/X _23822_/Q _21482_/X VGND VGND VPWR VPWR _21486_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24274_ _24240_/CLK _19337_/X HRESETn VGND VGND VPWR VPWR _24274_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20437_ _20231_/X _20423_/Y _20435_/X _20436_/Y _20255_/X VGND VGND VPWR VPWR _20438_/B
+ sky130_fd_sc_hd__a32o_4
X_23225_ _23641_/CLK _22531_/X VGND VGND VPWR VPWR _14753_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20368_ _20273_/X _20367_/X _24305_/Q _20349_/X VGND VGND VPWR VPWR _20368_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21461__A2 _21455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23156_ _23476_/CLK _22642_/X VGND VGND VPWR VPWR _11824_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20016__A _18670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22107_ _22105_/X _22099_/X _16476_/B _22106_/X VGND VGND VPWR VPWR _22107_/X sky130_fd_sc_hd__o22a_4
X_23087_ _18625_/X _19977_/X _24500_/Q _18625_/X VGND VGND VPWR VPWR _23087_/X sky130_fd_sc_hd__a2bb2o_4
X_20299_ _21526_/A VGND VGND VPWR VPWR _20299_/X sky130_fd_sc_hd__buf_2
XANTENNA__21213__A2 _21212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22038_ _11841_/B VGND VGND VPWR VPWR _22038_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14949__A _14663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13853__A _13853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14860_ _11895_/X VGND VGND VPWR VPWR _14881_/A sky130_fd_sc_hd__buf_2
XANTENNA__17325__A _15380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20972__A1 _20343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13811_ _13656_/A _13811_/B VGND VGND VPWR VPWR _13812_/C sky130_fd_sc_hd__or2_4
XFILLER_60_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14791_ _14675_/A _14717_/B VGND VGND VPWR VPWR _14792_/C sky130_fd_sc_hd__or2_4
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23989_ _23203_/CLK _23989_/D VGND VGND VPWR VPWR _23989_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12469__A _12469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18917__A1 _13266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22713__A2 _22708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16530_ _16527_/X _16529_/Y VGND VGND VPWR VPWR _16530_/Y sky130_fd_sc_hd__nor2_4
X_13742_ _13742_/A _23998_/Q VGND VGND VPWR VPWR _13743_/C sky130_fd_sc_hd__or2_4
XFILLER_56_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16461_ _16474_/A _16458_/X _16460_/X VGND VGND VPWR VPWR _16462_/C sky130_fd_sc_hd__and3_4
XFILLER_43_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23412__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13673_ _15411_/A _13673_/B _13673_/C VGND VGND VPWR VPWR _13673_/X sky130_fd_sc_hd__and3_4
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18200_ _17847_/A VGND VGND VPWR VPWR _18200_/X sky130_fd_sc_hd__buf_2
X_15412_ _15412_/A _15412_/B _15412_/C VGND VGND VPWR VPWR _15412_/X sky130_fd_sc_hd__or3_4
XANTENNA__17060__A _17060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12624_ _12973_/A _12520_/B VGND VGND VPWR VPWR _12624_/X sky130_fd_sc_hd__or2_4
X_19180_ _24331_/Q _19151_/X _19179_/Y VGND VGND VPWR VPWR _24331_/D sky130_fd_sc_hd__o21a_4
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16392_ _16011_/A _16390_/X _16391_/X VGND VGND VPWR VPWR _16392_/X sky130_fd_sc_hd__and3_4
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22477__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18131_ _17873_/X VGND VGND VPWR VPWR _18131_/X sky130_fd_sc_hd__buf_2
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15343_ _13704_/A _15343_/B VGND VGND VPWR VPWR _15343_/X sky130_fd_sc_hd__or2_4
X_12555_ _12511_/A _12668_/B VGND VGND VPWR VPWR _12555_/X sky130_fd_sc_hd__or2_4
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18062_ _18035_/X _18043_/Y _18056_/X _18059_/X _18061_/Y VGND VGND VPWR VPWR _18062_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15274_ _14165_/A _23928_/Q VGND VGND VPWR VPWR _15276_/B sky130_fd_sc_hd__or2_4
X_12486_ _13010_/A VGND VGND VPWR VPWR _12487_/A sky130_fd_sc_hd__buf_2
XFILLER_172_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12717__A1 _13339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17013_ _16939_/X VGND VGND VPWR VPWR _17013_/X sky130_fd_sc_hd__buf_2
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14225_ _14225_/A _23903_/Q VGND VGND VPWR VPWR _14228_/B sky130_fd_sc_hd__or2_4
XFILLER_171_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16404__A _12561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14156_ _14170_/A VGND VGND VPWR VPWR _14269_/A sky130_fd_sc_hd__buf_2
XANTENNA__12651__B _12548_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13107_ _13091_/A _13107_/B _13106_/X VGND VGND VPWR VPWR _13107_/X sky130_fd_sc_hd__or3_4
XANTENNA__20660__B1 _15702_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18964_ _18964_/A VGND VGND VPWR VPWR _18964_/Y sky130_fd_sc_hd__inv_2
X_14087_ _14086_/X VGND VGND VPWR VPWR _14088_/B sky130_fd_sc_hd__inv_2
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17408__A1 _13692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21204__A2 _21198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13038_ _11935_/A _13038_/B _13037_/X VGND VGND VPWR VPWR _13038_/X sky130_fd_sc_hd__or3_4
XANTENNA__22401__A1 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17408__B2 _17407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17915_ _18461_/A _17915_/B VGND VGND VPWR VPWR _17916_/D sky130_fd_sc_hd__and2_4
XANTENNA__22401__B2 _22366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18895_ _18894_/X VGND VGND VPWR VPWR _18896_/A sky130_fd_sc_hd__buf_2
XANTENNA__22141__A _20744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17846_ _17811_/X _17830_/X _17833_/X _17845_/Y VGND VGND VPWR VPWR _17846_/X sky130_fd_sc_hd__o22a_4
XFILLER_93_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12379__A _13529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17777_ _17673_/X _18013_/B _17671_/A _18013_/C VGND VGND VPWR VPWR _17777_/X sky130_fd_sc_hd__or4_4
XFILLER_47_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14989_ _15017_/A _23733_/Q VGND VGND VPWR VPWR _14990_/C sky130_fd_sc_hd__or2_4
XANTENNA__18908__A1 _16381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22704__A2 _22701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19516_ _19806_/A VGND VGND VPWR VPWR _19516_/X sky130_fd_sc_hd__buf_2
XANTENNA__19450__A _19450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16728_ _16724_/A _23857_/Q VGND VGND VPWR VPWR _16729_/C sky130_fd_sc_hd__or2_4
XFILLER_35_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16919__B1 _16911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24398__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18384__A2 _17188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16659_ _16659_/A _16657_/X _16658_/X VGND VGND VPWR VPWR _16660_/C sky130_fd_sc_hd__and3_4
X_19447_ _19438_/B VGND VGND VPWR VPWR _19447_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14594__A _15400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_54_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19378_ _18724_/X VGND VGND VPWR VPWR _19378_/Y sky130_fd_sc_hd__inv_2
X_18329_ _18307_/X _18328_/X _24487_/Q _18307_/X VGND VGND VPWR VPWR _24487_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13003__A _12506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21340_ _21266_/X _21334_/X _12809_/B _21338_/X VGND VGND VPWR VPWR _21340_/X sky130_fd_sc_hd__o22a_4
X_21271_ _20575_/A VGND VGND VPWR VPWR _21271_/X sky130_fd_sc_hd__buf_2
XANTENNA__12842__A _13566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16314__A _13377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23010_ _18325_/X _23003_/B VGND VGND VPWR VPWR _23010_/X sky130_fd_sc_hd__or2_4
X_20222_ _20221_/X VGND VGND VPWR VPWR _20772_/A sky130_fd_sc_hd__buf_2
XANTENNA__12184__A2 _12180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21443__A2 _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12561__B _12672_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20153_ _19906_/X _18628_/X _20152_/X VGND VGND VPWR VPWR _24134_/D sky130_fd_sc_hd__o21ai_4
XFILLER_170_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20084_ _24478_/Q VGND VGND VPWR VPWR _20084_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18886__D _17427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23912_ _23592_/CLK _21343_/X VGND VGND VPWR VPWR _13018_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18072__A1 _18022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17145__A _12419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21890__A _21923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23843_ _23939_/CLK _23843_/D VGND VGND VPWR VPWR _15827_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12289__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23774_ _23678_/CLK _21581_/X VGND VGND VPWR VPWR _13722_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _20863_/A _20984_/X _20985_/X VGND VGND VPWR VPWR _20986_/X sky130_fd_sc_hd__a21o_4
XPHY_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22725_ _20841_/A _22722_/X _13929_/B _22719_/X VGND VGND VPWR VPWR _23101_/D sky130_fd_sc_hd__o22a_4
XPHY_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16386__A1 _16309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11921__A _11891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22656_ _22432_/X _22651_/X _12548_/B _22655_/X VGND VGND VPWR VPWR _22656_/X sky130_fd_sc_hd__o22a_4
XFILLER_167_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21607_ _21607_/A VGND VGND VPWR VPWR _21608_/A sky130_fd_sc_hd__buf_2
XFILLER_22_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22587_ _21603_/A _22173_/B _21319_/A _22637_/D VGND VGND VPWR VPWR _22587_/X sky130_fd_sc_hd__or4_4
XFILLER_167_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21131__B2 _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12340_ _11712_/X _12204_/B VGND VGND VPWR VPWR _12340_/X sky130_fd_sc_hd__or2_4
X_24326_ _24287_/CLK _24326_/D HRESETn VGND VGND VPWR VPWR _19147_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21682__A2 _21677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21538_ _21536_/X _21530_/X _16395_/B _21537_/X VGND VGND VPWR VPWR _23792_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22226__A _22226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12271_ _12691_/A _12268_/X _12271_/C VGND VGND VPWR VPWR _12275_/B sky130_fd_sc_hd__and3_4
X_24257_ _24137_/CLK _24257_/D HRESETn VGND VGND VPWR VPWR _24257_/Q sky130_fd_sc_hd__dfrtp_4
X_21469_ _23828_/Q VGND VGND VPWR VPWR _21469_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14010_ _12233_/A _14008_/X _14010_/C VGND VGND VPWR VPWR _14011_/C sky130_fd_sc_hd__and3_4
X_23208_ _23496_/CLK _23208_/D VGND VGND VPWR VPWR _12995_/B sky130_fd_sc_hd__dfxtp_4
X_24188_ _23862_/CLK _19872_/Y HRESETn VGND VGND VPWR VPWR _22039_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22631__B2 _22626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23139_ _23303_/CLK _23139_/D VGND VGND VPWR VPWR _15826_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15961_ _15961_/A _15961_/B _15961_/C VGND VGND VPWR VPWR _15962_/C sky130_fd_sc_hd__and3_4
XFILLER_89_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17700_ _17699_/Y _17681_/X _17679_/A VGND VGND VPWR VPWR _17700_/X sky130_fd_sc_hd__a21o_4
X_14912_ _11659_/A _14912_/B VGND VGND VPWR VPWR _14915_/B sky130_fd_sc_hd__or2_4
XFILLER_62_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18063__B2 _18062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15892_ _13496_/A _15830_/B VGND VGND VPWR VPWR _15893_/C sky130_fd_sc_hd__or2_4
X_18680_ _17318_/A _18679_/B _17648_/X VGND VGND VPWR VPWR _18680_/X sky130_fd_sc_hd__o21a_4
XFILLER_48_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17631_ _17294_/X _17631_/B VGND VGND VPWR VPWR _17632_/D sky130_fd_sc_hd__nor2_4
X_14843_ _11666_/X _14811_/X _14843_/C VGND VGND VPWR VPWR _14843_/X sky130_fd_sc_hd__and3_4
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12199__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17562_ _17562_/A VGND VGND VPWR VPWR _18041_/B sky130_fd_sc_hd__inv_2
XFILLER_17_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23928__CLK _23864_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14774_ _15103_/A _14774_/B VGND VGND VPWR VPWR _14774_/X sky130_fd_sc_hd__or2_4
X_11986_ _16742_/A _21183_/A VGND VGND VPWR VPWR _11987_/C sky130_fd_sc_hd__or2_4
XFILLER_17_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16513_ _16481_/X _16436_/B VGND VGND VPWR VPWR _16514_/C sky130_fd_sc_hd__or2_4
X_19301_ _19236_/B VGND VGND VPWR VPWR _19301_/Y sky130_fd_sc_hd__inv_2
X_13725_ _15457_/A VGND VGND VPWR VPWR _13753_/A sky130_fd_sc_hd__buf_2
XFILLER_44_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21305__A _21238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17493_ _17493_/A _17492_/X VGND VGND VPWR VPWR _17493_/X sky130_fd_sc_hd__or2_4
XFILLER_147_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12927__A _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16444_ _11882_/X _16442_/X _16443_/X VGND VGND VPWR VPWR _16444_/X sky130_fd_sc_hd__and3_4
X_19232_ _24283_/Q _19231_/X VGND VGND VPWR VPWR _19233_/B sky130_fd_sc_hd__and2_4
XANTENNA__15303__A _14301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13656_ _13656_/A _23966_/Q VGND VGND VPWR VPWR _13657_/C sky130_fd_sc_hd__or2_4
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12646__B _12646_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12607_ _12623_/A VGND VGND VPWR VPWR _12646_/A sky130_fd_sc_hd__buf_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19163_ _19161_/A _19160_/X _20266_/A _19162_/Y VGND VGND VPWR VPWR _19163_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11550__B IRQ[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16375_ _16454_/A _16297_/B VGND VGND VPWR VPWR _16375_/X sky130_fd_sc_hd__or2_4
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13587_ _11928_/A VGND VGND VPWR VPWR _15029_/A sky130_fd_sc_hd__buf_2
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ _18037_/X _18114_/B VGND VGND VPWR VPWR _18119_/B sky130_fd_sc_hd__nor2_4
X_15326_ _15326_/A _24024_/Q VGND VGND VPWR VPWR _15326_/X sky130_fd_sc_hd__or2_4
X_12538_ _12905_/A VGND VGND VPWR VPWR _12894_/A sky130_fd_sc_hd__buf_2
XANTENNA__21673__A2 _21670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22870__A1 _17480_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19094_ _19094_/A VGND VGND VPWR VPWR _19094_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18045_ _17878_/A _17179_/X _17823_/A _17210_/X VGND VGND VPWR VPWR _18046_/A sky130_fd_sc_hd__o22a_4
XFILLER_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13758__A _12583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15257_ _15257_/A _23736_/Q VGND VGND VPWR VPWR _15258_/C sky130_fd_sc_hd__or2_4
X_12469_ _12469_/A VGND VGND VPWR VPWR _12470_/A sky130_fd_sc_hd__buf_2
X_14208_ _11708_/A VGND VGND VPWR VPWR _14254_/A sky130_fd_sc_hd__buf_2
X_15188_ _14771_/A _15188_/B _15188_/C VGND VGND VPWR VPWR _15188_/X sky130_fd_sc_hd__and3_4
XFILLER_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14139_ _14103_/A _14139_/B _14139_/C VGND VGND VPWR VPWR _14143_/B sky130_fd_sc_hd__and3_4
XFILLER_154_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19996_ _19992_/X _17780_/A _19956_/X _19995_/X VGND VGND VPWR VPWR _19997_/A sky130_fd_sc_hd__o22a_4
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18947_ _24370_/Q VGND VGND VPWR VPWR _18948_/C sky130_fd_sc_hd__inv_2
XANTENNA__22386__B1 _15466_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21189__B2 _21188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14589__A _14310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13493__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18878_ _18842_/A VGND VGND VPWR VPWR _18878_/X sky130_fd_sc_hd__buf_2
XFILLER_27_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17829_ _17828_/X VGND VGND VPWR VPWR _17829_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22138__B1 _15869_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14101__B _23199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20840_ _20840_/A VGND VGND VPWR VPWR _20841_/A sky130_fd_sc_hd__buf_2
XFILLER_130_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20771_ _20635_/X _20770_/X _24096_/Q _20746_/X VGND VGND VPWR VPWR _24096_/D sky130_fd_sc_hd__o22a_4
XFILLER_35_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21361__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22510_ _22440_/X _22508_/X _13035_/B _22505_/X VGND VGND VPWR VPWR _23240_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15213__A _14677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23490_ _23587_/CLK _23490_/D VGND VGND VPWR VPWR _15508_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12556__B _12669_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22441_ _22440_/X _22438_/X _12988_/B _22433_/X VGND VGND VPWR VPWR _23272_/D sky130_fd_sc_hd__o22a_4
XFILLER_149_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21113__B2 _21108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22372_ _22115_/X _22369_/X _12223_/B _22366_/X VGND VGND VPWR VPWR _22372_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21664__A2 _21663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22861__A1 _13049_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22046__A _22060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24111_ _23983_/CLK _24111_/D VGND VGND VPWR VPWR _16294_/B sky130_fd_sc_hd__dfxtp_4
X_21323_ _21338_/A VGND VGND VPWR VPWR _21331_/A sky130_fd_sc_hd__buf_2
XANTENNA__13668__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12572__A _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16044__A _11759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24233__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24042_ _24074_/CLK _24042_/D VGND VGND VPWR VPWR _24042_/Q sky130_fd_sc_hd__dfxtp_4
X_21254_ _21824_/A VGND VGND VPWR VPWR _21254_/X sky130_fd_sc_hd__buf_2
XANTENNA__21416__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22613__B2 _22612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15883__A _12402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20205_ _20205_/A VGND VGND VPWR VPWR _20205_/Y sky130_fd_sc_hd__inv_2
X_21185_ _21184_/X VGND VGND VPWR VPWR _21219_/A sky130_fd_sc_hd__buf_2
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20136_ _11566_/X _20134_/Y _20135_/Y VGND VGND VPWR VPWR _20136_/X sky130_fd_sc_hd__o21a_4
XFILLER_89_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11916__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24131__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20067_ _18475_/X _20055_/X _20065_/Y _20066_/X VGND VGND VPWR VPWR _20067_/X sky130_fd_sc_hd__o22a_4
XFILLER_58_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15107__B _23477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23826_ _23728_/CLK _23826_/D VGND VGND VPWR VPWR _23826_/Q sky130_fd_sc_hd__dfxtp_4
X_11840_ _11768_/X VGND VGND VPWR VPWR _12166_/A sky130_fd_sc_hd__buf_2
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21125__A _21118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23757_ _24045_/CLK _23757_/D VGND VGND VPWR VPWR _16102_/B sky130_fd_sc_hd__dfxtp_4
X_11771_ _16033_/A VGND VGND VPWR VPWR _16049_/A sky130_fd_sc_hd__buf_2
XPHY_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12747__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20969_ _20470_/A _20968_/X _19120_/A _18893_/A VGND VGND VPWR VPWR _20969_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24381__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16219__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13564_/A _13498_/X _13510_/C VGND VGND VPWR VPWR _13510_/X sky130_fd_sc_hd__and3_4
XANTENNA__15123__A _11898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11651__A _15321_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22708_ _22708_/A VGND VGND VPWR VPWR _22708_/X sky130_fd_sc_hd__buf_2
XFILLER_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14490_ _14513_/A _14490_/B _14490_/C VGND VGND VPWR VPWR _14490_/X sky130_fd_sc_hd__or3_4
XPHY_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23688_ _23337_/CLK _23688_/D VGND VGND VPWR VPWR _23688_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _13441_/A _22337_/A VGND VGND VPWR VPWR _13444_/B sky130_fd_sc_hd__or2_4
XFILLER_158_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22639_ _22672_/A VGND VGND VPWR VPWR _22655_/A sky130_fd_sc_hd__inv_2
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15582__A2 _11629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16160_ _16160_/A _16159_/X VGND VGND VPWR VPWR _16160_/X sky130_fd_sc_hd__and2_4
X_13372_ _13413_/A _13372_/B _13372_/C VGND VGND VPWR VPWR _13373_/C sky130_fd_sc_hd__and3_4
XFILLER_107_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15111_ _15080_/A _23637_/Q VGND VGND VPWR VPWR _15112_/C sky130_fd_sc_hd__or2_4
X_12323_ _13052_/A VGND VGND VPWR VPWR _13230_/A sky130_fd_sc_hd__buf_2
XFILLER_126_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24309_ _24342_/CLK _24309_/D HRESETn VGND VGND VPWR VPWR _24309_/Q sky130_fd_sc_hd__dfrtp_4
X_16091_ _15969_/A _16167_/B VGND VGND VPWR VPWR _16091_/X sky130_fd_sc_hd__or2_4
XFILLER_6_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15042_ _12233_/A _15042_/B _15041_/X VGND VGND VPWR VPWR _15043_/C sky130_fd_sc_hd__and3_4
X_12254_ _12269_/A _23596_/Q VGND VGND VPWR VPWR _12255_/C sky130_fd_sc_hd__or2_4
XANTENNA__18808__B1 _11573_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21407__A2 _21405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22604__B2 _22598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15793__A _12848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19850_ _19767_/A _19712_/B _19507_/B _19849_/X VGND VGND VPWR VPWR _19850_/X sky130_fd_sc_hd__a211o_4
X_12185_ _13046_/A VGND VGND VPWR VPWR _12912_/A sky130_fd_sc_hd__buf_2
XANTENNA__22080__A2 _22074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18801_ _12419_/X _18796_/X _24460_/Q _18797_/X VGND VGND VPWR VPWR _18801_/X sky130_fd_sc_hd__o22a_4
X_19781_ _19781_/A _19787_/A _19780_/X VGND VGND VPWR VPWR _19781_/X sky130_fd_sc_hd__or3_4
X_16993_ _17667_/A _18107_/A VGND VGND VPWR VPWR _16994_/B sky130_fd_sc_hd__or2_4
XFILLER_89_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11826__A _11705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18732_ _18518_/A _17341_/A VGND VGND VPWR VPWR _18732_/X sky130_fd_sc_hd__and2_4
X_15944_ _15944_/A _23374_/Q VGND VGND VPWR VPWR _15946_/B sky130_fd_sc_hd__or2_4
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23750__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21711__A2_N _21710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11545__B IRQ[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15875_ _13543_/X _23331_/Q VGND VGND VPWR VPWR _15877_/B sky130_fd_sc_hd__or2_4
X_18663_ _17013_/X _18658_/Y _16943_/A _18662_/X VGND VGND VPWR VPWR _18663_/X sky130_fd_sc_hd__o22a_4
XFILLER_49_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15017__B _23957_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21591__A1 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21591__B2 _21585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17614_ _17429_/X _17613_/Y _17423_/B _17433_/Y VGND VGND VPWR VPWR _17614_/X sky130_fd_sc_hd__a211o_4
X_14826_ _14682_/A _14826_/B _14825_/X VGND VGND VPWR VPWR _14826_/X sky130_fd_sc_hd__and3_4
X_18594_ _18574_/X _18593_/X _20088_/A _18574_/X VGND VGND VPWR VPWR _24477_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13760__B _13760_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21035__A _21042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17545_ _17452_/X _17528_/Y _17536_/Y _17544_/Y VGND VGND VPWR VPWR _17545_/X sky130_fd_sc_hd__a211o_4
X_14757_ _12495_/A _14827_/B VGND VGND VPWR VPWR _14757_/X sky130_fd_sc_hd__or2_4
XANTENNA__12657__A _12943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11969_ _11969_/A VGND VGND VPWR VPWR _11970_/A sky130_fd_sc_hd__buf_2
XANTENNA__21343__B2 _21338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13708_ _14543_/A _13702_/X _13708_/C VGND VGND VPWR VPWR _13708_/X sky130_fd_sc_hd__and3_4
X_17476_ _17640_/A VGND VGND VPWR VPWR _18154_/B sky130_fd_sc_hd__inv_2
X_14688_ _15620_/A _14688_/B VGND VGND VPWR VPWR _14689_/C sky130_fd_sc_hd__or2_4
XFILLER_20_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19215_ _19215_/A VGND VGND VPWR VPWR _19215_/Y sky130_fd_sc_hd__inv_2
X_16427_ _16129_/A _16423_/X _16426_/X VGND VGND VPWR VPWR _16427_/X sky130_fd_sc_hd__or3_4
X_13639_ _13639_/A _23550_/Q VGND VGND VPWR VPWR _13640_/C sky130_fd_sc_hd__or2_4
XFILLER_60_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24256__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13584__A1 _13485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16358_ _16342_/A _16290_/B VGND VGND VPWR VPWR _16358_/X sky130_fd_sc_hd__or2_4
X_19146_ _24325_/Q _19145_/X VGND VGND VPWR VPWR _19146_/X sky130_fd_sc_hd__and2_4
XFILLER_34_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21646__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15309_ _15018_/A _15309_/B _15308_/X VGND VGND VPWR VPWR _15310_/C sky130_fd_sc_hd__and3_4
X_16289_ _11890_/X _16289_/B VGND VGND VPWR VPWR _16289_/X sky130_fd_sc_hd__or2_4
X_19077_ _19075_/Y _19076_/Y _11525_/X VGND VGND VPWR VPWR _19077_/X sky130_fd_sc_hd__o21a_4
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18028_ _16995_/B VGND VGND VPWR VPWR _18028_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19979_ _19951_/X VGND VGND VPWR VPWR _19979_/X sky130_fd_sc_hd__buf_2
XFILLER_45_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11736__A _11736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15208__A _14635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22990_ _22922_/A _22990_/B _22990_/C VGND VGND VPWR VPWR _22990_/X sky130_fd_sc_hd__or3_4
XFILLER_80_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19775__A1 _19773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21941_ _21941_/A VGND VGND VPWR VPWR _21957_/A sky130_fd_sc_hd__inv_2
XFILLER_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17786__B1 _17653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21872_ _20892_/A VGND VGND VPWR VPWR _21872_/X sky130_fd_sc_hd__buf_2
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _23323_/CLK _23611_/D VGND VGND VPWR VPWR _14455_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _20664_/A _20821_/X _20822_/X VGND VGND VPWR VPWR _20824_/B sky130_fd_sc_hd__and3_4
XFILLER_23_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12567__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23542_ _23511_/CLK _23542_/D VGND VGND VPWR VPWR _14946_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20754_ _20754_/A VGND VGND VPWR VPWR _20754_/X sky130_fd_sc_hd__buf_2
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23473_ _23409_/CLK _22104_/X VGND VGND VPWR VPWR _16776_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_24_0_HCLK clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20685_ _20501_/A _20685_/B VGND VGND VPWR VPWR _20685_/Y sky130_fd_sc_hd__nor2_4
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14782__A _15106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22424_ _22423_/X _22414_/X _16247_/B _22421_/X VGND VGND VPWR VPWR _22424_/X sky130_fd_sc_hd__o22a_4
XFILLER_109_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21637__A2 _21634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13398__A _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22355_ _22090_/A _21656_/B _21319_/A _21030_/A VGND VGND VPWR VPWR _22355_/X sky130_fd_sc_hd__or4_4
XFILLER_152_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21306_ _21304_/X _21305_/X _14644_/B _21300_/X VGND VGND VPWR VPWR _21306_/X sky130_fd_sc_hd__o22a_4
X_22286_ _22108_/X _22280_/X _16251_/B _22284_/X VGND VGND VPWR VPWR _22286_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24025_ _24057_/CLK _21127_/X VGND VGND VPWR VPWR _14716_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22062__A2 _22060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21237_ _21236_/X VGND VGND VPWR VPWR _21238_/A sky130_fd_sc_hd__buf_2
XFILLER_104_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21168_ _20770_/X _21162_/X _24000_/Q _21166_/X VGND VGND VPWR VPWR _24000_/D sky130_fd_sc_hd__o22a_4
XFILLER_46_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11646__A _11646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15118__A _14983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20119_ _20119_/A VGND VGND VPWR VPWR _20119_/Y sky130_fd_sc_hd__inv_2
X_21099_ _20464_/X _21097_/X _24045_/Q _21094_/X VGND VGND VPWR VPWR _21099_/X sky130_fd_sc_hd__o22a_4
X_13990_ _13990_/A _23136_/Q VGND VGND VPWR VPWR _13990_/X sky130_fd_sc_hd__or2_4
XANTENNA__14022__A _13705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12941_ _12941_/A _12939_/X _12941_/C VGND VGND VPWR VPWR _12941_/X sky130_fd_sc_hd__and3_4
XANTENNA__24129__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20376__A2 _20304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13861__A _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15660_ _12689_/A _15660_/B VGND VGND VPWR VPWR _15660_/X sky130_fd_sc_hd__or2_4
XANTENNA__17333__A _15251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12872_ _12872_/A _23561_/Q VGND VGND VPWR VPWR _12872_/X sky130_fd_sc_hd__or2_4
XFILLER_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18148__B _18148_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14611_ _15450_/A _14610_/X VGND VGND VPWR VPWR _14611_/X sky130_fd_sc_hd__and2_4
X_11823_ _12138_/A _11819_/X _11822_/X VGND VGND VPWR VPWR _11823_/X sky130_fd_sc_hd__or3_4
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23809_ _23744_/CLK _23809_/D VGND VGND VPWR VPWR _15574_/B sky130_fd_sc_hd__dfxtp_4
X_15591_ _15616_/A _15585_/X _15591_/C VGND VGND VPWR VPWR _15591_/X sky130_fd_sc_hd__or3_4
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__A _12477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21325__B2 _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23153__CLK _23281_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24279__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17330_ _17327_/Y _17018_/X _17025_/Y _17329_/X VGND VGND VPWR VPWR _17332_/B sky130_fd_sc_hd__o22a_4
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _13751_/A _14470_/B VGND VGND VPWR VPWR _14543_/C sky130_fd_sc_hd__or2_4
XFILLER_14_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _12596_/A VGND VGND VPWR VPWR _13063_/A sky130_fd_sc_hd__buf_2
XANTENNA__21876__A2 _21875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17261_ _16821_/A VGND VGND VPWR VPWR _17261_/Y sky130_fd_sc_hd__inv_2
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _15395_/A _14531_/B VGND VGND VPWR VPWR _14473_/X sky130_fd_sc_hd__or2_4
X_11685_ _11684_/X VGND VGND VPWR VPWR _16187_/A sky130_fd_sc_hd__buf_2
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16212_ _16231_/A _24077_/Q VGND VGND VPWR VPWR _16213_/C sky130_fd_sc_hd__or2_4
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19000_ _11538_/A _11538_/B _18995_/Y VGND VGND VPWR VPWR _19000_/Y sky130_fd_sc_hd__a21oi_4
X_13424_ _13327_/A _13422_/X _13424_/C VGND VGND VPWR VPWR _13424_/X sky130_fd_sc_hd__and3_4
XANTENNA__21628__A2 _21627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17192_ _17197_/A VGND VGND VPWR VPWR _17192_/X sky130_fd_sc_hd__buf_2
X_16143_ _16147_/A _16219_/B VGND VGND VPWR VPWR _16143_/X sky130_fd_sc_hd__or2_4
X_13355_ _13399_/A _13348_/X _13355_/C VGND VGND VPWR VPWR _13363_/B sky130_fd_sc_hd__or3_4
XFILLER_128_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ _13333_/A _23660_/Q VGND VGND VPWR VPWR _12307_/C sky130_fd_sc_hd__or2_4
XANTENNA__13101__A _13094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16074_ _16066_/A _16072_/X _16074_/C VGND VGND VPWR VPWR _16074_/X sky130_fd_sc_hd__and3_4
XFILLER_155_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13286_ _13309_/A _13286_/B VGND VGND VPWR VPWR _13288_/B sky130_fd_sc_hd__or2_4
XFILLER_136_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22414__A _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19902_ _19890_/A _19741_/B VGND VGND VPWR VPWR _19902_/X sky130_fd_sc_hd__or2_4
X_15025_ _13965_/A _15023_/X _15025_/C VGND VGND VPWR VPWR _15025_/X sky130_fd_sc_hd__and3_4
X_12237_ _12748_/A VGND VGND VPWR VPWR _12298_/A sky130_fd_sc_hd__buf_2
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_44_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR _23662_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19833_ _19687_/A _19832_/X _19815_/B VGND VGND VPWR VPWR _19833_/X sky130_fd_sc_hd__o21a_4
X_12168_ _12168_/A _12168_/B _12168_/C VGND VGND VPWR VPWR _12169_/C sky130_fd_sc_hd__and3_4
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19764_ _19823_/A _19763_/Y VGND VGND VPWR VPWR _19765_/B sky130_fd_sc_hd__or2_4
X_16976_ _17732_/A _16975_/X VGND VGND VPWR VPWR _16976_/X sky130_fd_sc_hd__or2_4
X_12099_ _12064_/X _23667_/Q VGND VGND VPWR VPWR _12100_/C sky130_fd_sc_hd__or2_4
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18715_ _17333_/X _18713_/X _18506_/A _18714_/X VGND VGND VPWR VPWR _18716_/A sky130_fd_sc_hd__a211o_4
X_15927_ _15914_/X VGND VGND VPWR VPWR _15927_/Y sky130_fd_sc_hd__inv_2
X_19695_ _19797_/A _19691_/Y _19895_/A _19694_/X VGND VGND VPWR VPWR _19695_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21564__B2 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18646_ _18622_/Y _18624_/X _18625_/X _18645_/X VGND VGND VPWR VPWR _18646_/X sky130_fd_sc_hd__o22a_4
XFILLER_65_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15858_ _15851_/A _15797_/B VGND VGND VPWR VPWR _15858_/X sky130_fd_sc_hd__or2_4
XFILLER_149_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14809_ _14660_/A _14809_/B _14809_/C VGND VGND VPWR VPWR _14810_/C sky130_fd_sc_hd__or3_4
XFILLER_80_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18577_ _16975_/X _18698_/B VGND VGND VPWR VPWR _18577_/X sky130_fd_sc_hd__or2_4
XFILLER_75_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15789_ _11888_/A _15789_/B VGND VGND VPWR VPWR _15789_/X sky130_fd_sc_hd__or2_4
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21316__B2 _21239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17528_ _17528_/A _17527_/X VGND VGND VPWR VPWR _17528_/Y sky130_fd_sc_hd__nor2_4
XFILLER_75_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15698__A _13145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17459_ _17459_/A VGND VGND VPWR VPWR _17459_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18074__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21619__A2 _21613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20470_ _20470_/A VGND VGND VPWR VPWR _20470_/X sky130_fd_sc_hd__buf_2
XFILLER_119_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19129_ _19129_/A VGND VGND VPWR VPWR _24341_/D sky130_fd_sc_hd__inv_2
XANTENNA__15210__B _15139_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22292__A2 _22287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14107__A _12287_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22140_ _22139_/X _22135_/X _15474_/B _22130_/X VGND VGND VPWR VPWR _23458_/D sky130_fd_sc_hd__o22a_4
XFILLER_134_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13946__A _13945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22071_ _22057_/A VGND VGND VPWR VPWR _22071_/X sky130_fd_sc_hd__buf_2
XANTENNA__17418__A _17418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12850__A _12236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19996__A1 _19992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21022_ _24213_/Q _20358_/A _21021_/Y VGND VGND VPWR VPWR _22169_/A sky130_fd_sc_hd__o21a_4
XFILLER_113_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_1_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22973_ _18494_/X _22973_/B VGND VGND VPWR VPWR _22974_/C sky130_fd_sc_hd__or2_4
XANTENNA__14777__A _15080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21555__B2 _21549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13681__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17153__A _17153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21924_ _21862_/X _21923_/X _23583_/Q _21920_/X VGND VGND VPWR VPWR _23583_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22994__A _22993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21855_ _21570_/A VGND VGND VPWR VPWR _21855_/X sky130_fd_sc_hd__buf_2
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12297__A _13145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _20641_/X _20805_/X _20639_/X VGND VGND VPWR VPWR _20806_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21786_ _21568_/X _21784_/X _15837_/B _21781_/X VGND VGND VPWR VPWR _21786_/X sky130_fd_sc_hd__o22a_4
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23525_ _23493_/CLK _23525_/D VGND VGND VPWR VPWR _13420_/B sky130_fd_sc_hd__dfxtp_4
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20737_ _20930_/A _20736_/X VGND VGND VPWR VPWR _20737_/Y sky130_fd_sc_hd__nor2_4
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15401__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23456_ _23456_/CLK _23456_/D VGND VGND VPWR VPWR _14039_/B sky130_fd_sc_hd__dfxtp_4
X_20668_ _20668_/A VGND VGND VPWR VPWR _20697_/A sky130_fd_sc_hd__buf_2
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22407_ _22462_/A VGND VGND VPWR VPWR _22433_/A sky130_fd_sc_hd__inv_2
XFILLER_52_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23387_ _23772_/CLK _23387_/D VGND VGND VPWR VPWR _14462_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22283__A2 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20599_ _20251_/A _20598_/X _20306_/X VGND VGND VPWR VPWR _20599_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__14017__A _15369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20961__B _19773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13140_ _13170_/A _13140_/B _13139_/X VGND VGND VPWR VPWR _13141_/C sky130_fd_sc_hd__and3_4
XFILLER_104_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22338_ _15746_/B VGND VGND VPWR VPWR _23332_/D sky130_fd_sc_hd__buf_2
XFILLER_87_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22234__A _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13856__A _11878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13071_ _13103_/A _13071_/B _13070_/X VGND VGND VPWR VPWR _13072_/C sky130_fd_sc_hd__and3_4
XANTENNA__18239__B2 _18238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22035__A2 _22031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17328__A _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22269_ _22165_/X _22265_/X _15165_/B _22226_/X VGND VGND VPWR VPWR _22269_/X sky130_fd_sc_hd__o22a_4
XFILLER_3_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24008_ _24073_/CLK _24008_/D VGND VGND VPWR VPWR _24008_/Q sky130_fd_sc_hd__dfxtp_4
X_12022_ _11851_/X _12021_/Y VGND VGND VPWR VPWR _12025_/A sky130_fd_sc_hd__and2_4
XFILLER_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21794__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22888__B _22887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16830_ _15931_/D VGND VGND VPWR VPWR _16830_/X sky130_fd_sc_hd__buf_2
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16761_ _16788_/A _16761_/B VGND VGND VPWR VPWR _16761_/X sky130_fd_sc_hd__or2_4
XFILLER_65_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13973_ _13663_/A _13973_/B _13973_/C VGND VGND VPWR VPWR _13973_/X sky130_fd_sc_hd__or3_4
XANTENNA__14687__A _15606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18500_ _18500_/A _18364_/X VGND VGND VPWR VPWR _18500_/Y sky130_fd_sc_hd__nand2_4
X_12924_ _12950_/A _12924_/B _12923_/X VGND VGND VPWR VPWR _12924_/X sky130_fd_sc_hd__and3_4
X_15712_ _12747_/A _15712_/B VGND VGND VPWR VPWR _15712_/X sky130_fd_sc_hd__or2_4
XFILLER_4_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17063__A _11595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19480_ _19480_/A VGND VGND VPWR VPWR _19480_/X sky130_fd_sc_hd__buf_2
X_16692_ _16702_/A _16692_/B _16692_/C VGND VGND VPWR VPWR _16692_/X sky130_fd_sc_hd__and3_4
XFILLER_61_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18431_ _18400_/X _18430_/X _24484_/Q _18400_/X VGND VGND VPWR VPWR _24484_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23669__CLK _23456_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12855_ _12860_/A _12919_/B VGND VGND VPWR VPWR _12855_/X sky130_fd_sc_hd__or2_4
X_15643_ _13886_/A _15641_/X _15643_/C VGND VGND VPWR VPWR _15643_/X sky130_fd_sc_hd__and3_4
XFILLER_146_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11806_ _16647_/A _11804_/X _11805_/X VGND VGND VPWR VPWR _11807_/C sky130_fd_sc_hd__and3_4
XFILLER_33_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21849__A2 _21839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18362_ _17726_/A VGND VGND VPWR VPWR _18553_/A sky130_fd_sc_hd__buf_2
X_15574_ _14421_/A _15574_/B VGND VGND VPWR VPWR _15574_/X sky130_fd_sc_hd__or2_4
X_12786_ _13343_/A _12782_/X _12786_/C VGND VGND VPWR VPWR _12786_/X sky130_fd_sc_hd__and3_4
XANTENNA__12000__A _16148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19911__A1 _19906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22409__A _22421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _12410_/A _14523_/X _14525_/C VGND VGND VPWR VPWR _14525_/X sky130_fd_sc_hd__and3_4
XANTENNA__21313__A _21313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17313_ _17304_/X VGND VGND VPWR VPWR _17351_/B sky130_fd_sc_hd__inv_2
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _12634_/A VGND VGND VPWR VPWR _13232_/A sky130_fd_sc_hd__buf_2
XANTENNA__19430__A2_N _18682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18293_ _18169_/Y _17499_/Y _17530_/Y VGND VGND VPWR VPWR _18293_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12935__A _12942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16407__A _15998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15311__A _13853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14456_ _12455_/A _24059_/Q VGND VGND VPWR VPWR _14457_/C sky130_fd_sc_hd__or2_4
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17244_ _12027_/X _17240_/B VGND VGND VPWR VPWR _17245_/A sky130_fd_sc_hd__or2_4
X_11668_ _11668_/A VGND VGND VPWR VPWR _12979_/A sky130_fd_sc_hd__buf_2
XFILLER_168_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _13407_/A _13407_/B _13407_/C VGND VGND VPWR VPWR _13415_/B sky130_fd_sc_hd__or3_4
XANTENNA__24234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15030__B _23477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17175_ _17160_/X _17171_/X _17838_/A _17174_/X VGND VGND VPWR VPWR _17175_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14387_ _14506_/A _14387_/B VGND VGND VPWR VPWR _14387_/X sky130_fd_sc_hd__or2_4
X_11599_ _17357_/A VGND VGND VPWR VPWR _17048_/A sky130_fd_sc_hd__buf_2
X_16126_ _16099_/X VGND VGND VPWR VPWR _16157_/A sky130_fd_sc_hd__buf_2
XFILLER_6_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13338_ _13338_/A _13334_/X _13338_/C VGND VGND VPWR VPWR _13339_/B sky130_fd_sc_hd__or3_4
XFILLER_128_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22144__A _22459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16057_ _16057_/A _16057_/B VGND VGND VPWR VPWR _16059_/B sky130_fd_sc_hd__or2_4
XANTENNA__22026__A2 _22024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13269_ _13269_/A _13269_/B VGND VGND VPWR VPWR _13269_/X sky130_fd_sc_hd__or2_4
XFILLER_142_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15008_ _12450_/X _23573_/Q VGND VGND VPWR VPWR _15009_/C sky130_fd_sc_hd__or2_4
XFILLER_116_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21785__B2 _21781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19816_ _19749_/X _19816_/B VGND VGND VPWR VPWR _19816_/X sky130_fd_sc_hd__and2_4
XFILLER_116_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19747_ _19848_/B VGND VGND VPWR VPWR _19748_/C sky130_fd_sc_hd__inv_2
XFILLER_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16959_ _24147_/Q VGND VGND VPWR VPWR _17905_/A sky130_fd_sc_hd__inv_2
XFILLER_42_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14597__A _12477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19678_ _19681_/A _19678_/B VGND VGND VPWR VPWR _19678_/X sky130_fd_sc_hd__and2_4
XFILLER_37_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18629_ _18698_/B VGND VGND VPWR VPWR _18630_/C sky130_fd_sc_hd__inv_2
XANTENNA__13006__A _12513_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21640_ _21575_/X _21634_/X _23744_/Q _21638_/X VGND VGND VPWR VPWR _23744_/D sky130_fd_sc_hd__o22a_4
XFILLER_162_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21223__A _21202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21571_ _21570_/X _21566_/X _23778_/Q _21561_/X VGND VGND VPWR VPWR _23778_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17420__B _17421_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16317__A _11727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23310_ _23438_/CLK _23310_/D VGND VGND VPWR VPWR _23310_/Q sky130_fd_sc_hd__dfxtp_4
X_20522_ _20352_/A VGND VGND VPWR VPWR _20522_/X sky130_fd_sc_hd__buf_2
XFILLER_123_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24290_ _24388_/CLK _24290_/D HRESETn VGND VGND VPWR VPWR _24290_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12564__B _12564_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23241_ _23241_/CLK _22509_/X VGND VGND VPWR VPWR _23241_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18469__A1 _18413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20453_ _20273_/A _20452_/Y _19250_/A _20323_/X VGND VGND VPWR VPWR _20453_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13950__A1 _13863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23172_ _23204_/CLK _22616_/X VGND VGND VPWR VPWR _15737_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_107_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20384_ _20277_/X _20383_/X _24400_/Q _18894_/B VGND VGND VPWR VPWR _20384_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17141__A1 _14549_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13676__A _13676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22123_ _22123_/A VGND VGND VPWR VPWR _22123_/X sky130_fd_sc_hd__buf_2
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17692__A2 _17520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16052__A _16222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12580__A _12580_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22989__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22054_ _21826_/X _22053_/X _16076_/B _22050_/X VGND VGND VPWR VPWR _23502_/D sky130_fd_sc_hd__o22a_4
XFILLER_99_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21776__B2 _21774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21005_ _20894_/X _21004_/X _14895_/B _20396_/A VGND VGND VPWR VPWR _24086_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_7_90_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR _23582_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_75_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20302__A _20533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11924__A _11905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22956_ _22947_/X _22954_/Y _22955_/X VGND VGND VPWR VPWR _22956_/X sky130_fd_sc_hd__and3_4
XANTENNA__14300__A _12469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21907_ _21833_/X _21902_/X _12619_/B _21906_/X VGND VGND VPWR VPWR _21907_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22887_ _17556_/Y _22885_/X _22875_/X _22886_/X VGND VGND VPWR VPWR _22887_/X sky130_fd_sc_hd__o22a_4
X_12640_ _12962_/A _12640_/B _12640_/C VGND VGND VPWR VPWR _12641_/C sky130_fd_sc_hd__and3_4
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21838_ _21268_/A VGND VGND VPWR VPWR _21838_/X sky130_fd_sc_hd__buf_2
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22229__A _22258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21133__A _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12571_ _12571_/A _12571_/B _12570_/X VGND VGND VPWR VPWR _12571_/X sky130_fd_sc_hd__or3_4
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12755__A _12975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21769_ _21539_/X _21763_/X _16297_/B _21767_/X VGND VGND VPWR VPWR _21769_/X sky130_fd_sc_hd__o22a_4
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16227__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _14310_/A _14310_/B _14310_/C VGND VGND VPWR VPWR _14310_/X sky130_fd_sc_hd__or3_4
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21700__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23508_ _23668_/CLK _23508_/D VGND VGND VPWR VPWR _11841_/B sky130_fd_sc_hd__dfxtp_4
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ _11522_/A _11521_/X VGND VGND VPWR VPWR _11523_/B sky130_fd_sc_hd__or2_4
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15290_ _14154_/A _23128_/Q VGND VGND VPWR VPWR _15290_/X sky130_fd_sc_hd__or2_4
XFILLER_8_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24488_ _24294_/CLK _24488_/D HRESETn VGND VGND VPWR VPWR _20036_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17380__A1 _16611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24317__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14241_ _14656_/A _14239_/X _14240_/X VGND VGND VPWR VPWR _14241_/X sky130_fd_sc_hd__and3_4
X_23439_ _23983_/CLK _23439_/D VGND VGND VPWR VPWR _16290_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22256__A2 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14172_ _14991_/A _14167_/X _14172_/C VGND VGND VPWR VPWR _14172_/X sky130_fd_sc_hd__or3_4
XANTENNA__15785__B _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13123_ _13123_/A _13123_/B _13122_/X VGND VGND VPWR VPWR _13124_/C sky130_fd_sc_hd__and3_4
XFILLER_124_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13586__A _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22008__A2 _22003_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17058__A _17017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12490__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18980_ _24367_/Q VGND VGND VPWR VPWR _18980_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18880__A1 _17290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13054_ _13094_/A _12988_/B VGND VGND VPWR VPWR _13054_/X sky130_fd_sc_hd__or2_4
X_17931_ _17811_/X _17925_/X _17833_/X _17930_/Y VGND VGND VPWR VPWR _17931_/X sky130_fd_sc_hd__o22a_4
XFILLER_3_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12005_ _12106_/A _24116_/Q VGND VGND VPWR VPWR _12006_/C sky130_fd_sc_hd__or2_4
X_17862_ _17922_/A _17860_/X _17814_/X _17861_/X VGND VGND VPWR VPWR _17862_/X sky130_fd_sc_hd__o22a_4
XFILLER_87_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19601_ _19582_/X _19601_/B _19597_/X _19600_/X VGND VGND VPWR VPWR _19601_/X sky130_fd_sc_hd__or4_4
XFILLER_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16813_ _16621_/A _16813_/B VGND VGND VPWR VPWR _16813_/X sky130_fd_sc_hd__or2_4
XFILLER_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20212__A _24129_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17793_ _17792_/X VGND VGND VPWR VPWR _17793_/X sky130_fd_sc_hd__buf_2
XANTENNA__21519__B2 _21482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19532_ _19532_/A VGND VGND VPWR VPWR _19533_/B sky130_fd_sc_hd__inv_2
XANTENNA__15306__A _14897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16744_ _16744_/A _23729_/Q VGND VGND VPWR VPWR _16746_/B sky130_fd_sc_hd__or2_4
X_13956_ _13983_/A _23360_/Q VGND VGND VPWR VPWR _13956_/X sky130_fd_sc_hd__or2_4
XANTENNA__17199__A1 _16821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22192__B2 _22191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12907_ _12472_/A _12907_/B _12907_/C VGND VGND VPWR VPWR _12907_/X sky130_fd_sc_hd__and3_4
X_19463_ _19506_/A VGND VGND VPWR VPWR _19839_/A sky130_fd_sc_hd__buf_2
XFILLER_98_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16675_ _16675_/A _16671_/X _16675_/C VGND VGND VPWR VPWR _16683_/B sky130_fd_sc_hd__or3_4
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13887_ _15595_/A VGND VGND VPWR VPWR _14385_/A sky130_fd_sc_hd__buf_2
XANTENNA__20866__B _20866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18414_ _17636_/B _17616_/B VGND VGND VPWR VPWR _18415_/C sky130_fd_sc_hd__and2_4
X_12838_ _13367_/A _12836_/X _12838_/C VGND VGND VPWR VPWR _12839_/C sky130_fd_sc_hd__and3_4
XANTENNA__24486__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15626_ _11710_/A _15559_/B VGND VGND VPWR VPWR _15628_/B sky130_fd_sc_hd__or2_4
X_19394_ _19392_/X _18031_/Y _19392_/X _24239_/Q VGND VGND VPWR VPWR _19394_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22139__A _20718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18345_ _17497_/X _17638_/Y VGND VGND VPWR VPWR _18345_/X sky130_fd_sc_hd__or2_4
XANTENNA__24415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ _12775_/A _23754_/Q VGND VGND VPWR VPWR _12769_/X sky130_fd_sc_hd__or2_4
X_15557_ _14418_/X _15555_/X _15557_/C VGND VGND VPWR VPWR _15557_/X sky130_fd_sc_hd__and3_4
XANTENNA__22495__A2 _22494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16137__A _16110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508_ _14520_/A _23995_/Q VGND VGND VPWR VPWR _14509_/C sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_2_1_0_HCLK_A clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15488_ _13774_/A _15488_/B _15487_/X VGND VGND VPWR VPWR _15488_/X sky130_fd_sc_hd__and3_4
X_18276_ _18244_/X _18275_/X _24489_/Q _18244_/X VGND VGND VPWR VPWR _24489_/D sky130_fd_sc_hd__a2bb2o_4
X_17227_ _17151_/X VGND VGND VPWR VPWR _17227_/X sky130_fd_sc_hd__buf_2
X_14439_ _12537_/A _23323_/Q VGND VGND VPWR VPWR _14441_/B sky130_fd_sc_hd__or2_4
XANTENNA__22247__A2 _22244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17158_ _17130_/X _17154_/X _17124_/X _17157_/X VGND VGND VPWR VPWR _17158_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24358__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16109_ _16109_/A _23309_/Q VGND VGND VPWR VPWR _16110_/C sky130_fd_sc_hd__or2_4
XFILLER_115_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17089_ _17089_/A _17912_/A VGND VGND VPWR VPWR _17089_/X sky130_fd_sc_hd__and2_4
XFILLER_157_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_14_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14104__B _24031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19820__B1 _16915_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16600__A _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11744__A _16079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22810_ _17284_/Y _22803_/X VGND VGND VPWR VPWR HWDATA[5] sky130_fd_sc_hd__nor2_4
XANTENNA__15216__A _14615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23790_ _23662_/CLK _23790_/D VGND VGND VPWR VPWR _23790_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14120__A _14131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12559__B _12671_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22183__B2 _22177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22741_ _23048_/A VGND VGND VPWR VPWR _22742_/A sky130_fd_sc_hd__buf_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_1_HCLK clkbuf_1_0_1_HCLK/A VGND VGND VPWR VPWR clkbuf_2_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__18527__A _18064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17431__A _17429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22672_ _22672_/A VGND VGND VPWR VPWR _22672_/X sky130_fd_sc_hd__buf_2
XANTENNA__18139__B1 _17648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24411_ _24445_/CLK _24411_/D HRESETn VGND VGND VPWR VPWR _24411_/Q sky130_fd_sc_hd__dfrtp_4
X_21623_ _21546_/X _21620_/X _23756_/Q _21617_/X VGND VGND VPWR VPWR _23756_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12575__A _11681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16047__A _16047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24342_ _24342_/CLK _24342_/D HRESETn VGND VGND VPWR VPWR _24342_/Q sky130_fd_sc_hd__dfstp_4
X_21554_ _21542_/A VGND VGND VPWR VPWR _21554_/X sky130_fd_sc_hd__buf_2
XFILLER_139_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20505_ _24267_/Q _20443_/X _20504_/X VGND VGND VPWR VPWR _20505_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22238__A2 _22237_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24273_ _24240_/CLK _24273_/D HRESETn VGND VGND VPWR VPWR _20373_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_53_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21485_ _21492_/A VGND VGND VPWR VPWR _21485_/X sky130_fd_sc_hd__buf_2
X_23224_ _23194_/CLK _23224_/D VGND VGND VPWR VPWR _15300_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20436_ _20436_/A VGND VGND VPWR VPWR _20436_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21997__B2 _21993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18862__A1 _17172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23155_ _23347_/CLK _23155_/D VGND VGND VPWR VPWR _12155_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_161_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20367_ _20277_/X _20366_/X _24401_/Q _18894_/B VGND VGND VPWR VPWR _20367_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22106_ _22106_/A VGND VGND VPWR VPWR _22106_/X sky130_fd_sc_hd__buf_2
XFILLER_134_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23086_ _23086_/A _23086_/B _23086_/C _23084_/Y VGND VGND VPWR VPWR HTRANS[1] sky130_fd_sc_hd__or4_4
XANTENNA__11638__B _11637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22512__A _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21749__A1 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20298_ _20298_/A VGND VGND VPWR VPWR _21526_/A sky130_fd_sc_hd__buf_2
XANTENNA__21749__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22037_ _21885_/X _22010_/A _23509_/Q _22000_/A VGND VGND VPWR VPWR _22037_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11654__A _11654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13810_ _12477_/A _24029_/Q VGND VGND VPWR VPWR _13812_/B sky130_fd_sc_hd__or2_4
X_14790_ _14674_/A _14716_/B VGND VGND VPWR VPWR _14790_/X sky130_fd_sc_hd__or2_4
X_23988_ _23668_/CLK _21189_/X VGND VGND VPWR VPWR _21183_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__14030__A _12580_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12111__B1 _11609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13741_ _13753_/A _13741_/B VGND VGND VPWR VPWR _13741_/X sky130_fd_sc_hd__or2_4
X_22939_ _22929_/A _22939_/B _22938_/X VGND VGND VPWR VPWR _22939_/X sky130_fd_sc_hd__and3_4
XFILLER_95_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14965__A _15362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18437__A _18483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21921__B2 _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16460_ _16491_/A _16391_/B VGND VGND VPWR VPWR _16460_/X sky130_fd_sc_hd__or2_4
X_13672_ _13639_/A _13761_/B VGND VGND VPWR VPWR _13673_/C sky130_fd_sc_hd__or2_4
XFILLER_16_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12623_ _12623_/A VGND VGND VPWR VPWR _12973_/A sky130_fd_sc_hd__buf_2
X_15411_ _15411_/A _15411_/B _15410_/X VGND VGND VPWR VPWR _15412_/C sky130_fd_sc_hd__and3_4
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16391_ _16009_/X _16391_/B VGND VGND VPWR VPWR _16391_/X sky130_fd_sc_hd__or2_4
XANTENNA__12485__A _12485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23707__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15342_ _13699_/A _22350_/A VGND VGND VPWR VPWR _15342_/X sky130_fd_sc_hd__or2_4
X_18130_ _18130_/A VGND VGND VPWR VPWR _18130_/Y sky130_fd_sc_hd__inv_2
X_12554_ _12874_/A _12550_/X _12554_/C VGND VGND VPWR VPWR _12554_/X sky130_fd_sc_hd__or3_4
XFILLER_12_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21798__A _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15273_ _13788_/A _15269_/X _15272_/X VGND VGND VPWR VPWR _15273_/X sky130_fd_sc_hd__or3_4
X_18061_ _17583_/B _18059_/B _18060_/X VGND VGND VPWR VPWR _18061_/Y sky130_fd_sc_hd__a21oi_4
X_12485_ _12485_/A VGND VGND VPWR VPWR _13010_/A sky130_fd_sc_hd__buf_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17012_ _23073_/B _17011_/A _16945_/X _17011_/Y VGND VGND VPWR VPWR _17012_/X sky130_fd_sc_hd__o22a_4
X_14224_ _15362_/A VGND VGND VPWR VPWR _14663_/A sky130_fd_sc_hd__buf_2
XFILLER_125_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23857__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14155_ _14155_/A VGND VGND VPWR VPWR _14170_/A sky130_fd_sc_hd__buf_2
XANTENNA__18853__A1 _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13106_ _13090_/A _13104_/X _13105_/X VGND VGND VPWR VPWR _13106_/X sky130_fd_sc_hd__and3_4
XANTENNA__20660__A1 _20635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20660__B2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18963_ _19016_/A VGND VGND VPWR VPWR _18963_/X sky130_fd_sc_hd__buf_2
X_14086_ _14086_/A _14084_/X VGND VGND VPWR VPWR _14086_/X sky130_fd_sc_hd__or2_4
XFILLER_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13037_ _11881_/A _13037_/B _13037_/C VGND VGND VPWR VPWR _13037_/X sky130_fd_sc_hd__and3_4
X_17914_ _17798_/A _17914_/B VGND VGND VPWR VPWR _17916_/C sky130_fd_sc_hd__and2_4
XFILLER_79_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22401__A2 _22397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18894_ _18837_/A _18894_/B VGND VGND VPWR VPWR _18894_/X sky130_fd_sc_hd__or2_4
XFILLER_6_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14859__B _14859_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21038__A _21045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17845_ _17845_/A VGND VGND VPWR VPWR _17845_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17776_ _17675_/X _17706_/Y _17768_/X _17775_/X VGND VGND VPWR VPWR _18013_/C sky130_fd_sc_hd__o22a_4
XFILLER_47_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14988_ _14988_/A _23349_/Q VGND VGND VPWR VPWR _14990_/B sky130_fd_sc_hd__or2_4
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19515_ _19719_/A VGND VGND VPWR VPWR _19515_/X sky130_fd_sc_hd__buf_2
XFILLER_47_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16727_ _16700_/A _16795_/B VGND VGND VPWR VPWR _16727_/X sky130_fd_sc_hd__or2_4
X_13939_ _13710_/A _13848_/B VGND VGND VPWR VPWR _13939_/X sky130_fd_sc_hd__or2_4
XANTENNA__16919__A1 _16918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21912__B2 _21906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17251__A _17251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19446_ _19446_/A VGND VGND VPWR VPWR _19518_/A sky130_fd_sc_hd__buf_2
X_16658_ _16658_/A _24082_/Q VGND VGND VPWR VPWR _16658_/X sky130_fd_sc_hd__or2_4
XANTENNA__17592__A1 _16821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_5_0_HCLK clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15609_ _15625_/A _15603_/X _15608_/X VGND VGND VPWR VPWR _15609_/X sky130_fd_sc_hd__or3_4
X_19377_ _19377_/A VGND VGND VPWR VPWR _19377_/X sky130_fd_sc_hd__buf_2
XANTENNA__12395__A _15894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16589_ _16586_/A _16679_/B VGND VGND VPWR VPWR _16589_/X sky130_fd_sc_hd__or2_4
XFILLER_163_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20479__A1 _18178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18328_ _18215_/X _18326_/X _18240_/X _18327_/X VGND VGND VPWR VPWR _18328_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18259_ _18378_/A _17459_/Y VGND VGND VPWR VPWR _18260_/D sky130_fd_sc_hd__and2_4
XFILLER_163_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21270_ _21268_/X _21269_/X _23945_/Q _21264_/X VGND VGND VPWR VPWR _21270_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21979__A1 _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21979__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11739__A _11739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20221_ _22487_/A _21184_/D VGND VGND VPWR VPWR _20221_/X sky130_fd_sc_hd__or2_4
XANTENNA__19906__A _19402_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18844__A1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20152_ _20200_/A _20152_/B VGND VGND VPWR VPWR _20152_/X sky130_fd_sc_hd__or2_4
XANTENNA__13954__A _13954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20083_ _20082_/X VGND VGND VPWR VPWR _24141_/D sky130_fd_sc_hd__inv_2
XFILLER_170_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23911_ _23111_/CLK _21344_/X VGND VGND VPWR VPWR _13161_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_111_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23842_ _23587_/CLK _23842_/D VGND VGND VPWR VPWR _15494_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24337__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23773_ _23678_/CLK _21583_/X VGND VGND VPWR VPWR _23773_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20985_ _19459_/Y _20873_/A _20598_/B _20697_/A VGND VGND VPWR VPWR _20985_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21903__B2 _21899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17161__A _14084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22724_ _20819_/A _22722_/X _13765_/B _22719_/X VGND VGND VPWR VPWR _22724_/X sky130_fd_sc_hd__o22a_4
XPHY_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16386__A2 _16383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22655_ _22655_/A VGND VGND VPWR VPWR _22655_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21606_ _21706_/A _21656_/B _21706_/C _21184_/D VGND VGND VPWR VPWR _21607_/A sky130_fd_sc_hd__or4_4
X_22586_ _11793_/B VGND VGND VPWR VPWR _22586_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21131__A2 _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24325_ _24292_/CLK _24325_/D HRESETn VGND VGND VPWR VPWR _24325_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21537_ _21524_/X VGND VGND VPWR VPWR _21537_/X sky130_fd_sc_hd__buf_2
X_12270_ _12690_/A _23980_/Q VGND VGND VPWR VPWR _12271_/C sky130_fd_sc_hd__or2_4
X_24256_ _24137_/CLK _24256_/D HRESETn VGND VGND VPWR VPWR _20765_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21468_ _21315_/X _21441_/A _23829_/Q _21431_/A VGND VGND VPWR VPWR _23829_/D sky130_fd_sc_hd__o22a_4
X_23207_ _24039_/CLK _23207_/D VGND VGND VPWR VPWR _13204_/B sky130_fd_sc_hd__dfxtp_4
X_20419_ _20226_/X VGND VGND VPWR VPWR _20895_/A sky130_fd_sc_hd__buf_2
XFILLER_49_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24187_ _24184_/CLK _19882_/X HRESETn VGND VGND VPWR VPWR _17414_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22631__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21399_ _21280_/X _21398_/X _15712_/B _21395_/X VGND VGND VPWR VPWR _21399_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14025__A _13888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23138_ _23303_/CLK _23138_/D VGND VGND VPWR VPWR _15493_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24341__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13864__A _11680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15960_ _15960_/A _23310_/Q VGND VGND VPWR VPWR _15961_/C sky130_fd_sc_hd__or2_4
XFILLER_122_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23069_ _17892_/X _23079_/B VGND VGND VPWR VPWR _23069_/X sky130_fd_sc_hd__or2_4
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16240__A _16239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22395__B2 _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14911_ _11853_/A _11625_/X _14879_/X _11603_/A _14910_/X VGND VGND VPWR VPWR _14911_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_76_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12883__A1 _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15891_ _15903_/A _15829_/B VGND VGND VPWR VPWR _15893_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_60_0_HCLK clkbuf_6_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17630_ _17630_/A _17630_/B VGND VGND VPWR VPWR _17631_/B sky130_fd_sc_hd__nand2_4
X_14842_ _15649_/A _14826_/X _14842_/C VGND VGND VPWR VPWR _14843_/C sky130_fd_sc_hd__or3_4
XFILLER_5_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23073__A _23078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17561_ _16383_/X _17561_/B VGND VGND VPWR VPWR _17562_/A sky130_fd_sc_hd__or2_4
X_14773_ _14773_/A VGND VGND VPWR VPWR _15103_/A sky130_fd_sc_hd__buf_2
X_11985_ _16741_/A _21317_/A VGND VGND VPWR VPWR _11985_/X sky130_fd_sc_hd__or2_4
XANTENNA__14695__A _15620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19300_ _24287_/Q _19236_/B _19299_/Y VGND VGND VPWR VPWR _24287_/D sky130_fd_sc_hd__o21a_4
X_16512_ _16479_/X _16435_/B VGND VGND VPWR VPWR _16512_/X sky130_fd_sc_hd__or2_4
XANTENNA__17071__A _17070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13724_ _13697_/A VGND VGND VPWR VPWR _13743_/A sky130_fd_sc_hd__buf_2
X_17492_ _16678_/A _17378_/X _17379_/X VGND VGND VPWR VPWR _17492_/X sky130_fd_sc_hd__o21a_4
XFILLER_95_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19231_ _19231_/A _19230_/X VGND VGND VPWR VPWR _19231_/X sky130_fd_sc_hd__and2_4
X_16443_ _16413_/A _16443_/B VGND VGND VPWR VPWR _16443_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13655_ _13655_/A VGND VGND VPWR VPWR _13656_/A sky130_fd_sc_hd__buf_2
XFILLER_20_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12606_ _13052_/A VGND VGND VPWR VPWR _12623_/A sky130_fd_sc_hd__buf_2
X_19162_ _19160_/X VGND VGND VPWR VPWR _19162_/Y sky130_fd_sc_hd__inv_2
X_16374_ _11715_/A _16296_/B VGND VGND VPWR VPWR _16374_/X sky130_fd_sc_hd__or2_4
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13586_ _13586_/A VGND VGND VPWR VPWR _14480_/A sky130_fd_sc_hd__buf_2
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18523__B1 _17890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18113_ _18310_/A _18113_/B VGND VGND VPWR VPWR _18113_/X sky130_fd_sc_hd__or2_4
X_12537_ _12537_/A VGND VGND VPWR VPWR _12905_/A sky130_fd_sc_hd__buf_2
X_15325_ _15325_/A VGND VGND VPWR VPWR _15326_/A sky130_fd_sc_hd__buf_2
XANTENNA__20330__B1 _20638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19093_ _11522_/A _11521_/X _19088_/Y VGND VGND VPWR VPWR _19093_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12943__A _12943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18044_ _17850_/X _17149_/X _17812_/X _17168_/X VGND VGND VPWR VPWR _18044_/Y sky130_fd_sc_hd__a22oi_4
X_15256_ _14140_/A _23352_/Q VGND VGND VPWR VPWR _15256_/X sky130_fd_sc_hd__or2_4
X_12468_ _12468_/A VGND VGND VPWR VPWR _12469_/A sky130_fd_sc_hd__buf_2
XANTENNA__12662__B _12565_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14207_ _11654_/A VGND VGND VPWR VPWR _14635_/A sky130_fd_sc_hd__buf_2
X_15187_ _15076_/A _15123_/B VGND VGND VPWR VPWR _15188_/C sky130_fd_sc_hd__or2_4
XANTENNA__18826__A1 _14548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12399_ _12363_/X _12399_/B VGND VGND VPWR VPWR _12400_/C sky130_fd_sc_hd__or2_4
XFILLER_126_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14138_ _14138_/A _23967_/Q VGND VGND VPWR VPWR _14139_/C sky130_fd_sc_hd__or2_4
X_19995_ _17961_/X _19983_/X _19993_/Y _19994_/X VGND VGND VPWR VPWR _19995_/X sky130_fd_sc_hd__o22a_4
XFILLER_154_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18946_ _11543_/B VGND VGND VPWR VPWR _18948_/B sky130_fd_sc_hd__inv_2
X_14069_ _11698_/A _14069_/B _14068_/X VGND VGND VPWR VPWR _14069_/X sky130_fd_sc_hd__and3_4
XANTENNA__22386__B2 _22380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21991__A _21991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24185__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24126__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18877_ _18838_/X VGND VGND VPWR VPWR _18877_/X sky130_fd_sc_hd__buf_2
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17828_ _17825_/X _17826_/X _17230_/X _17827_/X VGND VGND VPWR VPWR _17828_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22138__B2 _22130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17759_ _17737_/X _17739_/X _17758_/X VGND VGND VPWR VPWR _17760_/C sky130_fd_sc_hd__or3_4
XFILLER_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18077__A _18335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20770_ _20770_/A VGND VGND VPWR VPWR _20770_/X sky130_fd_sc_hd__buf_2
XFILLER_23_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21361__A2 _21355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19429_ _19425_/X _18662_/X _19428_/X _24218_/Q VGND VGND VPWR VPWR _24218_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13014__A _12492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22440_ _22440_/A VGND VGND VPWR VPWR _22440_/X sky130_fd_sc_hd__buf_2
XANTENNA__21113__A2 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22310__B2 _22305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22371_ _22113_/X _22369_/X _23309_/Q _22366_/X VGND VGND VPWR VPWR _23309_/D sky130_fd_sc_hd__o22a_4
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12853__A _12884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24110_ _24078_/CLK _24110_/D VGND VGND VPWR VPWR _24110_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_148_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_HCLK clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_2_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21322_ _21322_/A VGND VGND VPWR VPWR _21338_/A sky130_fd_sc_hd__inv_2
XFILLER_85_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24041_ _23337_/CLK _24041_/D VGND VGND VPWR VPWR _24041_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_151_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21253_ _21251_/X _21245_/X _16412_/B _21252_/X VGND VGND VPWR VPWR _23952_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19636__A HRDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14551__A1 _14483_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22613__A2 _22608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20204_ _19402_/A _17005_/X _20200_/A _20203_/X VGND VGND VPWR VPWR _20205_/A sky130_fd_sc_hd__o22a_4
XANTENNA__16828__B1 _16905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21184_ _21184_/A _21134_/B _21184_/C _21184_/D VGND VGND VPWR VPWR _21184_/X sky130_fd_sc_hd__or4_4
XFILLER_145_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13684__A _12299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14303__A1 _13689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17156__A _17156_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20135_ _11569_/B VGND VGND VPWR VPWR _20135_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16060__A _11759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22377__B2 _22373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20066_ _19950_/X VGND VGND VPWR VPWR _20066_/X sky130_fd_sc_hd__buf_2
XFILLER_86_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_4_0_HCLK_A clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23825_ _23889_/CLK _23825_/D VGND VGND VPWR VPWR _23825_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__A _11932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23756_ _24045_/CLK _23756_/D VGND VGND VPWR VPWR _23756_/Q sky130_fd_sc_hd__dfxtp_4
X_11770_ _11832_/A _21080_/A VGND VGND VPWR VPWR _11770_/X sky130_fd_sc_hd__or2_4
X_20968_ _24407_/Q _20427_/A _24439_/Q _20282_/A VGND VGND VPWR VPWR _20968_/X sky130_fd_sc_hd__o22a_4
XPHY_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _20531_/A _22701_/X _12824_/B _22705_/X VGND VGND VPWR VPWR _23114_/D sky130_fd_sc_hd__o22a_4
XPHY_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23687_ _23750_/CLK _23687_/D VGND VGND VPWR VPWR _23687_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20899_ _20943_/A _20898_/X VGND VGND VPWR VPWR _20899_/X sky130_fd_sc_hd__and2_4
XPHY_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13440_ _12871_/A VGND VGND VPWR VPWR _13441_/A sky130_fd_sc_hd__buf_2
XFILLER_55_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22638_ _22637_/X VGND VGND VPWR VPWR _22672_/A sky130_fd_sc_hd__buf_2
XANTENNA__22237__A _22244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21141__A _21155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13371_ _13379_/A _23462_/Q VGND VGND VPWR VPWR _13372_/C sky130_fd_sc_hd__or2_4
XFILLER_167_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13859__A _12251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22569_ _22555_/A VGND VGND VPWR VPWR _22569_/X sky130_fd_sc_hd__buf_2
X_12322_ _12322_/A VGND VGND VPWR VPWR _13052_/A sky130_fd_sc_hd__buf_2
X_15110_ _15103_/A _15033_/B VGND VGND VPWR VPWR _15110_/X sky130_fd_sc_hd__or2_4
X_16090_ _15967_/A _16090_/B VGND VGND VPWR VPWR _16092_/B sky130_fd_sc_hd__or2_4
XFILLER_6_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24308_ _24368_/CLK _19259_/X HRESETn VGND VGND VPWR VPWR _24308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20980__A _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15041_ _13606_/A _15104_/B VGND VGND VPWR VPWR _15041_/X sky130_fd_sc_hd__or2_4
X_12253_ _12228_/A _12357_/B VGND VGND VPWR VPWR _12253_/X sky130_fd_sc_hd__or2_4
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24239_ _24158_/CLK _19394_/X HRESETn VGND VGND VPWR VPWR _24239_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18808__A1 _13262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22604__A2 _22601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20615__A1 _20533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20615__B2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23068__A _23078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12184_ _12112_/Y _12180_/X _12183_/X VGND VGND VPWR VPWR _16905_/B sky130_fd_sc_hd__o21ai_4
XFILLER_150_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18800_ _16240_/X _18796_/X _11575_/A _18797_/X VGND VGND VPWR VPWR _18800_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19780_ _19776_/X _19779_/X _19537_/B _19705_/X VGND VGND VPWR VPWR _19780_/X sky130_fd_sc_hd__o22a_4
X_16992_ _17675_/A _16992_/B VGND VGND VPWR VPWR _18107_/A sky130_fd_sc_hd__or2_4
XFILLER_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22368__B2 _22366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18731_ _18731_/A _18729_/X VGND VGND VPWR VPWR _18731_/X sky130_fd_sc_hd__or2_4
X_15943_ _16011_/A VGND VGND VPWR VPWR _15993_/A sky130_fd_sc_hd__buf_2
XANTENNA__24259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21040__B2 _21035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18662_ _22931_/B _18661_/X _22931_/B _18661_/X VGND VGND VPWR VPWR _18662_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15874_ _13521_/X _15872_/X _15873_/X VGND VGND VPWR VPWR _15874_/X sky130_fd_sc_hd__and3_4
XANTENNA__12003__A _11905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17613_ _18587_/B _17612_/Y _17412_/B VGND VGND VPWR VPWR _17613_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14825_ _15106_/A _14821_/X _14825_/C VGND VGND VPWR VPWR _14825_/X sky130_fd_sc_hd__or3_4
X_18593_ _18499_/X _18591_/X _18527_/X _18592_/X VGND VGND VPWR VPWR _18593_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17513__B _17515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12938__A _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11842__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15314__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17544_ _17544_/A VGND VGND VPWR VPWR _17544_/Y sky130_fd_sc_hd__inv_2
X_14756_ _12288_/A _14756_/B _14755_/X VGND VGND VPWR VPWR _14756_/X sky130_fd_sc_hd__or3_4
X_11968_ _15420_/A VGND VGND VPWR VPWR _11969_/A sky130_fd_sc_hd__buf_2
XANTENNA__12657__B _12657_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21343__A2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13707_ _13751_/A _13707_/B VGND VGND VPWR VPWR _13708_/C sky130_fd_sc_hd__or2_4
XANTENNA__15033__B _15033_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17475_ _17145_/Y _17475_/B VGND VGND VPWR VPWR _17640_/A sky130_fd_sc_hd__or2_4
X_11899_ _14421_/A VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_67_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR _23862_/CLK sky130_fd_sc_hd__clkbuf_1
X_14687_ _15606_/A VGND VGND VPWR VPWR _15620_/A sky130_fd_sc_hd__buf_2
X_19214_ _19135_/A _19215_/A _19213_/Y VGND VGND VPWR VPWR _19214_/X sky130_fd_sc_hd__o21a_4
X_16426_ _15998_/X _16424_/X _16425_/X VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__and3_4
X_13638_ _15447_/A VGND VGND VPWR VPWR _13639_/A sky130_fd_sc_hd__buf_2
XFILLER_20_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22147__A _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13769__A _12610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19145_ _24324_/Q _19144_/X VGND VGND VPWR VPWR _19145_/X sky130_fd_sc_hd__and2_4
X_16357_ _16333_/A _16289_/B VGND VGND VPWR VPWR _16359_/B sky130_fd_sc_hd__or2_4
XFILLER_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16145__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12673__A _12975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13569_ _13485_/X _13583_/A VGND VGND VPWR VPWR _13570_/A sky130_fd_sc_hd__or2_4
XFILLER_34_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15308_ _15017_/A _23864_/Q VGND VGND VPWR VPWR _15308_/X sky130_fd_sc_hd__or2_4
X_19076_ _19076_/A VGND VGND VPWR VPWR _19076_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16288_ _15936_/X _16286_/X _16287_/X VGND VGND VPWR VPWR _16292_/B sky130_fd_sc_hd__and3_4
X_18027_ _18026_/X VGND VGND VPWR VPWR _18027_/X sky130_fd_sc_hd__buf_2
X_15239_ _12336_/A _15239_/B _15239_/C VGND VGND VPWR VPWR _15240_/C sky130_fd_sc_hd__and3_4
XFILLER_126_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19978_ _24500_/Q VGND VGND VPWR VPWR _19978_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18929_ _17161_/X _18927_/X _24384_/Q _18928_/X VGND VGND VPWR VPWR _18929_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_0_HCLK HCLK VGND VGND VPWR VPWR clkbuf_0_HCLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13009__A _12537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21940_ _21939_/X VGND VGND VPWR VPWR _21941_/A sky130_fd_sc_hd__buf_2
XANTENNA__17786__A1 _16935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21226__A _21219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21871_ _21869_/X _21863_/X _14380_/B _21870_/X VGND VGND VPWR VPWR _21871_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12848__A _12848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11752__A _11752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23610_ _24090_/CLK _23610_/D VGND VGND VPWR VPWR _23610_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20822_ _21007_/B _20671_/A VGND VGND VPWR VPWR _20822_/X sky130_fd_sc_hd__or2_4
XANTENNA__15224__A _14201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18735__B1 _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22531__B2 _22526_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23541_ _23617_/CLK _23541_/D VGND VGND VPWR VPWR _23541_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20753_ _20261_/X VGND VGND VPWR VPWR _20753_/X sky130_fd_sc_hd__buf_2
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24200__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23472_ _23728_/CLK _22107_/X VGND VGND VPWR VPWR _16476_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20684_ _20539_/X _20683_/X _19144_/A _20549_/X VGND VGND VPWR VPWR _20685_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22057__A _22057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22423_ _20415_/A VGND VGND VPWR VPWR _22423_/X sky130_fd_sc_hd__buf_2
XANTENNA__21098__B2 _21094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13679__A _13676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12583__A _12583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22354_ _11774_/B VGND VGND VPWR VPWR _22354_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21305_ _21238_/A VGND VGND VPWR VPWR _21305_/X sky130_fd_sc_hd__buf_2
XANTENNA__15894__A _15894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22285_ _22105_/X _22280_/X _16390_/B _22284_/X VGND VGND VPWR VPWR _22285_/X sky130_fd_sc_hd__o22a_4
XFILLER_163_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24024_ _23290_/CLK _24024_/D VGND VGND VPWR VPWR _24024_/Q sky130_fd_sc_hd__dfxtp_4
X_21236_ _21134_/A _21134_/B _21184_/C _21236_/D VGND VGND VPWR VPWR _21236_/X sky130_fd_sc_hd__or4_4
XANTENNA__11927__A _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21270__B2 _21264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21167_ _20745_/X _21162_/X _24001_/Q _21166_/X VGND VGND VPWR VPWR _24001_/D sky130_fd_sc_hd__o22a_4
XFILLER_160_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20118_ NMI VGND VGND VPWR VPWR _20118_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21098_ _20441_/X _21097_/X _24046_/Q _21094_/X VGND VGND VPWR VPWR _21098_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12940_ _12940_/A _24009_/Q VGND VGND VPWR VPWR _12941_/C sky130_fd_sc_hd__or2_4
X_20049_ _20040_/X _16986_/A _20046_/X _20048_/X VGND VGND VPWR VPWR _20050_/A sky130_fd_sc_hd__o22a_4
XFILLER_74_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21136__A _21136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12871_ _12871_/A _23337_/Q VGND VGND VPWR VPWR _12871_/X sky130_fd_sc_hd__or2_4
XANTENNA__20040__A _18670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12758__A _12758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14610_ _13589_/A _14606_/X _14610_/C VGND VGND VPWR VPWR _14610_/X sky130_fd_sc_hd__or3_4
X_11822_ _11834_/A _11822_/B _11821_/X VGND VGND VPWR VPWR _11822_/X sky130_fd_sc_hd__and3_4
X_23808_ _23649_/CLK _21505_/X VGND VGND VPWR VPWR _14068_/B sky130_fd_sc_hd__dfxtp_4
X_15590_ _12337_/A _15587_/X _15590_/C VGND VGND VPWR VPWR _15591_/C sky130_fd_sc_hd__and3_4
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14541_/A _14469_/B VGND VGND VPWR VPWR _14541_/X sky130_fd_sc_hd__or2_4
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11753_ _11753_/A VGND VGND VPWR VPWR _12596_/A sky130_fd_sc_hd__buf_2
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23739_ _23675_/CLK _23739_/D VGND VGND VPWR VPWR _14488_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17260_/A VGND VGND VPWR VPWR _17260_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11684_ _13415_/A VGND VGND VPWR VPWR _11684_/X sky130_fd_sc_hd__buf_2
X_14472_ _12266_/A _14472_/B _14471_/X VGND VGND VPWR VPWR _14472_/X sky130_fd_sc_hd__or3_4
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _16181_/X _23629_/Q VGND VGND VPWR VPWR _16211_/X sky130_fd_sc_hd__or2_4
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _13427_/A _23749_/Q VGND VGND VPWR VPWR _13424_/C sky130_fd_sc_hd__or2_4
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13589__A _13589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17191_ _17140_/Y _17144_/A _14549_/Y _17146_/A VGND VGND VPWR VPWR _17191_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12493__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16142_ _16142_/A _16142_/B VGND VGND VPWR VPWR _16142_/X sky130_fd_sc_hd__or2_4
X_13354_ _13410_/A _13354_/B _13354_/C VGND VGND VPWR VPWR _13355_/C sky130_fd_sc_hd__and3_4
XFILLER_155_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12305_ _12747_/A VGND VGND VPWR VPWR _13333_/A sky130_fd_sc_hd__buf_2
XFILLER_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13285_ _13321_/A _13285_/B _13284_/X VGND VGND VPWR VPWR _13285_/X sky130_fd_sc_hd__and3_4
X_16073_ _16049_/A _16010_/B VGND VGND VPWR VPWR _16074_/C sky130_fd_sc_hd__or2_4
XFILLER_6_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18180__A _17768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12236_ _12236_/A VGND VGND VPWR VPWR _12748_/A sky130_fd_sc_hd__buf_2
X_19901_ _19900_/X VGND VGND VPWR VPWR _19901_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_9_0_HCLK clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15024_ _13953_/A _23829_/Q VGND VGND VPWR VPWR _15025_/C sky130_fd_sc_hd__or2_4
XFILLER_155_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11837__A _16647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19832_ _19647_/Y _19823_/X _19831_/Y VGND VGND VPWR VPWR _19832_/X sky130_fd_sc_hd__o21a_4
X_12167_ _12167_/A _23891_/Q VGND VGND VPWR VPWR _12168_/C sky130_fd_sc_hd__or2_4
XANTENNA__15309__A _15018_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14213__A _13882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19763_ _19752_/B VGND VGND VPWR VPWR _19763_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11556__B IRQ[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16975_ _17740_/A _16973_/X _17734_/A VGND VGND VPWR VPWR _16975_/X sky130_fd_sc_hd__or3_4
XFILLER_1_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12098_ _12097_/X _12173_/B VGND VGND VPWR VPWR _12098_/X sky130_fd_sc_hd__or2_4
XANTENNA__22430__A _20485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18714_ _18565_/A _18714_/B VGND VGND VPWR VPWR _18714_/X sky130_fd_sc_hd__and2_4
XANTENNA__17524__A _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15926_ _15920_/X _16842_/B _15925_/Y VGND VGND VPWR VPWR _15926_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__22210__B1 _13761_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19694_ _19849_/A _19839_/A _19879_/D _19687_/C VGND VGND VPWR VPWR _19694_/X sky130_fd_sc_hd__and4_4
XANTENNA__21564__A2 _21554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_30_0_HCLK clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18645_ _17652_/X _18626_/X _16935_/A _18644_/X VGND VGND VPWR VPWR _18645_/X sky130_fd_sc_hd__o22a_4
X_15857_ _12373_/X _15796_/B VGND VGND VPWR VPWR _15857_/X sky130_fd_sc_hd__or2_4
XFILLER_65_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12668__A _12942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15044__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24223__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14808_ _14680_/A _14806_/X _14808_/C VGND VGND VPWR VPWR _14809_/C sky130_fd_sc_hd__and3_4
X_18576_ _24212_/Q _18576_/B VGND VGND VPWR VPWR _18698_/B sky130_fd_sc_hd__or2_4
XFILLER_80_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15788_ _15788_/A _15787_/X VGND VGND VPWR VPWR _16855_/A sky130_fd_sc_hd__or2_4
XFILLER_33_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18717__B1 _18712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21316__A2 _21269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22513__B2 _22512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17527_ _17499_/Y _17509_/Y _17517_/Y _17527_/D VGND VGND VPWR VPWR _17527_/X sky130_fd_sc_hd__or4_4
XFILLER_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15979__A _11971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14739_ _13652_/A _14739_/B VGND VGND VPWR VPWR _14741_/B sky130_fd_sc_hd__or2_4
XFILLER_71_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17458_ _12982_/X _17460_/B VGND VGND VPWR VPWR _17459_/A sky130_fd_sc_hd__or2_4
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13499__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16409_ _16409_/A _16409_/B VGND VGND VPWR VPWR _16409_/X sky130_fd_sc_hd__or2_4
XFILLER_119_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17389_ _17360_/A _17389_/B VGND VGND VPWR VPWR _17389_/X sky130_fd_sc_hd__or2_4
X_19128_ _18948_/D _19126_/Y _19124_/X _19127_/Y VGND VGND VPWR VPWR _19129_/A sky130_fd_sc_hd__o22a_4
XFILLER_134_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19059_ _11528_/A _11528_/B _19054_/Y VGND VGND VPWR VPWR _19059_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_173_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22070_ _21855_/X _22067_/X _15508_/B _22064_/X VGND VGND VPWR VPWR _23490_/D sky130_fd_sc_hd__o22a_4
XFILLER_114_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21021_ _20977_/A _21020_/X VGND VGND VPWR VPWR _21021_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15219__A _14225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14123__A _13788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17208__B1 _17162_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22972_ _22910_/X VGND VGND VPWR VPWR _22973_/B sky130_fd_sc_hd__buf_2
XFILLER_110_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21555__A2 _21554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21923_ _21923_/A VGND VGND VPWR VPWR _21923_/X sky130_fd_sc_hd__buf_2
XFILLER_28_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21854_ _21853_/X _21851_/X _15822_/B _21846_/X VGND VGND VPWR VPWR _21854_/X sky130_fd_sc_hd__o22a_4
XFILLER_167_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12297__B _24108_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18708__B1 _17919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22504__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20805_ _20845_/A _20803_/X _20804_/X VGND VGND VPWR VPWR _20805_/X sky130_fd_sc_hd__and3_4
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21785_ _21565_/X _21784_/X _15705_/B _21781_/X VGND VGND VPWR VPWR _23652_/D sky130_fd_sc_hd__o22a_4
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18265__A _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14793__A _15091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23524_ _23588_/CLK _22018_/X VGND VGND VPWR VPWR _15658_/B sky130_fd_sc_hd__dfxtp_4
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20736_ _20539_/X _20735_/X _24321_/Q _20549_/X VGND VGND VPWR VPWR _20736_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_50_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR _23728_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17931__A1 _17811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23455_ _23101_/CLK _23455_/D VGND VGND VPWR VPWR _23455_/Q sky130_fd_sc_hd__dfxtp_4
X_20667_ _20670_/A VGND VGND VPWR VPWR _20668_/A sky130_fd_sc_hd__inv_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22406_ _22405_/X VGND VGND VPWR VPWR _22462_/A sky130_fd_sc_hd__buf_2
XFILLER_104_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23386_ _23772_/CLK _22266_/X VGND VGND VPWR VPWR _23386_/Q sky130_fd_sc_hd__dfxtp_4
X_20598_ _20307_/X _20598_/B VGND VGND VPWR VPWR _20598_/X sky130_fd_sc_hd__and2_4
XFILLER_164_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22515__A _22508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22337_ _22337_/A VGND VGND VPWR VPWR _23333_/D sky130_fd_sc_hd__buf_2
XFILLER_139_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21491__B2 _21489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13070_ _13085_/A _12999_/B VGND VGND VPWR VPWR _13070_/X sky130_fd_sc_hd__or2_4
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22268_ _22163_/X _22265_/X _23384_/Q _22262_/X VGND VGND VPWR VPWR _23384_/D sky130_fd_sc_hd__o22a_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24007_ _24039_/CLK _21158_/X VGND VGND VPWR VPWR _24007_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_133_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12021_ _12020_/X VGND VGND VPWR VPWR _12021_/Y sky130_fd_sc_hd__inv_2
X_21219_ _21219_/A VGND VGND VPWR VPWR _21219_/X sky130_fd_sc_hd__buf_2
XFILLER_120_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22199_ _22129_/X _22194_/X _23430_/Q _22198_/X VGND VGND VPWR VPWR _23430_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14033__A _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21794__A2 _21791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13872__A _13719_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16760_ _16606_/A _16760_/B _16759_/X VGND VGND VPWR VPWR _16760_/X sky130_fd_sc_hd__or3_4
XANTENNA__24246__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13484__A1 _11971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13972_ _12250_/A _13970_/X _13972_/C VGND VGND VPWR VPWR _13973_/C sky130_fd_sc_hd__and3_4
XFILLER_93_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15711_ _11887_/A _23716_/Q VGND VGND VPWR VPWR _15713_/B sky130_fd_sc_hd__or2_4
X_12923_ _12923_/A _23785_/Q VGND VGND VPWR VPWR _12923_/X sky130_fd_sc_hd__or2_4
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16691_ _16691_/A _23537_/Q VGND VGND VPWR VPWR _16692_/C sky130_fd_sc_hd__or2_4
XANTENNA__12488__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18430_ _18356_/X _18427_/X _18396_/X _18429_/X VGND VGND VPWR VPWR _18430_/X sky130_fd_sc_hd__o22a_4
X_15642_ _15642_/A _24097_/Q VGND VGND VPWR VPWR _15643_/C sky130_fd_sc_hd__or2_4
X_12854_ _12854_/A VGND VGND VPWR VPWR _12860_/A sky130_fd_sc_hd__buf_2
XFILLER_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15799__A _12847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11805_ _11836_/A _21937_/A VGND VGND VPWR VPWR _11805_/X sky130_fd_sc_hd__or2_4
X_18361_ _16964_/Y VGND VGND VPWR VPWR _18500_/A sky130_fd_sc_hd__buf_2
X_15573_ _12434_/A _15634_/B VGND VGND VPWR VPWR _15573_/X sky130_fd_sc_hd__or2_4
X_12785_ _12801_/A _12785_/B VGND VGND VPWR VPWR _12786_/C sky130_fd_sc_hd__or2_4
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17312_ _18603_/B _17305_/X _17311_/Y VGND VGND VPWR VPWR _17312_/Y sky130_fd_sc_hd__a21oi_4
X_14524_ _14517_/A _14460_/B VGND VGND VPWR VPWR _14525_/C sky130_fd_sc_hd__or2_4
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _11736_/A VGND VGND VPWR VPWR _12634_/A sky130_fd_sc_hd__buf_2
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18292_ _17605_/D _18291_/X VGND VGND VPWR VPWR _18292_/X sky130_fd_sc_hd__or2_4
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _17227_/X _17241_/X _17880_/A VGND VGND VPWR VPWR _17243_/X sky130_fd_sc_hd__o21a_4
XFILLER_159_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14455_ _12531_/A _14455_/B VGND VGND VPWR VPWR _14455_/X sky130_fd_sc_hd__or2_4
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11667_ _11666_/X VGND VGND VPWR VPWR _11668_/A sky130_fd_sc_hd__buf_2
XANTENNA__14208__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _13398_/A _13406_/B _13406_/C VGND VGND VPWR VPWR _13407_/C sky130_fd_sc_hd__and3_4
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17174_ _15913_/Y _17107_/X _17173_/Y _17074_/X VGND VGND VPWR VPWR _17174_/X sky130_fd_sc_hd__o22a_4
X_14386_ _14386_/A VGND VGND VPWR VPWR _14506_/A sky130_fd_sc_hd__buf_2
X_11598_ _11592_/X _11647_/B _17017_/A _11598_/D VGND VGND VPWR VPWR _11598_/X sky130_fd_sc_hd__or4_4
XANTENNA__22425__A _22110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16125_ _16156_/A _16193_/B VGND VGND VPWR VPWR _16125_/X sky130_fd_sc_hd__or2_4
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13337_ _13324_/A _13335_/X _13336_/X VGND VGND VPWR VPWR _13338_/C sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_4_7_0_HCLK_A clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16056_ _16056_/A _16054_/X _16056_/C VGND VGND VPWR VPWR _16056_/X sky130_fd_sc_hd__and3_4
XANTENNA__13766__B _13766_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13268_ _13126_/X VGND VGND VPWR VPWR _13269_/B sky130_fd_sc_hd__inv_2
XFILLER_97_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20037__A2 _20031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15007_ _15007_/A _23925_/Q VGND VGND VPWR VPWR _15009_/B sky130_fd_sc_hd__or2_4
XANTENNA__24203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15039__A _12467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12219_ _13637_/A VGND VGND VPWR VPWR _12294_/A sky130_fd_sc_hd__buf_2
X_13199_ _13220_/A _13199_/B VGND VGND VPWR VPWR _13199_/X sky130_fd_sc_hd__or2_4
XFILLER_124_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21785__A2 _21784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19815_ _19889_/A _19815_/B VGND VGND VPWR VPWR _19815_/X sky130_fd_sc_hd__or2_4
XANTENNA__22798__C _20218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14878__A _13981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13782__A _13692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19746_ _19743_/Y _19745_/X _19819_/A VGND VGND VPWR VPWR _19746_/X sky130_fd_sc_hd__o21a_4
X_16958_ _16958_/A VGND VGND VPWR VPWR _16986_/A sky130_fd_sc_hd__inv_2
XFILLER_110_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22734__A1 _21313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22734__B2 _22698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15909_ _13520_/A _15909_/B _15909_/C VGND VGND VPWR VPWR _15910_/C sky130_fd_sc_hd__or3_4
X_19677_ _19677_/A VGND VGND VPWR VPWR _19894_/C sky130_fd_sc_hd__buf_2
XFILLER_53_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16889_ _15933_/X _16246_/B _16243_/X VGND VGND VPWR VPWR _16889_/X sky130_fd_sc_hd__o21a_4
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18628_ _17748_/A VGND VGND VPWR VPWR _18628_/X sky130_fd_sc_hd__buf_2
XFILLER_64_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18559_ _18413_/X _17401_/X _18557_/Y _18467_/X _18558_/Y VGND VGND VPWR VPWR _18560_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_36_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21570_ _21570_/A VGND VGND VPWR VPWR _21570_/X sky130_fd_sc_hd__buf_2
XFILLER_36_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21170__B1 _23999_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_37_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_74_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20521_ _20516_/X _20520_/X _11536_/A _20475_/X VGND VGND VPWR VPWR _20521_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19909__A _22846_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14118__A _12194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13022__A _12506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23240_ _23656_/CLK _23240_/D VGND VGND VPWR VPWR _13035_/B sky130_fd_sc_hd__dfxtp_4
X_20452_ _20452_/A VGND VGND VPWR VPWR _20452_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22335__A _13148_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24119__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23171_ _23203_/CLK _22617_/X VGND VGND VPWR VPWR _15868_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17429__A _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12861__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20383_ _24432_/Q _18837_/B _24464_/Q _20282_/X VGND VGND VPWR VPWR _20383_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13950__A2 _13947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22122_ _20558_/A VGND VGND VPWR VPWR _22122_/X sky130_fd_sc_hd__buf_2
XFILLER_133_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13676__B _24094_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22053_ _22060_/A VGND VGND VPWR VPWR _22053_/X sky130_fd_sc_hd__buf_2
XANTENNA__21225__B2 _21223_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19644__A _19811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24269__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21776__A2 _21770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21004_ _21313_/A VGND VGND VPWR VPWR _21004_/X sky130_fd_sc_hd__buf_2
XFILLER_173_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20984__B1 HRDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22725__A1 _20841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22725__B2 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22955_ _18568_/X _22938_/B VGND VGND VPWR VPWR _22955_/X sky130_fd_sc_hd__or2_4
XFILLER_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21906_ _21906_/A VGND VGND VPWR VPWR _21906_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_119_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR _23323_/CLK sky130_fd_sc_hd__clkbuf_1
X_22886_ _22876_/X _22826_/X _17425_/Y _22877_/X VGND VGND VPWR VPWR _22886_/X sky130_fd_sc_hd__o22a_4
X_21837_ _21836_/X _21827_/X _12723_/B _21834_/X VGND VGND VPWR VPWR _21837_/X sky130_fd_sc_hd__o22a_4
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11940__A _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12570_ _12570_/A _12568_/X _12569_/X VGND VGND VPWR VPWR _12570_/X sky130_fd_sc_hd__and3_4
X_21768_ _21536_/X _21763_/X _16439_/B _21767_/X VGND VGND VPWR VPWR _23664_/D sky130_fd_sc_hd__o22a_4
XFILLER_106_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20719_ _21570_/A VGND VGND VPWR VPWR _20719_/X sky130_fd_sc_hd__buf_2
X_23507_ _23764_/CLK _23507_/D VGND VGND VPWR VPWR _23507_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _11521_/A _19099_/A VGND VGND VPWR VPWR _11521_/X sky130_fd_sc_hd__or2_4
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24487_ _24495_/CLK _24487_/D HRESETn VGND VGND VPWR VPWR _24487_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21699_ _21589_/X _21698_/X _14686_/B _21695_/X VGND VGND VPWR VPWR _23706_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14028__A _11659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14240_ _14240_/A _23423_/Q VGND VGND VPWR VPWR _14240_/X sky130_fd_sc_hd__or2_4
XFILLER_172_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23438_ _23438_/CLK _22188_/X VGND VGND VPWR VPWR _23438_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14171_ _14171_/A _14171_/B _14171_/C VGND VGND VPWR VPWR _14172_/C sky130_fd_sc_hd__and3_4
XANTENNA__13867__A _13884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23369_ _23561_/CLK _22295_/X VGND VGND VPWR VPWR _23369_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_152_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17339__A _17339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21464__B2 _21459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12771__A _13556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16243__A _16162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13122_ _13100_/A _13122_/B _13122_/C VGND VGND VPWR VPWR _13122_/X sky130_fd_sc_hd__or3_4
XFILLER_125_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13053_ _13053_/A VGND VGND VPWR VPWR _13094_/A sky130_fd_sc_hd__buf_2
X_17930_ _17930_/A VGND VGND VPWR VPWR _17930_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12004_ _12015_/A VGND VGND VPWR VPWR _12106_/A sky130_fd_sc_hd__buf_2
X_17861_ _17233_/X _17215_/X _17231_/X _17191_/X VGND VGND VPWR VPWR _17861_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14698__A _13894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16812_ _16759_/A _16810_/X _16811_/X VGND VGND VPWR VPWR _16812_/X sky130_fd_sc_hd__and3_4
X_19600_ _19744_/A _19558_/A _19558_/X VGND VGND VPWR VPWR _19600_/X sky130_fd_sc_hd__o21a_4
XFILLER_120_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17792_ _17094_/Y VGND VGND VPWR VPWR _17792_/X sky130_fd_sc_hd__buf_2
XFILLER_59_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21519__A2 _21492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22716__B2 _22712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19531_ _19445_/A _19530_/X HRDATA[8] _19461_/A VGND VGND VPWR VPWR _19532_/A sky130_fd_sc_hd__o22a_4
X_16743_ _11943_/X _16743_/B _16743_/C VGND VGND VPWR VPWR _16747_/B sky130_fd_sc_hd__and3_4
X_13955_ _13955_/A VGND VGND VPWR VPWR _13985_/A sky130_fd_sc_hd__buf_2
XFILLER_98_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22192__A2 _22187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12906_ _12906_/A _12964_/B VGND VGND VPWR VPWR _12907_/C sky130_fd_sc_hd__or2_4
XANTENNA__13107__A _13091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19462_ _19518_/A _19458_/Y _19459_/Y _19461_/X VGND VGND VPWR VPWR _19506_/A sky130_fd_sc_hd__o22a_4
XANTENNA__17802__A _17801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12011__A _11960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16674_ _16678_/A _16674_/B _16674_/C VGND VGND VPWR VPWR _16675_/C sky130_fd_sc_hd__and3_4
XFILLER_59_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13886_ _13886_/A _13886_/B _13886_/C VGND VGND VPWR VPWR _13893_/B sky130_fd_sc_hd__and3_4
X_18413_ _18413_/A VGND VGND VPWR VPWR _18413_/X sky130_fd_sc_hd__buf_2
XFILLER_59_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21324__A _21331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15625_ _15625_/A _15625_/B _15625_/C VGND VGND VPWR VPWR _15633_/B sky130_fd_sc_hd__or3_4
X_12837_ _13370_/A _23658_/Q VGND VGND VPWR VPWR _12838_/C sky130_fd_sc_hd__or2_4
X_19393_ _19389_/X _17966_/X _19392_/X _24240_/Q VGND VGND VPWR VPWR _19393_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12946__A _12962_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16418__A _13475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11850__A _16684_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15322__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18344_ _17920_/X _18443_/B _18089_/X _18343_/X VGND VGND VPWR VPWR _18344_/X sky130_fd_sc_hd__a211o_4
X_15556_ _11900_/A _24065_/Q VGND VGND VPWR VPWR _15557_/C sky130_fd_sc_hd__or2_4
X_12768_ _12759_/A _12768_/B VGND VGND VPWR VPWR _12768_/X sky130_fd_sc_hd__or2_4
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12665__B _12665_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14507_/A VGND VGND VPWR VPWR _14520_/A sky130_fd_sc_hd__buf_2
X_18275_ _18215_/X _18273_/X _18240_/X _18274_/X VGND VGND VPWR VPWR _18275_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11719_ _11706_/A VGND VGND VPWR VPWR _11720_/A sky130_fd_sc_hd__inv_2
X_15487_ _15487_/A _15487_/B VGND VGND VPWR VPWR _15487_/X sky130_fd_sc_hd__or2_4
X_12699_ _11935_/A _12699_/B _12698_/X VGND VGND VPWR VPWR _12699_/X sky130_fd_sc_hd__or3_4
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17226_ _18538_/A VGND VGND VPWR VPWR _18320_/A sky130_fd_sc_hd__buf_2
X_14438_ _12492_/A _14438_/B _14438_/C VGND VGND VPWR VPWR _14442_/B sky130_fd_sc_hd__and3_4
XANTENNA__24455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17249__A _18538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17157_ _14262_/X _17144_/X _17539_/A _17146_/X VGND VGND VPWR VPWR _17157_/X sky130_fd_sc_hd__o22a_4
X_14369_ _14369_/A _22346_/A VGND VGND VPWR VPWR _14369_/X sky130_fd_sc_hd__or2_4
XANTENNA__12681__A _12574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16108_ _16108_/A _24045_/Q VGND VGND VPWR VPWR _16110_/B sky130_fd_sc_hd__or2_4
XFILLER_116_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17088_ _17088_/A VGND VGND VPWR VPWR _17912_/A sky130_fd_sc_hd__inv_2
XFILLER_157_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21207__B2 _21202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16039_ _16062_/A _16039_/B VGND VGND VPWR VPWR _16039_/X sky130_fd_sc_hd__or2_4
XFILLER_69_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20966__B1 _19773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22707__A1 _20531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22707__B2 _22705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19729_ _19659_/Y _19727_/X _19859_/A _19728_/X VGND VGND VPWR VPWR _19729_/X sky130_fd_sc_hd__a211o_4
XFILLER_38_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22183__A2 _22180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22740_ _19223_/A VGND VGND VPWR VPWR _23048_/A sky130_fd_sc_hd__inv_2
XFILLER_168_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22671_ _22459_/X _22665_/X _23136_/Q _22669_/X VGND VGND VPWR VPWR _22671_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12856__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16328__A _11684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11760__A _11759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21622_ _21544_/X _21620_/X _16102_/B _21617_/X VGND VGND VPWR VPWR _23757_/D sky130_fd_sc_hd__o22a_4
X_24410_ _24419_/CLK _24410_/D HRESETn VGND VGND VPWR VPWR _24410_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21553_ _21268_/A VGND VGND VPWR VPWR _21553_/X sky130_fd_sc_hd__buf_2
X_24341_ _24357_/CLK _24341_/D HRESETn VGND VGND VPWR VPWR _19126_/A sky130_fd_sc_hd__dfstp_4
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23509__CLK _23509_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20504_ _20398_/X _20488_/X _20714_/A _20503_/Y VGND VGND VPWR VPWR _20504_/X sky130_fd_sc_hd__a211o_4
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24272_ _24158_/CLK _19341_/X HRESETn VGND VGND VPWR VPWR _24272_/Q sky130_fd_sc_hd__dfrtp_4
X_21484_ _21254_/X _21478_/X _16301_/B _21482_/X VGND VGND VPWR VPWR _23823_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19639__A1 _20776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14790__B _14716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23223_ _23904_/CLK _22533_/X VGND VGND VPWR VPWR _15172_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13687__A _13687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20435_ _18101_/X _20260_/X _20341_/X _20434_/Y VGND VGND VPWR VPWR _20435_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17159__A _12093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21446__B2 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24125__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16063__A _16047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24091__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21997__A2 _21996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23154_ _23537_/CLK _23154_/D VGND VGND VPWR VPWR _16661_/B sky130_fd_sc_hd__dfxtp_4
X_20366_ _24433_/Q _18837_/B _24465_/Q _20282_/X VGND VGND VPWR VPWR _20366_/X sky130_fd_sc_hd__o22a_4
XFILLER_134_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22105_ _22420_/A VGND VGND VPWR VPWR _22105_/X sky130_fd_sc_hd__buf_2
XFILLER_134_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23085_ _20216_/D _23084_/Y VGND VGND VPWR VPWR HWRITE sky130_fd_sc_hd__and2_4
X_20297_ _20358_/A _20232_/X _20295_/X _24244_/Q _20334_/A VGND VGND VPWR VPWR _20298_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21749__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22036_ _21883_/X _22031_/X _14850_/B _22000_/A VGND VGND VPWR VPWR _23510_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21409__A _21388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20313__A _20257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11935__A _11935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17822__B1 _17820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15407__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23987_ _23889_/CLK _23987_/D VGND VGND VPWR VPWR _23987_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12111__A1 _12027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13740_ _12597_/A _13734_/X _13739_/X VGND VGND VPWR VPWR _13740_/X sky130_fd_sc_hd__or3_4
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22938_ _18643_/X _22938_/B VGND VGND VPWR VPWR _22938_/X sky130_fd_sc_hd__or2_4
XFILLER_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20185__A1 _24462_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21921__A2 _21916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13671_ _12191_/A _13760_/B VGND VGND VPWR VPWR _13673_/B sky130_fd_sc_hd__or2_4
X_22869_ _14483_/Y _22800_/Y _22815_/X VGND VGND VPWR VPWR _22869_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16238__A _11815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11670__A _13566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15410_ _13639_/A _15481_/B VGND VGND VPWR VPWR _15410_/X sky130_fd_sc_hd__or2_4
XFILLER_25_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15142__A _14574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12622_ _12621_/X VGND VGND VPWR VPWR _12975_/A sky130_fd_sc_hd__buf_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16390_ _16007_/X _16390_/B VGND VGND VPWR VPWR _16390_/X sky130_fd_sc_hd__or2_4
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24364__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20488__A2 _20866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15341_ _13695_/A _15339_/X _15341_/C VGND VGND VPWR VPWR _15345_/B sky130_fd_sc_hd__and3_4
X_12553_ _12515_/A _12551_/X _12553_/C VGND VGND VPWR VPWR _12554_/C sky130_fd_sc_hd__and3_4
XANTENNA__21685__B2 _21681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14981__A _11812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23189__CLK _23904_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18453__A _18399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_20_0_HCLK clkbuf_6_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_20_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18060_ _18008_/A VGND VGND VPWR VPWR _18060_/X sky130_fd_sc_hd__buf_2
XANTENNA__24434__CLK _23409_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15796__B _15796_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15272_ _14272_/A _15270_/X _15271_/X VGND VGND VPWR VPWR _15272_/X sky130_fd_sc_hd__and3_4
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ _12484_/A VGND VGND VPWR VPWR _12485_/A sky130_fd_sc_hd__buf_2
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17011_ _17011_/A VGND VGND VPWR VPWR _17011_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14223_ _11674_/A _14223_/B _14222_/X VGND VGND VPWR VPWR _14223_/X sky130_fd_sc_hd__or3_4
XANTENNA__21437__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14154_ _14154_/A _23487_/Q VGND VGND VPWR VPWR _14154_/X sky130_fd_sc_hd__or2_4
XFILLER_98_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14205__B _23583_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13105_ _13089_/A _13105_/B VGND VGND VPWR VPWR _13105_/X sky130_fd_sc_hd__or2_4
XFILLER_152_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18962_ _20192_/A VGND VGND VPWR VPWR _19016_/A sky130_fd_sc_hd__buf_2
X_14085_ _14086_/A _14084_/X VGND VGND VPWR VPWR _14085_/X sky130_fd_sc_hd__and2_4
XANTENNA__12006__A _12001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13036_ _12569_/A _23656_/Q VGND VGND VPWR VPWR _13037_/C sky130_fd_sc_hd__or2_4
X_17913_ _18406_/A _17913_/B VGND VGND VPWR VPWR _17913_/X sky130_fd_sc_hd__and2_4
X_18893_ _18893_/A VGND VGND VPWR VPWR _18894_/B sky130_fd_sc_hd__buf_2
XANTENNA__20223__A _20772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11845__A _11792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20412__A2 _20305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15317__A _11654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17844_ _17229_/X _17840_/X _17823_/X _17843_/X VGND VGND VPWR VPWR _17845_/A sky130_fd_sc_hd__o22a_4
XANTENNA__14221__A _13865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17775_ _17769_/X _17770_/Y _17775_/C _17775_/D VGND VGND VPWR VPWR _17775_/X sky130_fd_sc_hd__or4_4
X_14987_ _14897_/X _14985_/X _14986_/X VGND VGND VPWR VPWR _14987_/X sky130_fd_sc_hd__and3_4
X_19514_ _19514_/A VGND VGND VPWR VPWR _19514_/Y sky130_fd_sc_hd__inv_2
X_16726_ _16592_/A _16726_/B _16726_/C VGND VGND VPWR VPWR _16726_/X sky130_fd_sc_hd__or3_4
X_13938_ _14375_/A _13936_/X _13938_/C VGND VGND VPWR VPWR _13942_/B sky130_fd_sc_hd__and3_4
XFILLER_75_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21912__A2 _21909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20715__A3 _20712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19445_ _19445_/A VGND VGND VPWR VPWR _19446_/A sky130_fd_sc_hd__buf_2
X_16657_ _16676_/A _23634_/Q VGND VGND VPWR VPWR _16657_/X sky130_fd_sc_hd__or2_4
XANTENNA__17251__B _17251_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12676__A _12676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13869_ _13877_/A VGND VGND VPWR VPWR _13885_/A sky130_fd_sc_hd__buf_2
XANTENNA__16148__A _16148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_102_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR _23523_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__11580__A _24468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15608_ _13923_/A _15605_/X _15607_/X VGND VGND VPWR VPWR _15608_/X sky130_fd_sc_hd__and3_4
X_19376_ _19324_/A VGND VGND VPWR VPWR _19377_/A sky130_fd_sc_hd__buf_2
X_16588_ _16588_/A _16588_/B _16588_/C VGND VGND VPWR VPWR _16592_/B sky130_fd_sc_hd__and3_4
XFILLER_76_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18327_ _17697_/B _18302_/X _17697_/B _18302_/X VGND VGND VPWR VPWR _18327_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15539_ _14420_/A _15539_/B VGND VGND VPWR VPWR _15541_/B sky130_fd_sc_hd__or2_4
XANTENNA__19459__A HRDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21676__B2 _21674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22873__B1 _22799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14891__A _14110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18258_ _18377_/A _17460_/X VGND VGND VPWR VPWR _18258_/Y sky130_fd_sc_hd__nor2_4
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17209_ _17114_/X _17207_/X _17119_/X _17208_/X VGND VGND VPWR VPWR _17209_/X sky130_fd_sc_hd__o22a_4
XFILLER_159_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21428__B2 _21424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18189_ _18189_/A VGND VGND VPWR VPWR _18217_/C sky130_fd_sc_hd__inv_2
XFILLER_128_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13300__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21979__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20220_ _20220_/A VGND VGND VPWR VPWR _21184_/D sky130_fd_sc_hd__buf_2
X_20151_ _18706_/Y _19959_/A _20150_/X VGND VGND VPWR VPWR _20152_/B sky130_fd_sc_hd__o21a_4
XFILLER_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16611__A _16611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20082_ _20064_/X _18533_/A _20070_/X _20081_/X VGND VGND VPWR VPWR _20082_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20939__B1 _14751_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23910_ _23397_/CLK _23910_/D VGND VGND VPWR VPWR _13309_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_131_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19922__A _19438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14131__A _14131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23841_ _23744_/CLK _23841_/D VGND VGND VPWR VPWR _15560_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18538__A _18538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20984_ _20864_/A _20982_/X _20983_/X HRDATA[9] _20869_/A VGND VGND VPWR VPWR _20984_/X
+ sky130_fd_sc_hd__a32o_4
X_23772_ _23772_/CLK _21586_/X VGND VGND VPWR VPWR _23772_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21903__A2 _21902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22723_ _20801_/A _22722_/X _23103_/Q _22719_/X VGND VGND VPWR VPWR _23103_/D sky130_fd_sc_hd__o22a_4
XPHY_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__A _12634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23331__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21899__A _21899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22654_ _22430_/X _22651_/X _12389_/B _22648_/X VGND VGND VPWR VPWR _22654_/X sky130_fd_sc_hd__o22a_4
XFILLER_142_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21605_ _21133_/A VGND VGND VPWR VPWR _21706_/C sky130_fd_sc_hd__buf_2
XANTENNA__24306__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22585_ _22484_/X _22558_/A _15059_/B _22548_/A VGND VGND VPWR VPWR _22585_/X sky130_fd_sc_hd__o22a_4
XFILLER_21_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24324_ _24292_/CLK _19194_/X HRESETn VGND VGND VPWR VPWR _24324_/Q sky130_fd_sc_hd__dfrtp_4
X_21536_ _21821_/A VGND VGND VPWR VPWR _21536_/X sky130_fd_sc_hd__buf_2
XFILLER_21_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24255_ _24137_/CLK _24255_/D HRESETn VGND VGND VPWR VPWR _24255_/Q sky130_fd_sc_hd__dfrtp_4
X_21467_ _21313_/X _21462_/X _14959_/B _21431_/A VGND VGND VPWR VPWR _23830_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14306__A _12445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20418_ _20533_/A VGND VGND VPWR VPWR _20418_/X sky130_fd_sc_hd__buf_2
X_23206_ _24039_/CLK _23206_/D VGND VGND VPWR VPWR _13283_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18296__B1 _18168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21398_ _21391_/A VGND VGND VPWR VPWR _21398_/X sky130_fd_sc_hd__buf_2
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24186_ _24182_/CLK _19887_/X HRESETn VGND VGND VPWR VPWR _17016_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14025__B _23200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23137_ _23617_/CLK _23137_/D VGND VGND VPWR VPWR _15559_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20642__A2 HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20349_ _20349_/A VGND VGND VPWR VPWR _20349_/X sky130_fd_sc_hd__buf_2
XFILLER_150_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16521__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23068_ _23078_/A _17788_/Y VGND VGND VPWR VPWR _23070_/B sky130_fd_sc_hd__or2_4
XFILLER_122_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22395__A2 _22390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22019_ _21853_/X _22017_/X _15790_/B _22014_/X VGND VGND VPWR VPWR _22019_/X sky130_fd_sc_hd__o22a_4
X_14910_ _15281_/A _14886_/X _14893_/X _14901_/X _14909_/X VGND VGND VPWR VPWR _14910_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11665__A _15616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15890_ _13542_/A _15890_/B _15889_/X VGND VGND VPWR VPWR _15894_/B sky130_fd_sc_hd__and3_4
XFILLER_76_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14041__A _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14841_ _14841_/A _14833_/X _14841_/C VGND VGND VPWR VPWR _14842_/C sky130_fd_sc_hd__and3_4
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13880__A _14335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17560_ _17556_/Y _17024_/A _17031_/A _17660_/B VGND VGND VPWR VPWR _17561_/B sky130_fd_sc_hd__o22a_4
X_14772_ _14772_/A VGND VGND VPWR VPWR _14773_/A sky130_fd_sc_hd__buf_2
XFILLER_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11984_ _11973_/X VGND VGND VPWR VPWR _11984_/X sky130_fd_sc_hd__buf_2
X_16511_ _16362_/X _16511_/B _16511_/C VGND VGND VPWR VPWR _16519_/B sky130_fd_sc_hd__or3_4
X_13723_ _13752_/A _13721_/X _13722_/X VGND VGND VPWR VPWR _13723_/X sky130_fd_sc_hd__and3_4
XFILLER_95_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17491_ _13485_/X VGND VGND VPWR VPWR _17491_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12496__A _13666_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19230_ _19230_/A _19313_/A VGND VGND VPWR VPWR _19230_/X sky130_fd_sc_hd__and2_4
X_16442_ _16401_/X _16442_/B VGND VGND VPWR VPWR _16442_/X sky130_fd_sc_hd__or2_4
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13654_ _12502_/A VGND VGND VPWR VPWR _13655_/A sky130_fd_sc_hd__buf_2
XANTENNA__15303__C _15302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12605_ _12650_/A VGND VGND VPWR VPWR _12953_/A sky130_fd_sc_hd__buf_2
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19161_ _19161_/A VGND VGND VPWR VPWR _20266_/A sky130_fd_sc_hd__inv_2
X_16373_ _16314_/X _16371_/X _16372_/X VGND VGND VPWR VPWR _16373_/X sky130_fd_sc_hd__and3_4
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _16831_/A _16831_/B VGND VGND VPWR VPWR _13585_/X sky130_fd_sc_hd__or2_4
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18112_ _23043_/B _18111_/X _23043_/B _18111_/X VGND VGND VPWR VPWR _18112_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19720__B1 _17811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15324_ _15324_/A _15324_/B _15324_/C VGND VGND VPWR VPWR _15324_/X sky130_fd_sc_hd__and3_4
XANTENNA__15600__A _13894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12536_ _12536_/A _12536_/B _12536_/C VGND VGND VPWR VPWR _12536_/X sky130_fd_sc_hd__and3_4
X_19092_ _19082_/X _19091_/X _19082_/X _11523_/A VGND VGND VPWR VPWR _24349_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20330__A1 _17650_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20218__A _20218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18043_ _18043_/A VGND VGND VPWR VPWR _18043_/Y sky130_fd_sc_hd__inv_2
X_15255_ _14003_/A _15253_/X _15255_/C VGND VGND VPWR VPWR _15259_/B sky130_fd_sc_hd__and3_4
X_12467_ _12467_/A VGND VGND VPWR VPWR _12468_/A sky130_fd_sc_hd__buf_2
XFILLER_173_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13120__A _12762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14206_ _14191_/A _14206_/B _14205_/X VGND VGND VPWR VPWR _14213_/B sky130_fd_sc_hd__and3_4
XFILLER_144_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12020__B1 _11608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15186_ _14773_/A _15122_/B VGND VGND VPWR VPWR _15188_/B sky130_fd_sc_hd__or2_4
XANTENNA__22083__B2 _22078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22433__A _22433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12398_ _12407_/A _12398_/B VGND VGND VPWR VPWR _12398_/X sky130_fd_sc_hd__or2_4
XFILLER_158_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14137_ _14137_/A _23903_/Q VGND VGND VPWR VPWR _14139_/B sky130_fd_sc_hd__or2_4
XANTENNA__21830__B2 _21822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19994_ _19950_/X VGND VGND VPWR VPWR _19994_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_27_0_HCLK clkbuf_6_13_0_HCLK/X VGND VGND VPWR VPWR _24368_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__23204__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18945_ _24369_/Q VGND VGND VPWR VPWR _18948_/A sky130_fd_sc_hd__inv_2
X_14068_ _14056_/A _14068_/B VGND VGND VPWR VPWR _14068_/X sky130_fd_sc_hd__or2_4
XANTENNA__22386__A2 _22383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13019_ _12487_/A _23976_/Q VGND VGND VPWR VPWR _13019_/X sky130_fd_sc_hd__or2_4
XFILLER_100_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20397__A1 _20302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18876_ _17272_/X _18870_/X _24412_/Q _18871_/X VGND VGND VPWR VPWR _18876_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20397__B2 _20396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17827_ _17233_/X _17147_/X _17231_/X _17154_/X VGND VGND VPWR VPWR _17827_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22138__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13790__A _13954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17262__A _17398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17758_ _17758_/A _17744_/X _17757_/X VGND VGND VPWR VPWR _17758_/X sky130_fd_sc_hd__and3_4
XFILLER_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16709_ _16732_/A _16707_/X _16709_/C VGND VGND VPWR VPWR _16710_/C sky130_fd_sc_hd__and3_4
XANTENNA__21897__B2 _21892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17689_ _17691_/A _17688_/X VGND VGND VPWR VPWR _17689_/X sky130_fd_sc_hd__or2_4
XFILLER_63_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19428_ _19428_/A VGND VGND VPWR VPWR _19428_/X sky130_fd_sc_hd__buf_2
XANTENNA__24470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22608__A _22608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21649__A1 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19359_ _19354_/X _18429_/X _19358_/X _20654_/A VGND VGND VPWR VPWR _24260_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21649__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22310__A2 _22308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22370_ _22110_/X _22369_/X _23310_/Q _22366_/X VGND VGND VPWR VPWR _23310_/D sky130_fd_sc_hd__o22a_4
XFILLER_148_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21321_ _21320_/X VGND VGND VPWR VPWR _21322_/A sky130_fd_sc_hd__buf_2
XFILLER_136_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13030__A _12570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24040_ _23337_/CLK _24040_/D VGND VGND VPWR VPWR _24040_/Q sky130_fd_sc_hd__dfxtp_4
X_21252_ _21239_/X VGND VGND VPWR VPWR _21252_/X sky130_fd_sc_hd__buf_2
XFILLER_117_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14551__A2 _14548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20203_ _18742_/X _20079_/X _20202_/Y _19951_/X VGND VGND VPWR VPWR _20203_/X sky130_fd_sc_hd__o22a_4
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13965__A _13965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21183_ _21183_/A VGND VGND VPWR VPWR _21183_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20134_ _20133_/Y _11553_/X _11549_/B VGND VGND VPWR VPWR _20134_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__22377__A2 _22376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20065_ _24482_/Q VGND VGND VPWR VPWR _20065_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17253__A1 _16687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17172__A _13417_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23824_ _23728_/CLK _23824_/D VGND VGND VPWR VPWR _16443_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ _23467_/CLK _23755_/D VGND VGND VPWR VPWR _23755_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _20964_/X _20966_/X _20262_/X VGND VGND VPWR VPWR _20967_/Y sky130_fd_sc_hd__o21ai_4
XPHY_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22706_ _20509_/A _22701_/X _12564_/B _22705_/X VGND VGND VPWR VPWR _23115_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13205__A _13205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17900__A _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20560__A1 _20533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23686_ _23397_/CLK _23686_/D VGND VGND VPWR VPWR _23686_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20560__B2 _20510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _20864_/X _20896_/X _20897_/X HRDATA[13] _20869_/X VGND VGND VPWR VPWR _20898_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_55_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21422__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24140__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22637_ _21806_/A _22173_/B _22637_/C _22637_/D VGND VGND VPWR VPWR _22637_/X sky130_fd_sc_hd__or4_4
XFILLER_139_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15420__A _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13370_ _13370_/A VGND VGND VPWR VPWR _13379_/A sky130_fd_sc_hd__buf_2
XFILLER_127_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22568_ _22454_/X _22565_/X _15399_/B _22562_/X VGND VGND VPWR VPWR _23202_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24307_ _24368_/CLK _24307_/D HRESETn VGND VGND VPWR VPWR _24307_/Q sky130_fd_sc_hd__dfrtp_4
X_12321_ _11659_/A VGND VGND VPWR VPWR _12322_/A sky130_fd_sc_hd__buf_2
XFILLER_166_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21519_ _21315_/X _21492_/A _15038_/B _21482_/A VGND VGND VPWR VPWR _21519_/X sky130_fd_sc_hd__o22a_4
XFILLER_154_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22499_ _22420_/X _22494_/X _16438_/B _22498_/X VGND VGND VPWR VPWR _22499_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15040_ _12474_/A _23701_/Q VGND VGND VPWR VPWR _15042_/B sky130_fd_sc_hd__or2_4
XANTENNA__22065__B2 _22064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12252_ _13677_/A VGND VGND VPWR VPWR _12279_/A sky130_fd_sc_hd__buf_2
X_24238_ _24158_/CLK _24238_/D HRESETn VGND VGND VPWR VPWR _24238_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13875__A _13888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12183_ _12183_/A VGND VGND VPWR VPWR _12183_/X sky130_fd_sc_hd__buf_2
XANTENNA__21812__B2 _21810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24169_ _23383_/CLK _24169_/D HRESETn VGND VGND VPWR VPWR _24169_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17492__A1 _16678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16991_ _17703_/A _16991_/B VGND VGND VPWR VPWR _16992_/B sky130_fd_sc_hd__or2_4
XANTENNA__22368__A2 _22362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15942_ _13327_/A VGND VGND VPWR VPWR _16011_/A sky130_fd_sc_hd__buf_2
X_18730_ _18731_/A _18729_/X VGND VGND VPWR VPWR _18730_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__23377__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20379__A1 _20302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20379__B2 _20225_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21576__B1 _23776_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21040__A2 _21038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18661_ _18661_/A _18630_/C VGND VGND VPWR VPWR _18661_/X sky130_fd_sc_hd__and2_4
XFILLER_23_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15873_ _13540_/X _15804_/B VGND VGND VPWR VPWR _15873_/X sky130_fd_sc_hd__or2_4
XFILLER_110_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17612_ _17412_/A VGND VGND VPWR VPWR _17612_/Y sky130_fd_sc_hd__inv_2
X_14824_ _14693_/A _14824_/B _14824_/C VGND VGND VPWR VPWR _14825_/C sky130_fd_sc_hd__and3_4
XANTENNA__24299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18592_ _17760_/X _17731_/X _17760_/X _17731_/X VGND VGND VPWR VPWR _18592_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17543_ _17145_/Y _17537_/Y _17490_/C _17542_/X VGND VGND VPWR VPWR _17544_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15314__B _15253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14755_ _12299_/A _14755_/B _14754_/X VGND VGND VPWR VPWR _14755_/X sky130_fd_sc_hd__and3_4
X_11967_ _11967_/A VGND VGND VPWR VPWR _15420_/A sky130_fd_sc_hd__buf_2
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13115__A _13091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13706_ _13706_/A VGND VGND VPWR VPWR _13751_/A sky130_fd_sc_hd__buf_2
X_17474_ _12320_/Y _17022_/X _17031_/A _17473_/Y VGND VGND VPWR VPWR _17475_/B sky130_fd_sc_hd__o22a_4
X_14686_ _14657_/A _14686_/B VGND VGND VPWR VPWR _14689_/B sky130_fd_sc_hd__or2_4
XANTENNA__22428__A _22113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11898_ _11898_/A VGND VGND VPWR VPWR _14421_/A sky130_fd_sc_hd__buf_2
XFILLER_32_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16425_ _16409_/A _16425_/B VGND VGND VPWR VPWR _16425_/X sky130_fd_sc_hd__or2_4
X_19213_ _19213_/A VGND VGND VPWR VPWR _19213_/Y sky130_fd_sc_hd__inv_2
X_13637_ _13637_/A VGND VGND VPWR VPWR _15447_/A sky130_fd_sc_hd__buf_2
XANTENNA__12954__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16426__A _15998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19144_ _19144_/A _19143_/X VGND VGND VPWR VPWR _19144_/X sky130_fd_sc_hd__and2_4
X_16356_ _16313_/A _16356_/B _16355_/X VGND VGND VPWR VPWR _16356_/X sky130_fd_sc_hd__and3_4
XFILLER_73_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13568_ _13567_/X VGND VGND VPWR VPWR _13583_/A sky130_fd_sc_hd__inv_2
XFILLER_9_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15307_ _13952_/A _15307_/B VGND VGND VPWR VPWR _15309_/B sky130_fd_sc_hd__or2_4
X_12519_ _12870_/A _12517_/X _12518_/X VGND VGND VPWR VPWR _12523_/B sky130_fd_sc_hd__and3_4
X_19075_ _19075_/A VGND VGND VPWR VPWR _19075_/Y sky130_fd_sc_hd__inv_2
X_16287_ _16287_/A _16287_/B VGND VGND VPWR VPWR _16287_/X sky130_fd_sc_hd__or2_4
XFILLER_173_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13499_ _12954_/A VGND VGND VPWR VPWR _13520_/A sky130_fd_sc_hd__buf_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18026_ _24212_/Q VGND VGND VPWR VPWR _18026_/X sky130_fd_sc_hd__buf_2
X_15238_ _14248_/A _15180_/B VGND VGND VPWR VPWR _15239_/C sky130_fd_sc_hd__or2_4
XANTENNA__22056__B2 _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22163__A _20958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24152__CLK _24302_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17257__A _17255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15169_ _14295_/A _15169_/B VGND VGND VPWR VPWR _15169_/X sky130_fd_sc_hd__or2_4
XANTENNA__21803__B2 _21767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18680__B1 _17648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19977_ _16935_/X _19976_/X _17653_/X _19331_/X VGND VGND VPWR VPWR _19977_/X sky130_fd_sc_hd__o22a_4
XFILLER_80_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18928_ _18928_/A VGND VGND VPWR VPWR _18928_/X sky130_fd_sc_hd__buf_2
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21567__B1 _23780_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22178__A2_N _22177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18859_ _12980_/X _18856_/X _20541_/A _18857_/X VGND VGND VPWR VPWR _18859_/X sky130_fd_sc_hd__o22a_4
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15505__A _12626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21870_ _21834_/A VGND VGND VPWR VPWR _21870_/X sky130_fd_sc_hd__buf_2
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20821_ HRDATA[8] _20668_/A VGND VGND VPWR VPWR _20821_/X sky130_fd_sc_hd__or2_4
XFILLER_51_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13025__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23540_ _23668_/CLK _21994_/X VGND VGND VPWR VPWR _23540_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20752_ _20641_/X _20751_/X _20639_/X VGND VGND VPWR VPWR _20752_/Y sky130_fd_sc_hd__o21ai_4
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23471_ _23119_/CLK _22109_/X VGND VGND VPWR VPWR _16274_/B sky130_fd_sc_hd__dfxtp_4
X_20683_ _20540_/X _20682_/X _19053_/A _20547_/X VGND VGND VPWR VPWR _20683_/X sky130_fd_sc_hd__o22a_4
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12864__A _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15240__A _14615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21098__A2 _21097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22422_ _22420_/X _22414_/X _16387_/B _22421_/X VGND VGND VPWR VPWR _22422_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22295__B2 _22291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19647__A _19888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22353_ _15003_/B VGND VGND VPWR VPWR _23317_/D sky130_fd_sc_hd__buf_2
XANTENNA__17171__B1 _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21304_ _21304_/A VGND VGND VPWR VPWR _21304_/X sky130_fd_sc_hd__buf_2
X_22284_ _22284_/A VGND VGND VPWR VPWR _22284_/X sky130_fd_sc_hd__buf_2
XANTENNA__22047__B2 _22043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24023_ _23416_/CLK _24023_/D VGND VGND VPWR VPWR _15134_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13695__A _13695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21235_ _22537_/D VGND VGND VPWR VPWR _21236_/D sky130_fd_sc_hd__buf_2
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17474__A1 _12320_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21270__A2 _21269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21166_ _21152_/A VGND VGND VPWR VPWR _21166_/X sky130_fd_sc_hd__buf_2
XANTENNA__17474__B2 _17473_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20117_ _19433_/X _20116_/X _19399_/X _24136_/Q VGND VGND VPWR VPWR _24136_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_10_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR _23476_/CLK sky130_fd_sc_hd__clkbuf_1
X_21097_ _21104_/A VGND VGND VPWR VPWR _21097_/X sky130_fd_sc_hd__buf_2
XANTENNA__12104__A _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_73_0_HCLK clkbuf_7_72_0_HCLK/A VGND VGND VPWR VPWR _23192_/CLK sky130_fd_sc_hd__clkbuf_1
X_20048_ _18354_/X _20031_/X _20047_/Y _20042_/X VGND VGND VPWR VPWR _20048_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21022__A2 _20358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18423__B1 _18168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11943__A _16116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15415__A _15415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12870_ _12870_/A VGND VGND VPWR VPWR _12873_/A sky130_fd_sc_hd__buf_2
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11821_ _11833_/A _24084_/Q VGND VGND VPWR VPWR _11821_/X sky130_fd_sc_hd__or2_4
X_23807_ _23101_/CLK _23807_/D VGND VGND VPWR VPWR _23807_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24321__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21999_ _21819_/X _21996_/X _23537_/Q _21993_/X VGND VGND VPWR VPWR _21999_/X sky130_fd_sc_hd__o22a_4
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14540_/A _14540_/B _14540_/C VGND VGND VPWR VPWR _14544_/B sky130_fd_sc_hd__and3_4
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11752_/A VGND VGND VPWR VPWR _11753_/A sky130_fd_sc_hd__buf_2
X_23738_ _24090_/CLK _23738_/D VGND VGND VPWR VPWR _14627_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21325__A2_N _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22248__A _22226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21152__A _21152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _11880_/A _14469_/X _14470_/X VGND VGND VPWR VPWR _14471_/X sky130_fd_sc_hd__and3_4
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _13123_/A VGND VGND VPWR VPWR _13415_/A sky130_fd_sc_hd__buf_2
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23669_ _23456_/CLK _23669_/D VGND VGND VPWR VPWR _23669_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16210_/A _16208_/X _16210_/C VGND VGND VPWR VPWR _16210_/X sky130_fd_sc_hd__and3_4
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _13455_/A _23365_/Q VGND VGND VPWR VPWR _13422_/X sky130_fd_sc_hd__or2_4
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15150__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17190_ _17113_/X _17185_/X _17128_/X _17189_/X VGND VGND VPWR VPWR _17190_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__22286__B2 _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24175__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16141_ _16110_/A _16139_/X _16141_/C VGND VGND VPWR VPWR _16145_/B sky130_fd_sc_hd__and3_4
X_13353_ _13375_/A _13280_/B VGND VGND VPWR VPWR _13354_/C sky130_fd_sc_hd__or2_4
XFILLER_154_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12304_ _12304_/A VGND VGND VPWR VPWR _12747_/A sky130_fd_sc_hd__buf_2
X_16072_ _16048_/A _23726_/Q VGND VGND VPWR VPWR _16072_/X sky130_fd_sc_hd__or2_4
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13284_ _12561_/A _23782_/Q VGND VGND VPWR VPWR _13284_/X sky130_fd_sc_hd__or2_4
XFILLER_170_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19900_ _19700_/A _19898_/X _19899_/X _16927_/Y _19552_/X VGND VGND VPWR VPWR _19900_/X
+ sky130_fd_sc_hd__a32o_4
X_15023_ _15000_/A _23125_/Q VGND VGND VPWR VPWR _15023_/X sky130_fd_sc_hd__or2_4
XFILLER_155_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12235_ _13687_/A VGND VGND VPWR VPWR _12236_/A sky130_fd_sc_hd__buf_2
XANTENNA__17077__A _17077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19831_ _19831_/A VGND VGND VPWR VPWR _19831_/Y sky130_fd_sc_hd__inv_2
X_12166_ _12166_/A _23731_/Q VGND VGND VPWR VPWR _12168_/B sky130_fd_sc_hd__or2_4
XFILLER_111_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17465__B2 _17464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19762_ _19890_/A _19742_/X VGND VGND VPWR VPWR _19762_/X sky130_fd_sc_hd__or2_4
XANTENNA__17805__A _17109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12014__A _11960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16974_ _24137_/Q VGND VGND VPWR VPWR _17734_/A sky130_fd_sc_hd__inv_2
X_12097_ _12105_/A VGND VGND VPWR VPWR _12097_/X sky130_fd_sc_hd__buf_2
XANTENNA__21327__A _21341_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18713_ _18518_/X _17623_/A _18519_/X VGND VGND VPWR VPWR _18713_/X sky130_fd_sc_hd__a21o_4
XANTENNA__19611__C1 _19576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17524__B _17522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15925_ _15518_/X _15655_/Y _15519_/X VGND VGND VPWR VPWR _15925_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__22210__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20231__A _20231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19693_ _19744_/A VGND VGND VPWR VPWR _19879_/D sky130_fd_sc_hd__buf_2
XANTENNA__24409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12949__A _12949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15856_ _15894_/A _15852_/X _15856_/C VGND VGND VPWR VPWR _15856_/X sky130_fd_sc_hd__or3_4
X_18644_ _16943_/A _18633_/X _17013_/X _18643_/X VGND VGND VPWR VPWR _18644_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12668__B _12668_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14807_ _14679_/A _14724_/B VGND VGND VPWR VPWR _14808_/C sky130_fd_sc_hd__or2_4
X_18575_ _17006_/A _16976_/X _16977_/X VGND VGND VPWR VPWR _18575_/X sky130_fd_sc_hd__a21bo_4
X_15787_ _15717_/X _15786_/Y VGND VGND VPWR VPWR _15787_/X sky130_fd_sc_hd__and2_4
X_12999_ _12906_/A _12999_/B VGND VGND VPWR VPWR _12999_/X sky130_fd_sc_hd__or2_4
XANTENNA__14451__A1 _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22513__A2 _22508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17526_ _17605_/D VGND VGND VPWR VPWR _17527_/D sky130_fd_sc_hd__inv_2
X_14738_ _15415_/A _14736_/X _14737_/X VGND VGND VPWR VPWR _14738_/X sky130_fd_sc_hd__and3_4
XFILLER_33_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22158__A _22158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17457_ _17453_/Y _17021_/X _17029_/X _17456_/Y VGND VGND VPWR VPWR _17460_/B sky130_fd_sc_hd__o22a_4
XFILLER_20_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14669_ _14669_/A VGND VGND VPWR VPWR _14679_/A sky130_fd_sc_hd__buf_2
X_16408_ _16402_/X _22326_/A VGND VGND VPWR VPWR _16408_/X sky130_fd_sc_hd__or2_4
XANTENNA__15060__A _12329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17388_ _11643_/Y _17378_/A _17358_/Y VGND VGND VPWR VPWR _17389_/B sky130_fd_sc_hd__o21a_4
XANTENNA__11568__A2 IRQ[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15995__A _15967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16339_ _16318_/A _16339_/B VGND VGND VPWR VPWR _16339_/X sky130_fd_sc_hd__or2_4
X_19127_ _24373_/Q _19106_/X VGND VGND VPWR VPWR _19127_/Y sky130_fd_sc_hd__nor2_4
XFILLER_158_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22029__A1 _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19058_ _19052_/X _19057_/X _19052_/X _19053_/A VGND VGND VPWR VPWR _24355_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22029__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18009_ _18176_/A VGND VGND VPWR VPWR _18009_/X sky130_fd_sc_hd__buf_2
XFILLER_145_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21020_ _20305_/X _21011_/Y _21018_/X _21019_/Y _20255_/A VGND VGND VPWR VPWR _21020_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15219__B _15155_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17208__A1 _12982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22971_ _22961_/A _18480_/X VGND VGND VPWR VPWR _22974_/B sky130_fd_sc_hd__nand2_4
XANTENNA__12859__A _12884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21922_ _21860_/X _21916_/X _23584_/Q _21920_/X VGND VGND VPWR VPWR _23584_/D sky130_fd_sc_hd__o22a_4
XFILLER_83_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21853_ _21283_/A VGND VGND VPWR VPWR _21853_/X sky130_fd_sc_hd__buf_2
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18708__A1 _17974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22504__A2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19905__B1 _17087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20804_ _20422_/B _20844_/B VGND VGND VPWR VPWR _20804_/X sky130_fd_sc_hd__or2_4
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21784_ _21770_/A VGND VGND VPWR VPWR _21784_/X sky130_fd_sc_hd__buf_2
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23523_ _23523_/CLK _22019_/X VGND VGND VPWR VPWR _15790_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20735_ _20540_/X _20734_/X _19063_/A _20547_/X VGND VGND VPWR VPWR _20735_/X sky130_fd_sc_hd__o22a_4
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22268__B2 _22262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23454_ _23101_/CLK _23454_/D VGND VGND VPWR VPWR _13738_/B sky130_fd_sc_hd__dfxtp_4
X_20666_ _20871_/A _20665_/X VGND VGND VPWR VPWR _20670_/A sky130_fd_sc_hd__or2_4
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22405_ _22090_/A _22687_/B _22637_/C _22487_/B VGND VGND VPWR VPWR _22405_/X sky130_fd_sc_hd__or4_4
XFILLER_164_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19377__A _19377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20597_ _20533_/X _20596_/X _24103_/Q _20510_/X VGND VGND VPWR VPWR _20597_/X sky130_fd_sc_hd__o22a_4
X_23385_ _23772_/CLK _22267_/X VGND VGND VPWR VPWR _23385_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18281__A _18407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22336_ _13296_/B VGND VGND VPWR VPWR _23334_/D sky130_fd_sc_hd__buf_2
XANTENNA__21491__A2 _21485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22267_ _22161_/X _22265_/X _23385_/Q _22262_/X VGND VGND VPWR VPWR _22267_/X sky130_fd_sc_hd__o22a_4
X_24006_ _24102_/CLK _24006_/D VGND VGND VPWR VPWR _13294_/B sky130_fd_sc_hd__dfxtp_4
X_12020_ _11858_/X _11632_/X _11983_/X _11608_/X _12019_/X VGND VGND VPWR VPWR _12020_/X
+ sky130_fd_sc_hd__a32o_4
X_21218_ _20770_/X _21212_/X _23968_/Q _21216_/X VGND VGND VPWR VPWR _21218_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22198_ _22176_/A VGND VGND VPWR VPWR _22198_/X sky130_fd_sc_hd__buf_2
XANTENNA__15129__B _15129_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17625__A _18744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21149_ _20441_/X _21148_/X _24014_/Q _21145_/X VGND VGND VPWR VPWR _24014_/D sky130_fd_sc_hd__o22a_4
XFILLER_63_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13971_ _13630_/A _23552_/Q VGND VGND VPWR VPWR _13972_/C sky130_fd_sc_hd__or2_4
XFILLER_4_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15710_ _12301_/A _15708_/X _15710_/C VGND VGND VPWR VPWR _15710_/X sky130_fd_sc_hd__and3_4
XFILLER_4_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11673__A _11673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12922_ _12948_/A _12922_/B VGND VGND VPWR VPWR _12924_/B sky130_fd_sc_hd__or2_4
XANTENNA__15145__A _13589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16690_ _16586_/A _16751_/B VGND VGND VPWR VPWR _16692_/B sky130_fd_sc_hd__or2_4
XANTENNA__12488__B _12611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23415__CLK _23864_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15641_ _15641_/A _15566_/B VGND VGND VPWR VPWR _15641_/X sky130_fd_sc_hd__or2_4
X_12853_ _12884_/A _23369_/Q VGND VGND VPWR VPWR _12856_/B sky130_fd_sc_hd__or2_4
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_3_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR _24388_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11804_ _11792_/X _11804_/B VGND VGND VPWR VPWR _11804_/X sky130_fd_sc_hd__or2_4
X_18360_ _16982_/A VGND VGND VPWR VPWR _18367_/A sky130_fd_sc_hd__buf_2
XANTENNA__17360__A _17360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15572_ _12461_/A _15568_/X _15572_/C VGND VGND VPWR VPWR _15572_/X sky130_fd_sc_hd__or3_4
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12783_/X VGND VGND VPWR VPWR _12801_/A sky130_fd_sc_hd__buf_2
XFILLER_42_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17310_/X VGND VGND VPWR VPWR _17311_/Y sky130_fd_sc_hd__inv_2
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14516_/A _14523_/B VGND VGND VPWR VPWR _14523_/X sky130_fd_sc_hd__or2_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18291_ _17601_/X _18290_/X VGND VGND VPWR VPWR _18291_/X sky130_fd_sc_hd__and2_4
X_11735_ _11735_/A VGND VGND VPWR VPWR _11736_/A sky130_fd_sc_hd__buf_2
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _12077_/X _17240_/B VGND VGND VPWR VPWR _17880_/A sky130_fd_sc_hd__or2_4
X_14454_ _13011_/A _14452_/X _14454_/C VGND VGND VPWR VPWR _14454_/X sky130_fd_sc_hd__and3_4
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11665_/X VGND VGND VPWR VPWR _11666_/X sky130_fd_sc_hd__buf_2
XANTENNA__22259__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13379_/A _13405_/B VGND VGND VPWR VPWR _13406_/C sky130_fd_sc_hd__or2_4
XFILLER_128_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21610__A _21617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17173_ _17172_/X VGND VGND VPWR VPWR _17173_/Y sky130_fd_sc_hd__inv_2
X_14385_ _14385_/A VGND VGND VPWR VPWR _14509_/A sky130_fd_sc_hd__buf_2
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11597_ _11646_/A VGND VGND VPWR VPWR _11598_/D sky130_fd_sc_hd__inv_2
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12009__A _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16124_ _16096_/A VGND VGND VPWR VPWR _16156_/A sky130_fd_sc_hd__buf_2
X_13336_ _11902_/A _13405_/B VGND VGND VPWR VPWR _13336_/X sky130_fd_sc_hd__or2_4
XFILLER_143_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16055_ _16062_/A _23982_/Q VGND VGND VPWR VPWR _16056_/C sky130_fd_sc_hd__or2_4
XFILLER_115_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11848__A _16768_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13267_ _13049_/Y _13266_/X VGND VGND VPWR VPWR _13269_/A sky130_fd_sc_hd__and2_4
XANTENNA__14224__A _15362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15006_ _13663_/A _15002_/X _15005_/X VGND VGND VPWR VPWR _15006_/X sky130_fd_sc_hd__or3_4
XFILLER_68_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12218_ _12218_/A VGND VGND VPWR VPWR _13637_/A sky130_fd_sc_hd__buf_2
XANTENNA__11567__B IRQ[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22431__B2 _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13198_ _13052_/A VGND VGND VPWR VPWR _13220_/A sky130_fd_sc_hd__buf_2
XANTENNA__19734__B HRDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19814_ _19732_/X _19806_/X _19813_/X _16672_/A _19719_/X VGND VGND VPWR VPWR _19814_/X
+ sky130_fd_sc_hd__a32o_4
X_12149_ _16775_/A _23987_/Q VGND VGND VPWR VPWR _12150_/C sky130_fd_sc_hd__or2_4
XFILLER_155_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19745_ _19879_/C _19744_/X VGND VGND VPWR VPWR _19745_/X sky130_fd_sc_hd__and2_4
XANTENNA__13782__B _13781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16957_ _18250_/A VGND VGND VPWR VPWR _16987_/A sky130_fd_sc_hd__inv_2
XANTENNA__24243__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12679__A _12678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18938__A1 _14844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22734__A2 _22729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15055__A _15076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15908_ _13503_/X _15906_/X _15907_/X VGND VGND VPWR VPWR _15909_/C sky130_fd_sc_hd__and3_4
X_19676_ _19538_/A VGND VGND VPWR VPWR _19677_/A sky130_fd_sc_hd__inv_2
X_16888_ _16533_/X _16823_/X _16533_/X _16823_/X VGND VGND VPWR VPWR _16888_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18627_ _17743_/A VGND VGND VPWR VPWR _18627_/X sky130_fd_sc_hd__buf_2
X_15839_ _12890_/A _15835_/X _15839_/C VGND VGND VPWR VPWR _15839_/X sky130_fd_sc_hd__or3_4
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18558_ _18509_/X VGND VGND VPWR VPWR _18558_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17509_ _17508_/X VGND VGND VPWR VPWR _17509_/Y sky130_fd_sc_hd__inv_2
X_18489_ _18198_/A _18287_/X VGND VGND VPWR VPWR _18489_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21170__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13303__A _13303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20520_ _20425_/X _20518_/X _19247_/A _20519_/X VGND VGND VPWR VPWR _20520_/X sky130_fd_sc_hd__o22a_4
XFILLER_165_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20451_ _20447_/X _20448_/Y _20450_/X _18997_/Y _20275_/X VGND VGND VPWR VPWR _20452_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_146_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17126__B1 _17015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16614__A _11792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23170_ _23204_/CLK _23170_/D VGND VGND VPWR VPWR _15473_/B sky130_fd_sc_hd__dfxtp_4
X_20382_ _20847_/A VGND VGND VPWR VPWR _20388_/A sky130_fd_sc_hd__buf_2
XANTENNA__22670__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17429__B _17429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11758__A _13414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22121_ _22120_/X _22111_/X _12797_/B _22118_/X VGND VGND VPWR VPWR _23466_/D sky130_fd_sc_hd__o22a_4
XFILLER_134_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19925__A _22745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14134__A _15281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22052_ _21824_/X _22046_/X _16293_/B _22050_/X VGND VGND VPWR VPWR _22052_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22422__B2 _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21003_ _22482_/A VGND VGND VPWR VPWR _21313_/A sky130_fd_sc_hd__buf_2
XFILLER_102_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17445__A _15651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12589__A _12925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18929__A1 _17161_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22725__A2 _22722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22954_ _22738_/A _18554_/Y VGND VGND VPWR VPWR _22954_/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21905_ _21831_/X _21902_/X _23596_/Q _21899_/X VGND VGND VPWR VPWR _23596_/D sky130_fd_sc_hd__o22a_4
XFILLER_83_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22885_ _22801_/X VGND VGND VPWR VPWR _22885_/X sky130_fd_sc_hd__buf_2
X_21836_ _20531_/A VGND VGND VPWR VPWR _21836_/X sky130_fd_sc_hd__buf_2
XFILLER_110_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21767_ _21767_/A VGND VGND VPWR VPWR _21767_/X sky130_fd_sc_hd__buf_2
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21161__B2 _21159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14309__A _12470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23506_ _23204_/CLK _23506_/D VGND VGND VPWR VPWR _23506_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _11520_/A _11519_/X VGND VGND VPWR VPWR _19099_/A sky130_fd_sc_hd__or2_4
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20718_ _20718_/A VGND VGND VPWR VPWR _21570_/A sky130_fd_sc_hd__buf_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24486_ _24271_/CLK _24486_/D HRESETn VGND VGND VPWR VPWR _20047_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22526__A _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21698_ _21658_/A VGND VGND VPWR VPWR _21698_/X sky130_fd_sc_hd__buf_2
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23437_ _23501_/CLK _22189_/X VGND VGND VPWR VPWR _16219_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20649_ _20644_/X _20648_/X _24292_/Q _20519_/X VGND VGND VPWR VPWR _20649_/X sky130_fd_sc_hd__o22a_4
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17117__B1 _16821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16524__A _16452_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14170_ _14170_/A _23871_/Q VGND VGND VPWR VPWR _14171_/C sky130_fd_sc_hd__or2_4
XANTENNA__21464__A2 _21462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23368_ _23656_/CLK _23368_/D VGND VGND VPWR VPWR _12991_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17339__B _17339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13867__B _13796_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22661__B2 _22655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20046__A _19956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13121_ _13099_/A _13119_/X _13120_/X VGND VGND VPWR VPWR _13122_/C sky130_fd_sc_hd__and3_4
XANTENNA__11668__A _11668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22319_ _22165_/X _22315_/X _15125_/B _22284_/A VGND VGND VPWR VPWR _23351_/D sky130_fd_sc_hd__o22a_4
X_23299_ _23523_/CLK _23299_/D VGND VGND VPWR VPWR _15800_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14044__A _13696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24213__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13052_ _13052_/A VGND VGND VPWR VPWR _13053_/A sky130_fd_sc_hd__buf_2
XFILLER_133_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12003_ _11905_/X VGND VGND VPWR VPWR _12015_/A sky130_fd_sc_hd__buf_2
XFILLER_65_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17355__A _17418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13883__A _12336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17860_ _17837_/X _17212_/X _17838_/X _17214_/X VGND VGND VPWR VPWR _17860_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24387__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16811_ _16811_/A _24113_/Q VGND VGND VPWR VPWR _16811_/X sky130_fd_sc_hd__or2_4
XFILLER_66_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12499__A _12499_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24363__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17791_ _18150_/A _17260_/A VGND VGND VPWR VPWR _17791_/X sky130_fd_sc_hd__or2_4
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22716__A2 _22715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19530_ _24172_/Q _19457_/A HRDATA[24] _19454_/A VGND VGND VPWR VPWR _19530_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_6_43_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_86_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13954_ _13954_/A _13952_/X _13954_/C VGND VGND VPWR VPWR _13954_/X sky130_fd_sc_hd__and3_4
X_16742_ _16742_/A _23825_/Q VGND VGND VPWR VPWR _16743_/C sky130_fd_sc_hd__or2_4
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21924__B1 _23583_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12905_ _12905_/A _12963_/B VGND VGND VPWR VPWR _12907_/B sky130_fd_sc_hd__or2_4
XANTENNA__23092__A _17060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16673_ _16677_/A _23890_/Q VGND VGND VPWR VPWR _16674_/C sky130_fd_sc_hd__or2_4
X_19461_ _19461_/A VGND VGND VPWR VPWR _19461_/X sky130_fd_sc_hd__buf_2
XANTENNA__21605__A _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13885_ _13885_/A _23773_/Q VGND VGND VPWR VPWR _13886_/C sky130_fd_sc_hd__or2_4
X_18412_ _17920_/X _18388_/Y _17944_/X _18411_/X VGND VGND VPWR VPWR _18412_/X sky130_fd_sc_hd__a211o_4
X_12836_ _13387_/A _12836_/B VGND VGND VPWR VPWR _12836_/X sky130_fd_sc_hd__or2_4
X_15624_ _15612_/A _15624_/B _15624_/C VGND VGND VPWR VPWR _15625_/C sky130_fd_sc_hd__and3_4
X_19392_ _19377_/A VGND VGND VPWR VPWR _19392_/X sky130_fd_sc_hd__buf_2
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15555_ _11886_/A _15555_/B VGND VGND VPWR VPWR _15555_/X sky130_fd_sc_hd__or2_4
XANTENNA__15322__B _15260_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18343_ _18411_/A _18343_/B VGND VGND VPWR VPWR _18343_/X sky130_fd_sc_hd__and2_4
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12767_ _12766_/X VGND VGND VPWR VPWR _13349_/A sky130_fd_sc_hd__buf_2
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19896__A2 _19724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13123__A _13123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14506_/A _14436_/B VGND VGND VPWR VPWR _14506_/X sky130_fd_sc_hd__or2_4
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18274_ _17683_/B _18181_/X _17683_/B _18181_/X VGND VGND VPWR VPWR _18274_/X sky130_fd_sc_hd__a2bb2o_4
X_11718_ _11717_/X _11718_/B VGND VGND VPWR VPWR _11718_/X sky130_fd_sc_hd__or2_4
X_15486_ _15486_/A _23906_/Q VGND VGND VPWR VPWR _15488_/B sky130_fd_sc_hd__or2_4
X_12698_ _12698_/A _12698_/B _12697_/X VGND VGND VPWR VPWR _12698_/X sky130_fd_sc_hd__and3_4
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14437_ _13010_/A _23995_/Q VGND VGND VPWR VPWR _14438_/C sky130_fd_sc_hd__or2_4
X_17225_ _17075_/X VGND VGND VPWR VPWR _18538_/A sky130_fd_sc_hd__buf_2
X_11649_ _11648_/X VGND VGND VPWR VPWR _16899_/A sky130_fd_sc_hd__inv_2
XANTENNA__12962__A _12962_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16434__A _15934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17156_ _17156_/A VGND VGND VPWR VPWR _17539_/A sky130_fd_sc_hd__inv_2
X_14368_ _14383_/A _14368_/B _14367_/X VGND VGND VPWR VPWR _14368_/X sky130_fd_sc_hd__and3_4
XFILLER_156_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22652__B2 _22648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16107_ _16144_/A _16107_/B _16107_/C VGND VGND VPWR VPWR _16107_/X sky130_fd_sc_hd__and3_4
XFILLER_116_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13319_ _13319_/A _23398_/Q VGND VGND VPWR VPWR _13319_/X sky130_fd_sc_hd__or2_4
X_17087_ _17087_/A _17188_/A _17075_/X VGND VGND VPWR VPWR _17088_/A sky130_fd_sc_hd__or3_4
XANTENNA__24495__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14299_ _13823_/A _14363_/B VGND VGND VPWR VPWR _14300_/C sky130_fd_sc_hd__or2_4
XANTENNA__21207__A2 _21205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16038_ _16061_/A _16038_/B VGND VGND VPWR VPWR _16038_/X sky130_fd_sc_hd__or2_4
XFILLER_112_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14889__A _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_125_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR _23592_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_112_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17989_ _17922_/X _17842_/X _17945_/X _17857_/X VGND VGND VPWR VPWR _17989_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22707__A2 _22701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19728_ _19724_/A _19691_/Y VGND VGND VPWR VPWR _19728_/X sky130_fd_sc_hd__and2_4
XANTENNA__12202__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19659_ _19649_/A VGND VGND VPWR VPWR _19659_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22670_ _22456_/X _22665_/X _15559_/B _22669_/X VGND VGND VPWR VPWR _23137_/D sky130_fd_sc_hd__o22a_4
X_21621_ _21541_/X _21620_/X _23758_/Q _21617_/X VGND VGND VPWR VPWR _21621_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21143__B2 _21138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13033__A _12569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24340_ _24277_/CLK _19163_/X HRESETn VGND VGND VPWR VPWR _19161_/A sky130_fd_sc_hd__dfrtp_4
X_21552_ _21551_/X _21542_/X _23786_/Q _21549_/X VGND VGND VPWR VPWR _21552_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21694__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20503_ _20502_/X VGND VGND VPWR VPWR _20503_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24271_ _24271_/CLK _24271_/D HRESETn VGND VGND VPWR VPWR _24271_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12872__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21483_ _21251_/X _21478_/X _16443_/B _21482_/X VGND VGND VPWR VPWR _23824_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16570__A1 _11868_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16344__A _13407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24236__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23222_ _23192_/CLK _22534_/X VGND VGND VPWR VPWR _23222_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21446__A2 _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20434_ _20388_/A _20433_/X VGND VGND VPWR VPWR _20434_/Y sky130_fd_sc_hd__nor2_4
XFILLER_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23153_ _23281_/CLK _23153_/D VGND VGND VPWR VPWR _16795_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_101_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20365_ _20251_/X _20364_/X _20235_/X VGND VGND VPWR VPWR _20365_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22104_ _22103_/X _22099_/X _16776_/B _22094_/X VGND VGND VPWR VPWR _22104_/X sky130_fd_sc_hd__o22a_4
XFILLER_134_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23084_ _23084_/A VGND VGND VPWR VPWR _23084_/Y sky130_fd_sc_hd__inv_2
X_20296_ _18597_/Y VGND VGND VPWR VPWR _20334_/A sky130_fd_sc_hd__buf_2
XFILLER_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22081__A _22041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24386__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22035_ _21881_/X _22031_/X _15123_/B _22000_/A VGND VGND VPWR VPWR _22035_/X sky130_fd_sc_hd__o22a_4
XFILLER_130_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14311__B _14387_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23986_ _23922_/CLK _23986_/D VGND VGND VPWR VPWR _23986_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12112__A _12111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12111__A2 _11633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22937_ _23079_/B VGND VGND VPWR VPWR _22938_/B sky130_fd_sc_hd__buf_2
XANTENNA__20185__A2 IRQ[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16519__A _11684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21382__B2 _21381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11951__A _11951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15423__A _15423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13670_ _12251_/A VGND VGND VPWR VPWR _15411_/A sky130_fd_sc_hd__buf_2
X_22868_ _22868_/A VGND VGND VPWR VPWR HWDATA[21] sky130_fd_sc_hd__inv_2
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12621_ _12604_/A VGND VGND VPWR VPWR _12621_/X sky130_fd_sc_hd__buf_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21819_ _21534_/A VGND VGND VPWR VPWR _21819_/X sky130_fd_sc_hd__buf_2
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22799_ _22799_/A VGND VGND VPWR VPWR _22799_/X sky130_fd_sc_hd__buf_2
XANTENNA__14039__A _12581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20983__B _20422_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15340_ _15328_/A _23992_/Q VGND VGND VPWR VPWR _15341_/C sky130_fd_sc_hd__or2_4
X_12552_ _12514_/A _12657_/B VGND VGND VPWR VPWR _12553_/C sky130_fd_sc_hd__or2_4
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21685__A2 _21684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22882__A1 _16016_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15271_ _12453_/A _15343_/B VGND VGND VPWR VPWR _15271_/X sky130_fd_sc_hd__or2_4
XANTENNA__13878__A _14377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12782__A _12800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24469_ _23126_/CLK _18778_/X HRESETn VGND VGND VPWR VPWR _24469_/Q sky130_fd_sc_hd__dfrtp_4
X_12483_ _13964_/A VGND VGND VPWR VPWR _12484_/A sky130_fd_sc_hd__buf_2
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ _24160_/Q _17010_/B VGND VGND VPWR VPWR _17011_/A sky130_fd_sc_hd__and2_4
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ _11780_/A _14213_/X _14221_/X VGND VGND VPWR VPWR _14222_/X sky130_fd_sc_hd__and3_4
XANTENNA__21437__A2 _21434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13597__B _13702_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22634__B2 _22598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19565__A _19848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14153_ _14171_/A VGND VGND VPWR VPWR _14272_/A sky130_fd_sc_hd__buf_2
XFILLER_164_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13104_ _13088_/A _13028_/B VGND VGND VPWR VPWR _13104_/X sky130_fd_sc_hd__or2_4
X_18961_ _18960_/X VGND VGND VPWR VPWR _20192_/A sky130_fd_sc_hd__inv_2
X_14084_ _11666_/X _14084_/B _14084_/C VGND VGND VPWR VPWR _14084_/X sky130_fd_sc_hd__and3_4
X_13035_ _12568_/A _13035_/B VGND VGND VPWR VPWR _13037_/B sky130_fd_sc_hd__or2_4
X_17912_ _17912_/A VGND VGND VPWR VPWR _18406_/A sky130_fd_sc_hd__buf_2
XFILLER_156_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18892_ _18891_/X VGND VGND VPWR VPWR _18893_/A sky130_fd_sc_hd__buf_2
XANTENNA__14502__A _14510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23753__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17843_ _17825_/A _17841_/X _17836_/X _17842_/X VGND VGND VPWR VPWR _17843_/X sky130_fd_sc_hd__o22a_4
XFILLER_152_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17774_ _17697_/A _17697_/B _18301_/A _17773_/X VGND VGND VPWR VPWR _17775_/D sky130_fd_sc_hd__or4_4
XANTENNA__12022__A _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14986_ _14170_/A _23509_/Q VGND VGND VPWR VPWR _14986_/X sky130_fd_sc_hd__or2_4
XFILLER_94_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19513_ _19471_/X _19476_/X _19511_/Y _17037_/Y _19512_/X VGND VGND VPWR VPWR _19514_/A
+ sky130_fd_sc_hd__a32o_4
X_16725_ _16725_/A _16725_/B _16725_/C VGND VGND VPWR VPWR _16726_/C sky130_fd_sc_hd__and3_4
X_13937_ _13937_/A _24093_/Q VGND VGND VPWR VPWR _13938_/C sky130_fd_sc_hd__or2_4
XFILLER_170_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11861__A _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19444_ _19480_/A VGND VGND VPWR VPWR _19445_/A sky130_fd_sc_hd__buf_2
X_16656_ _16656_/A _16654_/X _16655_/X VGND VGND VPWR VPWR _16656_/X sky130_fd_sc_hd__and3_4
X_13868_ _13868_/A VGND VGND VPWR VPWR _13877_/A sky130_fd_sc_hd__buf_2
X_12819_ _12833_/A _12819_/B VGND VGND VPWR VPWR _12821_/B sky130_fd_sc_hd__or2_4
XANTENNA__11580__B IRQ[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15607_ _15642_/A _15607_/B VGND VGND VPWR VPWR _15607_/X sky130_fd_sc_hd__or2_4
X_19375_ _19372_/X _18704_/X _19372_/X _24248_/Q VGND VGND VPWR VPWR _19375_/X sky130_fd_sc_hd__a2bb2o_4
X_16587_ _16554_/X _24114_/Q VGND VGND VPWR VPWR _16588_/C sky130_fd_sc_hd__or2_4
X_13799_ _13799_/A VGND VGND VPWR VPWR _15393_/A sky130_fd_sc_hd__buf_2
XFILLER_76_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24259__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18326_ _18187_/X _18309_/X _18219_/X _18325_/X VGND VGND VPWR VPWR _18326_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21676__A2 _21670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15538_ _14418_/X _15536_/X _15537_/X VGND VGND VPWR VPWR _15538_/X sky130_fd_sc_hd__and3_4
XANTENNA__22873__A1 _12320_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18363__B _17906_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13788__A _13788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15469_ _12576_/A _15461_/X _15468_/X VGND VGND VPWR VPWR _15485_/B sky130_fd_sc_hd__and3_4
X_18257_ _18037_/X _17460_/B VGND VGND VPWR VPWR _18257_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16164__A _13408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12692__A _12571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17208_ _12982_/X _17197_/X _17162_/Y _17198_/X VGND VGND VPWR VPWR _17208_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21428__A2 _21427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18188_ _17703_/A _16991_/B _18148_/C VGND VGND VPWR VPWR _23030_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__22625__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17139_ _16085_/X VGND VGND VPWR VPWR _17139_/X sky130_fd_sc_hd__buf_2
XFILLER_144_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20150_ _20150_/A _20149_/X VGND VGND VPWR VPWR _20150_/X sky130_fd_sc_hd__or2_4
XFILLER_104_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17707__B _17381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22389__B1 _23296_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20081_ _18551_/X _20079_/X _20080_/Y _20066_/X VGND VGND VPWR VPWR _20081_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20939__A1 _20894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14412__A _15517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20939__B2 _20861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15227__B _15227_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24370__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14131__B _23455_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13028__A _12510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23840_ _23744_/CLK _23840_/D VGND VGND VPWR VPWR _23840_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21245__A _21269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23771_ _23675_/CLK _21588_/X VGND VGND VPWR VPWR _23771_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12867__A _12867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20983_ _20867_/A _20422_/B VGND VGND VPWR VPWR _20983_/X sky130_fd_sc_hd__or2_4
XANTENNA__21364__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22722_ _22722_/A VGND VGND VPWR VPWR _22722_/X sky130_fd_sc_hd__buf_2
XPHY_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22653_ _22428_/X _22651_/X _16139_/B _22648_/X VGND VGND VPWR VPWR _22653_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21116__B2 _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21604_ _22687_/B VGND VGND VPWR VPWR _21656_/B sky130_fd_sc_hd__buf_2
XANTENNA__22864__A1 _17453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22584_ _22482_/X _22579_/X _23190_/Q _22548_/A VGND VGND VPWR VPWR _23190_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24323_ _24292_/CLK _19196_/X HRESETn VGND VGND VPWR VPWR _19144_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21535_ _21534_/X _21530_/X _23793_/Q _21525_/X VGND VGND VPWR VPWR _21535_/X sky130_fd_sc_hd__o22a_4
XFILLER_90_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24254_ _24248_/CLK _19367_/X HRESETn VGND VGND VPWR VPWR _20814_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22616__B2 _22612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21466_ _21311_/X _21462_/X _15227_/B _21431_/A VGND VGND VPWR VPWR _23831_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_6_7_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23205_ _23750_/CLK _23205_/D VGND VGND VPWR VPWR _13500_/B sky130_fd_sc_hd__dfxtp_4
X_20417_ _20302_/X _20416_/X _16294_/B _20396_/X VGND VGND VPWR VPWR _24111_/D sky130_fd_sc_hd__o22a_4
X_24185_ _23383_/CLK _24185_/D HRESETn VGND VGND VPWR VPWR _11595_/A sky130_fd_sc_hd__dfrtp_4
X_21397_ _21278_/X _21391_/X _13480_/B _21395_/X VGND VGND VPWR VPWR _21397_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12107__A _12001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16802__A _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23136_ _23617_/CLK _22671_/X VGND VGND VPWR VPWR _23136_/Q sky130_fd_sc_hd__dfxtp_4
X_20348_ _20347_/X VGND VGND VPWR VPWR _20349_/A sky130_fd_sc_hd__buf_2
XFILLER_108_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11946__A _16742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15418__A _11878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23067_ _23086_/A _23067_/B VGND VGND VPWR VPWR HADDR[28] sky130_fd_sc_hd__nor2_4
XANTENNA__14322__A _12198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20279_ _18784_/B _20279_/B VGND VGND VPWR VPWR _20493_/A sky130_fd_sc_hd__or2_4
XFILLER_88_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22018_ _21850_/X _22017_/X _15658_/B _22014_/X VGND VGND VPWR VPWR _22018_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11665__B _12410_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14840_ _14840_/A _14840_/B _14839_/X VGND VGND VPWR VPWR _14841_/C sky130_fd_sc_hd__or3_4
XFILLER_84_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15282__A1 _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21155__A _21155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14771_ _14771_/A VGND VGND VPWR VPWR _15112_/A sky130_fd_sc_hd__buf_2
X_23969_ _23303_/CLK _23969_/D VGND VGND VPWR VPWR _23969_/Q sky130_fd_sc_hd__dfxtp_4
X_11983_ _11868_/X _11927_/X _11948_/X _11964_/X _11982_/X VGND VGND VPWR VPWR _11983_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12777__A _12604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11681__A _11681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23156__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16510_ _16210_/A _16510_/B _16510_/C VGND VGND VPWR VPWR _16511_/C sky130_fd_sc_hd__and3_4
X_13722_ _13751_/A _13722_/B VGND VGND VPWR VPWR _13722_/X sky130_fd_sc_hd__or2_4
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15153__A _15281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24401__CLK _23281_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17490_ _17490_/A _17490_/B _17490_/C _17490_/D VGND VGND VPWR VPWR _17528_/A sky130_fd_sc_hd__or4_4
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16441_ _16129_/A _16441_/B _16440_/X VGND VGND VPWR VPWR _16441_/X sky130_fd_sc_hd__or3_4
XFILLER_147_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13653_ _15402_/A _13750_/B VGND VGND VPWR VPWR _13653_/X sky130_fd_sc_hd__or2_4
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21107__B2 _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22304__B1 _15458_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14992__A _14988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18464__A _18411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12604_ _12604_/A VGND VGND VPWR VPWR _12650_/A sky130_fd_sc_hd__buf_2
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _16342_/A _16294_/B VGND VGND VPWR VPWR _16372_/X sky130_fd_sc_hd__or2_4
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19160_ _24339_/Q _19160_/B VGND VGND VPWR VPWR _19160_/X sky130_fd_sc_hd__and2_4
XFILLER_9_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22855__A1 _13342_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13584_ _13485_/X _13583_/X _13570_/Y VGND VGND VPWR VPWR _16831_/B sky130_fd_sc_hd__a21o_4
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18111_ _18111_/A _18148_/B _18111_/C VGND VGND VPWR VPWR _18111_/X sky130_fd_sc_hd__and3_4
X_15323_ _15319_/A _23768_/Q VGND VGND VPWR VPWR _15324_/C sky130_fd_sc_hd__or2_4
X_12535_ _12864_/A _23979_/Q VGND VGND VPWR VPWR _12536_/C sky130_fd_sc_hd__or2_4
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19091_ _19074_/X _19089_/X _19090_/Y _19079_/X VGND VGND VPWR VPWR _19091_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20330__A2 _20847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18042_ _17095_/X _18038_/Y _18042_/C _18042_/D VGND VGND VPWR VPWR _18043_/A sky130_fd_sc_hd__or4_4
X_15254_ _14138_/A _23512_/Q VGND VGND VPWR VPWR _15255_/C sky130_fd_sc_hd__or2_4
XANTENNA__22607__B2 _22605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12466_ _12466_/A VGND VGND VPWR VPWR _12467_/A sky130_fd_sc_hd__buf_2
X_14205_ _14200_/A _23583_/Q VGND VGND VPWR VPWR _14205_/X sky130_fd_sc_hd__or2_4
XANTENNA__14216__B _23999_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12020__A1 _11858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15185_ _13951_/X _11627_/A _15154_/X _11604_/A _15184_/X VGND VGND VPWR VPWR _15185_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22083__A2 _22081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12397_ _11682_/A VGND VGND VPWR VPWR _13564_/A sky130_fd_sc_hd__buf_2
XANTENNA__12017__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12020__B2 _12019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14136_ _15281_/A VGND VGND VPWR VPWR _14302_/A sky130_fd_sc_hd__buf_2
XFILLER_158_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21830__A2 _21827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19993_ _19993_/A VGND VGND VPWR VPWR _19993_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11856__A _11856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18944_ _11544_/D VGND VGND VPWR VPWR _18949_/A sky130_fd_sc_hd__inv_2
X_14067_ _14075_/A _23104_/Q VGND VGND VPWR VPWR _14069_/B sky130_fd_sc_hd__or2_4
XANTENNA__14232__A _14635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13018_ _12878_/A _13018_/B VGND VGND VPWR VPWR _13018_/X sky130_fd_sc_hd__or2_4
XANTENNA__11575__B IRQ[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18875_ _13945_/X _18870_/X _20825_/A _18871_/X VGND VGND VPWR VPWR _24413_/D sky130_fd_sc_hd__o22a_4
XFILLER_121_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17826_ _17233_/X _17141_/X _17231_/X _17143_/X VGND VGND VPWR VPWR _17826_/X sky130_fd_sc_hd__o22a_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17757_ _17746_/X _17747_/X _17756_/X VGND VGND VPWR VPWR _17757_/X sky130_fd_sc_hd__or3_4
XANTENNA__17262__B _17251_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12687__A _12687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_13_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14969_ _14976_/A _23702_/Q VGND VGND VPWR VPWR _14971_/B sky130_fd_sc_hd__or2_4
XANTENNA__21346__B2 _21345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16159__A _16159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24081__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16708_ _12041_/A _23569_/Q VGND VGND VPWR VPWR _16709_/C sky130_fd_sc_hd__or2_4
XANTENNA__21897__A2 _21895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18211__B2 _18210_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17688_ _17688_/A _17520_/X VGND VGND VPWR VPWR _17688_/X sky130_fd_sc_hd__or2_4
XANTENNA__15998__A _13474_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19427_ _19425_/X _18633_/X _19425_/X _24219_/Q VGND VGND VPWR VPWR _24219_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16639_ _16639_/A VGND VGND VPWR VPWR _16677_/A sky130_fd_sc_hd__buf_2
X_19358_ _19372_/A VGND VGND VPWR VPWR _19358_/X sky130_fd_sc_hd__buf_2
XANTENNA__21649__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18309_ _18249_/X _23009_/B _18251_/Y VGND VGND VPWR VPWR _18309_/X sky130_fd_sc_hd__o21a_4
X_19289_ _19289_/A VGND VGND VPWR VPWR _19289_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21320_ _21184_/A _21420_/B _21320_/C _21236_/D VGND VGND VPWR VPWR _21320_/X sky130_fd_sc_hd__or4_4
X_21251_ _21821_/A VGND VGND VPWR VPWR _21251_/X sky130_fd_sc_hd__buf_2
XFILLER_144_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21282__B1 _23940_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20202_ _24470_/Q VGND VGND VPWR VPWR _20202_/Y sky130_fd_sc_hd__inv_2
X_21182_ _21024_/X _21155_/A _23989_/Q _21137_/X VGND VGND VPWR VPWR _23989_/D sky130_fd_sc_hd__o22a_4
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20133_ _11549_/A VGND VGND VPWR VPWR _20133_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20064_ _18670_/A VGND VGND VPWR VPWR _20064_/X sky130_fd_sc_hd__buf_2
XFILLER_86_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13981__A _13981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17453__A _12914_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23823_ _23119_/CLK _23823_/D VGND VGND VPWR VPWR _16301_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21337__B2 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23754_ _23467_/CLK _21626_/X VGND VGND VPWR VPWR _23754_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ _20965_/Y _20873_/X _19773_/X _20697_/X VGND VGND VPWR VPWR _20966_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _22705_/A VGND VGND VPWR VPWR _22705_/X sky130_fd_sc_hd__buf_2
XPHY_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13205__B _23783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23685_ _23557_/CLK _23685_/D VGND VGND VPWR VPWR _23685_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _21007_/A _20339_/B VGND VGND VPWR VPWR _20897_/X sky130_fd_sc_hd__or2_4
XANTENNA__17961__B1 _17653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15701__A _13303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22636_ _11824_/B VGND VGND VPWR VPWR _22636_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_33_0_HCLK clkbuf_6_16_0_HCLK/X VGND VGND VPWR VPWR _23764_/CLK sky130_fd_sc_hd__clkbuf_1
X_22567_ _22452_/X _22565_/X _15796_/B _22562_/X VGND VGND VPWR VPWR _22567_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14317__A _14292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13221__A _12362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12320_ _12320_/A VGND VGND VPWR VPWR _12320_/Y sky130_fd_sc_hd__inv_2
X_24306_ _24306_/CLK _19262_/X HRESETn VGND VGND VPWR VPWR _24306_/Q sky130_fd_sc_hd__dfrtp_4
X_21518_ _21313_/X _21513_/X _14967_/B _21482_/A VGND VGND VPWR VPWR _23798_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_7_96_0_HCLK clkbuf_6_48_0_HCLK/X VGND VGND VPWR VPWR _23617_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_139_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22498_ _22498_/A VGND VGND VPWR VPWR _22498_/X sky130_fd_sc_hd__buf_2
XFILLER_154_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12251_ _12251_/A VGND VGND VPWR VPWR _13677_/A sky130_fd_sc_hd__buf_2
X_24237_ _24495_/CLK _24237_/D HRESETn VGND VGND VPWR VPWR _24237_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22065__A2 _22060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21449_ _21280_/X _21448_/X _15760_/B _21445_/X VGND VGND VPWR VPWR _21449_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24168_ _23991_/CLK _24168_/D HRESETn VGND VGND VPWR VPWR _24168_/Q sky130_fd_sc_hd__dfrtp_4
X_12182_ _12111_/X _12182_/B VGND VGND VPWR VPWR _12183_/A sky130_fd_sc_hd__or2_4
XFILLER_134_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11676__A _12641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23119_ _23119_/CLK _22700_/X VGND VGND VPWR VPWR _16300_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15148__A _14171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_122_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24099_ _23939_/CLK _20694_/X VGND VGND VPWR VPWR _15834_/B sky130_fd_sc_hd__dfxtp_4
X_16990_ _16954_/Y _18189_/A VGND VGND VPWR VPWR _16991_/B sky130_fd_sc_hd__or2_4
XFILLER_1_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14052__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21025__B1 _24085_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15941_ _15936_/X _15941_/B _15940_/X VGND VGND VPWR VPWR _15941_/X sky130_fd_sc_hd__and3_4
XFILLER_118_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14987__A _14897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21576__B2 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18459__A _18406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13891__A _14507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18660_ _17741_/A _16973_/X _24136_/Q _18661_/A VGND VGND VPWR VPWR _22931_/B sky130_fd_sc_hd__o22a_4
X_15872_ _13539_/A _15803_/B VGND VGND VPWR VPWR _15872_/X sky130_fd_sc_hd__or2_4
XFILLER_77_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17611_ _17401_/X VGND VGND VPWR VPWR _18587_/B sky130_fd_sc_hd__inv_2
XFILLER_63_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14823_ _14823_/A _23417_/Q VGND VGND VPWR VPWR _14824_/C sky130_fd_sc_hd__or2_4
XFILLER_91_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18591_ _18477_/X _18580_/X _18504_/X _18590_/X VGND VGND VPWR VPWR _18591_/X sky130_fd_sc_hd__o22a_4
XFILLER_76_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21328__B2 _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17542_ _17490_/D _17540_/X _17541_/Y VGND VGND VPWR VPWR _17542_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12300__A _12300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11966_ _13981_/A VGND VGND VPWR VPWR _11967_/A sky130_fd_sc_hd__buf_2
X_14754_ _12294_/A _14754_/B VGND VGND VPWR VPWR _14754_/X sky130_fd_sc_hd__or2_4
XFILLER_72_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21613__A _21620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19941__B2 _20917_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13705_ _13705_/A VGND VGND VPWR VPWR _13706_/A sky130_fd_sc_hd__buf_2
X_17473_ _17473_/A VGND VGND VPWR VPWR _17473_/Y sky130_fd_sc_hd__inv_2
X_14685_ _14685_/A _14683_/X _14685_/C VGND VGND VPWR VPWR _14685_/X sky130_fd_sc_hd__and3_4
X_11897_ _14110_/A VGND VGND VPWR VPWR _11898_/A sky130_fd_sc_hd__buf_2
XFILLER_44_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19212_ _19136_/A _19213_/A _19211_/Y VGND VGND VPWR VPWR _19212_/X sky130_fd_sc_hd__o21a_4
X_16424_ _16402_/X _16424_/B VGND VGND VPWR VPWR _16424_/X sky130_fd_sc_hd__or2_4
X_13636_ _13675_/A _23326_/Q VGND VGND VPWR VPWR _13636_/X sky130_fd_sc_hd__or2_4
XFILLER_73_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19143_ _24322_/Q _19142_/X VGND VGND VPWR VPWR _19143_/X sky130_fd_sc_hd__and2_4
XFILLER_160_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16355_ _16195_/A _16287_/B VGND VGND VPWR VPWR _16355_/X sky130_fd_sc_hd__or2_4
X_13567_ _13566_/X VGND VGND VPWR VPWR _13567_/X sky130_fd_sc_hd__buf_2
XANTENNA__21500__B2 _21496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13131__A _12273_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12518_ _12487_/A _12619_/B VGND VGND VPWR VPWR _12518_/X sky130_fd_sc_hd__or2_4
X_15306_ _14897_/X _15306_/B _15305_/X VGND VGND VPWR VPWR _15306_/X sky130_fd_sc_hd__and3_4
X_16286_ _16282_/A _16286_/B VGND VGND VPWR VPWR _16286_/X sky130_fd_sc_hd__or2_4
XFILLER_121_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19074_ _19016_/A VGND VGND VPWR VPWR _19074_/X sky130_fd_sc_hd__buf_2
X_13498_ _13528_/A _13491_/X _13497_/X VGND VGND VPWR VPWR _13498_/X sky130_fd_sc_hd__or3_4
XFILLER_145_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22444__A _20612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18025_ _17660_/A _18024_/X VGND VGND VPWR VPWR _18025_/Y sky130_fd_sc_hd__nand2_4
X_12449_ _12863_/A _23371_/Q VGND VGND VPWR VPWR _12458_/B sky130_fd_sc_hd__or2_4
XANTENNA__22056__A2 _22053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15237_ _14677_/A _15179_/B VGND VGND VPWR VPWR _15239_/B sky130_fd_sc_hd__or2_4
XANTENNA__17538__A _12980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12970__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15168_ _13589_/A _15168_/B _15168_/C VGND VGND VPWR VPWR _15168_/X sky130_fd_sc_hd__or3_4
XFILLER_119_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14119_ _14155_/A VGND VGND VPWR VPWR _14131_/A sky130_fd_sc_hd__buf_2
XANTENNA__15058__A _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19976_ _16943_/X _19386_/X _17014_/X _19975_/X VGND VGND VPWR VPWR _19976_/X sky130_fd_sc_hd__o22a_4
X_15099_ _14682_/A _15091_/X _15098_/X VGND VGND VPWR VPWR _15099_/X sky130_fd_sc_hd__and3_4
XFILLER_87_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18927_ _18896_/A VGND VGND VPWR VPWR _18927_/X sky130_fd_sc_hd__buf_2
XANTENNA__21567__B2 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17273__A _14334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18858_ _17156_/A _18856_/X _24426_/Q _18857_/X VGND VGND VPWR VPWR _24426_/D sky130_fd_sc_hd__o22a_4
XFILLER_68_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17809_ _17809_/A VGND VGND VPWR VPWR _17809_/X sky130_fd_sc_hd__buf_2
X_18789_ _18789_/A VGND VGND VPWR VPWR _18790_/A sky130_fd_sc_hd__buf_2
X_20820_ _20772_/X _20819_/X _24094_/Q _20746_/X VGND VGND VPWR VPWR _20820_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12210__A _12687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18735__A2 _17246_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21523__A _21523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20751_ _20845_/A _20751_/B _20750_/X VGND VGND VPWR VPWR _20751_/X sky130_fd_sc_hd__and3_4
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23470_ _23501_/CLK _22112_/X VGND VGND VPWR VPWR _23470_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20682_ _20490_/X _20681_/Y _19240_/A _20584_/X VGND VGND VPWR VPWR _20682_/X sky130_fd_sc_hd__o22a_4
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22421_ _22421_/A VGND VGND VPWR VPWR _22421_/X sky130_fd_sc_hd__buf_2
XFILLER_149_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22295__A2 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13041__A _12492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22352_ _14867_/B VGND VGND VPWR VPWR _22352_/X sky130_fd_sc_hd__buf_2
XANTENNA__17171__A1 _17170_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21303_ _21302_/X _21293_/X _14499_/B _21300_/X VGND VGND VPWR VPWR _21303_/X sky130_fd_sc_hd__o22a_4
XFILLER_163_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22047__A2 _22046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17448__A _15916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22283_ _22103_/X _22280_/X _16756_/B _22277_/X VGND VGND VPWR VPWR _22283_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20058__A1 _20040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24022_ _23416_/CLK _21130_/X VGND VGND VPWR VPWR _14859_/B sky130_fd_sc_hd__dfxtp_4
X_21234_ _21234_/A _21234_/B VGND VGND VPWR VPWR _22537_/D sky130_fd_sc_hd__or2_4
XFILLER_137_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21165_ _20719_/X _21162_/X _15478_/B _21159_/X VGND VGND VPWR VPWR _24002_/D sky130_fd_sc_hd__o22a_4
XFILLER_46_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20116_ _20150_/A _20114_/X _20115_/Y _19959_/A VGND VGND VPWR VPWR _20116_/X sky130_fd_sc_hd__o22a_4
X_21096_ _20416_/X _21090_/X _16259_/B _21094_/X VGND VGND VPWR VPWR _21096_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18423__A1 _18413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20047_ _20047_/A VGND VGND VPWR VPWR _20047_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14600__A _13658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11820_ _11832_/A _21805_/A VGND VGND VPWR VPWR _11822_/B sky130_fd_sc_hd__or2_4
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23806_ _23101_/CLK _21508_/X VGND VGND VPWR VPWR _13766_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23964__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12120__A _16080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _21817_/X _21996_/X _23538_/Q _21993_/X VGND VGND VPWR VPWR _23538_/D sky130_fd_sc_hd__o22a_4
XFILLER_61_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22529__A _22489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11751_ _15330_/A VGND VGND VPWR VPWR _11752_/A sky130_fd_sc_hd__buf_2
X_23737_ _23391_/CLK _23737_/D VGND VGND VPWR VPWR _14780_/B sky130_fd_sc_hd__dfxtp_4
X_20949_ _20425_/A _20948_/X _24280_/Q _20758_/X VGND VGND VPWR VPWR _20949_/X sky130_fd_sc_hd__o22a_4
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21730__B2 _21724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _12512_/A _14470_/B VGND VGND VPWR VPWR _14470_/X sky130_fd_sc_hd__or2_4
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11682_/A VGND VGND VPWR VPWR _13123_/A sky130_fd_sc_hd__buf_2
X_23668_ _23668_/CLK _21761_/X VGND VGND VPWR VPWR _23668_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13421_ _13330_/A _13419_/X _13421_/C VGND VGND VPWR VPWR _13421_/X sky130_fd_sc_hd__and3_4
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22619_ _22605_/A VGND VGND VPWR VPWR _22619_/X sky130_fd_sc_hd__buf_2
XANTENNA__22286__A2 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23599_ _23983_/CLK _23599_/D VGND VGND VPWR VPWR _16271_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14047__A _11736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16140_ _16109_/A _16140_/B VGND VGND VPWR VPWR _16141_/C sky130_fd_sc_hd__or2_4
XFILLER_128_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20297__A1 _20358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13352_ _13370_/A VGND VGND VPWR VPWR _13375_/A sky130_fd_sc_hd__buf_2
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20297__B2 _20334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12303_ _13332_/A _12303_/B VGND VGND VPWR VPWR _12303_/X sky130_fd_sc_hd__or2_4
XFILLER_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16071_ _16035_/A _16071_/B _16070_/X VGND VGND VPWR VPWR _16075_/B sky130_fd_sc_hd__and3_4
XFILLER_143_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13886__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13283_ _12559_/A _13283_/B VGND VGND VPWR VPWR _13285_/B sky130_fd_sc_hd__or2_4
XANTENNA__12790__A _12801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23079__B _23079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20049__A1 _20040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15022_ _15022_/A _15018_/X _15022_/C VGND VGND VPWR VPWR _15022_/X sky130_fd_sc_hd__or3_4
XFILLER_107_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12234_ _12250_/A VGND VGND VPWR VPWR _13687_/A sky130_fd_sc_hd__buf_2
XFILLER_30_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21797__B2 _21795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19830_ _19642_/Y _19808_/A VGND VGND VPWR VPWR _19830_/X sky130_fd_sc_hd__or2_4
XFILLER_155_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12165_ _12129_/A _12163_/X _12165_/C VGND VGND VPWR VPWR _12169_/B sky130_fd_sc_hd__and3_4
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19761_ _19849_/A VGND VGND VPWR VPWR _19890_/A sky130_fd_sc_hd__buf_2
XANTENNA__21608__A _21608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16973_ _17748_/A _17749_/A _17743_/A VGND VGND VPWR VPWR _16973_/X sky130_fd_sc_hd__or3_4
X_12096_ _12093_/X _12094_/X _12095_/X VGND VGND VPWR VPWR _12101_/B sky130_fd_sc_hd__and3_4
XFILLER_89_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22746__B1 HREADY VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18712_ _17920_/X _17885_/B _17944_/X _18711_/X VGND VGND VPWR VPWR _18712_/X sky130_fd_sc_hd__a211o_4
X_15924_ _15923_/X VGND VGND VPWR VPWR _16842_/B sky130_fd_sc_hd__inv_2
XANTENNA__15606__A _15606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19692_ _19507_/A VGND VGND VPWR VPWR _19849_/A sky130_fd_sc_hd__buf_2
XANTENNA__22210__A2 _22208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14510__A _14510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18643_ _17793_/X _18635_/X _18636_/Y _18638_/X _18642_/Y VGND VGND VPWR VPWR _18643_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15855_ _13514_/A _15855_/B _15855_/C VGND VGND VPWR VPWR _15856_/C sky130_fd_sc_hd__and3_4
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13126__A _13049_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14806_ _14691_/A _14723_/B VGND VGND VPWR VPWR _14806_/X sky130_fd_sc_hd__or2_4
XFILLER_149_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18574_ _18399_/X VGND VGND VPWR VPWR _18574_/X sky130_fd_sc_hd__buf_2
XANTENNA__12030__A _16595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15786_ _15783_/X VGND VGND VPWR VPWR _15786_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12998_ _12905_/A _24040_/Q VGND VGND VPWR VPWR _13000_/B sky130_fd_sc_hd__or2_4
XFILLER_17_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17525_ _17523_/Y _17524_/X VGND VGND VPWR VPWR _17605_/D sky130_fd_sc_hd__or2_4
XFILLER_73_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14737_ _12484_/A _14737_/B VGND VGND VPWR VPWR _14737_/X sky130_fd_sc_hd__or2_4
XANTENNA__12965__A _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11949_ _16145_/A VGND VGND VPWR VPWR _12108_/A sky130_fd_sc_hd__buf_2
XANTENNA__21721__B2 _21717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15341__A _13695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17456_ _17455_/X VGND VGND VPWR VPWR _17456_/Y sky130_fd_sc_hd__inv_2
X_14668_ _14653_/A _23610_/Q VGND VGND VPWR VPWR _14668_/X sky130_fd_sc_hd__or2_4
XFILLER_60_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16407_ _15998_/X _16403_/X _16406_/X VGND VGND VPWR VPWR _16407_/X sky130_fd_sc_hd__and3_4
XANTENNA__15060__B _23765_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13619_ _15423_/A _13722_/B VGND VGND VPWR VPWR _13619_/X sky130_fd_sc_hd__or2_4
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17387_ _17387_/A VGND VGND VPWR VPWR _17387_/Y sky130_fd_sc_hd__inv_2
X_14599_ _13657_/A _14597_/X _14598_/X VGND VGND VPWR VPWR _14599_/X sky130_fd_sc_hd__and3_4
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19126_ _19126_/A VGND VGND VPWR VPWR _19126_/Y sky130_fd_sc_hd__inv_2
X_16338_ _16316_/A _16338_/B VGND VGND VPWR VPWR _16338_/X sky130_fd_sc_hd__or2_4
XFILLER_125_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13796__A _14304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19057_ _19046_/X _19055_/X _19056_/Y _19049_/X VGND VGND VPWR VPWR _19057_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17268__A _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22029__A2 _22024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16269_ _15971_/A _16265_/X _16268_/X VGND VGND VPWR VPWR _16269_/X sky130_fd_sc_hd__or3_4
XANTENNA__16172__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18008_ _18008_/A VGND VGND VPWR VPWR _18176_/A sky130_fd_sc_hd__buf_2
XFILLER_160_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14911__B1 _11603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12205__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16900__A _17060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19959_ _19959_/A VGND VGND VPWR VPWR _20150_/A sky130_fd_sc_hd__inv_2
XFILLER_113_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15516__A _12978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22970_ _22969_/X VGND VGND VPWR VPWR HADDR[11] sky130_fd_sc_hd__inv_2
XFILLER_132_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21921_ _21857_/X _21916_/X _15602_/B _21920_/X VGND VGND VPWR VPWR _23585_/D sky130_fd_sc_hd__o22a_4
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15235__B _15177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13036__A _12569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21852_ _21850_/X _21851_/X _15755_/B _21846_/X VGND VGND VPWR VPWR _23620_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19905__A1 _19469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23217__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20803_ HRDATA[9] _20843_/B VGND VGND VPWR VPWR _20803_/X sky130_fd_sc_hd__or2_4
XFILLER_82_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21783_ _21563_/X _21777_/X _23653_/Q _21781_/X VGND VGND VPWR VPWR _21783_/X sky130_fd_sc_hd__o22a_4
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24119__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12875__A _12875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23522_ _23587_/CLK _22020_/X VGND VGND VPWR VPWR _15455_/B sky130_fd_sc_hd__dfxtp_4
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15251__A _15251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20734_ _20726_/X _20733_/Y _24289_/Q _20584_/X VGND VGND VPWR VPWR _20734_/X sky130_fd_sc_hd__o22a_4
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23453_ _23582_/CLK _23453_/D VGND VGND VPWR VPWR _13901_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_149_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20665_ _17077_/A VGND VGND VPWR VPWR _20665_/X sky130_fd_sc_hd__buf_2
XANTENNA__22268__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18562__A _18562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22404_ _11718_/B VGND VGND VPWR VPWR _22404_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23384_ _23290_/CLK _23384_/D VGND VGND VPWR VPWR _23384_/Q sky130_fd_sc_hd__dfxtp_4
X_20596_ _20596_/A VGND VGND VPWR VPWR _20596_/X sky130_fd_sc_hd__buf_2
XFILLER_149_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22335_ _13148_/B VGND VGND VPWR VPWR _22335_/X sky130_fd_sc_hd__buf_2
XANTENNA__16082__A _11759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22266_ _22158_/X _22265_/X _23386_/Q _22262_/X VGND VGND VPWR VPWR _22266_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14314__B _14391_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22812__A _17273_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24005_ _23493_/CLK _24005_/D VGND VGND VPWR VPWR _24005_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21779__B2 _21774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21217_ _20745_/X _21212_/X _23969_/Q _21216_/X VGND VGND VPWR VPWR _23969_/D sky130_fd_sc_hd__o22a_4
XFILLER_132_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22197_ _22127_/X _22194_/X _13241_/B _22191_/X VGND VGND VPWR VPWR _23431_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12115__A _16080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18644__B2 _18643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21148_ _21155_/A VGND VGND VPWR VPWR _21148_/X sky130_fd_sc_hd__buf_2
XFILLER_120_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17625__B _17346_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11954__A _11905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15426__A _14319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14330__A _11913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13970_ _13627_/A _22342_/A VGND VGND VPWR VPWR _13970_/X sky130_fd_sc_hd__or2_4
X_21079_ _21024_/X _21045_/A _24053_/Q _21042_/A VGND VGND VPWR VPWR _21079_/X sky130_fd_sc_hd__o22a_4
XFILLER_47_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20203__B2 _19951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12921_ _12659_/A _12917_/X _12921_/C VGND VGND VPWR VPWR _12921_/X sky130_fd_sc_hd__or3_4
XFILLER_19_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21951__B2 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15640_ _14335_/A _15636_/X _15639_/X VGND VGND VPWR VPWR _15640_/X sky130_fd_sc_hd__or3_4
X_12852_ _12852_/A VGND VGND VPWR VPWR _12884_/A sky130_fd_sc_hd__buf_2
X_11803_ _11742_/X VGND VGND VPWR VPWR _16647_/A sky130_fd_sc_hd__buf_2
XANTENNA__24142__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12783_ _13055_/A VGND VGND VPWR VPWR _12783_/X sky130_fd_sc_hd__buf_2
X_15571_ _12428_/A _15569_/X _15571_/C VGND VGND VPWR VPWR _15572_/C sky130_fd_sc_hd__and3_4
XANTENNA__12785__A _12801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21703__B2 _21667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15161__A _14277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17310_ _17307_/X _17310_/B VGND VGND VPWR VPWR _17310_/X sky130_fd_sc_hd__or2_4
X_14522_ _14522_/A _14518_/X _14522_/C VGND VGND VPWR VPWR _14522_/X sky130_fd_sc_hd__or3_4
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ _13717_/A VGND VGND VPWR VPWR _11735_/A sky130_fd_sc_hd__buf_2
XFILLER_159_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _18290_/A _17508_/X _17638_/Y VGND VGND VPWR VPWR _18290_/X sky130_fd_sc_hd__or3_4
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24347__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17229_/X _17237_/Y _17240_/X VGND VGND VPWR VPWR _17241_/X sky130_fd_sc_hd__o21a_4
X_14453_ _12455_/A _23963_/Q VGND VGND VPWR VPWR _14454_/C sky130_fd_sc_hd__or2_4
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11665_ _15616_/A _12410_/A _12955_/A _11665_/D VGND VGND VPWR VPWR _11665_/X sky130_fd_sc_hd__or4_4
XANTENNA__22259__A2 _22258_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24292__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _13378_/A _23718_/Q VGND VGND VPWR VPWR _13406_/B sky130_fd_sc_hd__or2_4
XFILLER_122_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _14522_/A _14379_/X _14383_/X VGND VGND VPWR VPWR _14384_/X sky130_fd_sc_hd__or3_4
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17172_ _13417_/X VGND VGND VPWR VPWR _17172_/X sky130_fd_sc_hd__buf_2
XFILLER_128_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11596_ _11596_/A VGND VGND VPWR VPWR _17017_/A sky130_fd_sc_hd__buf_2
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16123_ _16123_/A _16123_/B _16123_/C VGND VGND VPWR VPWR _16123_/X sky130_fd_sc_hd__and3_4
X_13335_ _11888_/A _23718_/Q VGND VGND VPWR VPWR _13335_/X sky130_fd_sc_hd__or2_4
XANTENNA__18883__A1 _15251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16054_ _16061_/A _16054_/B VGND VGND VPWR VPWR _16054_/X sky130_fd_sc_hd__or2_4
X_13266_ _13125_/X VGND VGND VPWR VPWR _13266_/X sky130_fd_sc_hd__buf_2
XANTENNA__22722__A _22722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12217_ _11895_/X VGND VGND VPWR VPWR _12218_/A sky130_fd_sc_hd__buf_2
X_15005_ _13985_/A _15005_/B _15005_/C VGND VGND VPWR VPWR _15005_/X sky130_fd_sc_hd__and3_4
XFILLER_124_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13197_ _13223_/A _13195_/X _13196_/X VGND VGND VPWR VPWR _13197_/X sky130_fd_sc_hd__and3_4
XANTENNA__22431__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20442__A1 _20418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19813_ _19644_/Y _19807_/Y _19767_/A _19812_/X VGND VGND VPWR VPWR _19813_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20442__B2 _20396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21338__A _21338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12148_ _16608_/A _23923_/Q VGND VGND VPWR VPWR _12148_/X sky130_fd_sc_hd__or2_4
XFILLER_111_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11864__A _11864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19744_ _19744_/A _19711_/A VGND VGND VPWR VPWR _19744_/X sky130_fd_sc_hd__or2_4
XANTENNA__15336__A _13704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16956_ _24150_/Q VGND VGND VPWR VPWR _16988_/A sky130_fd_sc_hd__inv_2
X_12079_ _16704_/A _23923_/Q VGND VGND VPWR VPWR _12081_/B sky130_fd_sc_hd__or2_4
XFILLER_38_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22195__B2 _22191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15907_ _13554_/A _15837_/B VGND VGND VPWR VPWR _15907_/X sky130_fd_sc_hd__or2_4
X_19675_ _19675_/A VGND VGND VPWR VPWR _19819_/A sky130_fd_sc_hd__buf_2
XFILLER_38_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12683__A1 _12574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16887_ _16858_/X _16884_/X _16885_/X _16887_/D VGND VGND VPWR VPWR _16887_/X sky130_fd_sc_hd__and4_4
XANTENNA__20896__B _20512_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18626_ _17758_/X _17739_/X _17758_/X _17739_/X VGND VGND VPWR VPWR _18626_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17551__A _17120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15838_ _12903_/A _15838_/B _15838_/C VGND VGND VPWR VPWR _15839_/C sky130_fd_sc_hd__and3_4
XFILLER_80_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22169__A _22169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21073__A _21033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18557_ _18557_/A _18557_/B VGND VGND VPWR VPWR _18557_/Y sky130_fd_sc_hd__nand2_4
XFILLER_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15769_ _12778_/X _15767_/X _15768_/X VGND VGND VPWR VPWR _15769_/X sky130_fd_sc_hd__and3_4
XANTENNA__24212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17508_ _18336_/B _17508_/B VGND VGND VPWR VPWR _17508_/X sky130_fd_sc_hd__or2_4
X_18488_ _18487_/X VGND VGND VPWR VPWR _18488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21170__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _17153_/Y _17439_/B VGND VGND VPWR VPWR _17439_/X sky130_fd_sc_hd__or2_4
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20450_ _20450_/A _20450_/B VGND VGND VPWR VPWR _20450_/X sky130_fd_sc_hd__or2_4
XANTENNA__17126__A1 _17339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19109_ _18957_/X VGND VGND VPWR VPWR _19109_/X sky130_fd_sc_hd__buf_2
X_20381_ _20251_/X _20380_/X _20235_/X VGND VGND VPWR VPWR _20381_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__18874__A1 _17153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22120_ _20530_/A VGND VGND VPWR VPWR _22120_/X sky130_fd_sc_hd__buf_2
XFILLER_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22051_ _21821_/X _22046_/X _16435_/B _22050_/X VGND VGND VPWR VPWR _23504_/D sky130_fd_sc_hd__o22a_4
XFILLER_133_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22422__A2 _22414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16630__A _16683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21002_ _24214_/Q _20895_/X _21001_/X VGND VGND VPWR VPWR _22482_/A sky130_fd_sc_hd__o21a_4
XFILLER_87_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17445__B _17445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20152__A _20200_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15246__A _14635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14150__A _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22186__B2 _22184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24165__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22953_ _22952_/X VGND VGND VPWR VPWR HADDR[8] sky130_fd_sc_hd__inv_2
XANTENNA__21933__B2 _21927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21904_ _21829_/X _21902_/X _16189_/B _21899_/X VGND VGND VPWR VPWR _21904_/X sky130_fd_sc_hd__o22a_4
X_22884_ _22884_/A VGND VGND VPWR VPWR _22897_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21835_ _21833_/X _21827_/X _12646_/B _21834_/X VGND VGND VPWR VPWR _23627_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16077__A _16049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21766_ _21534_/X _21763_/X _23665_/Q _21760_/X VGND VGND VPWR VPWR _23665_/D sky130_fd_sc_hd__o22a_4
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21161__A2 _21155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22807__A _17327_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23505_ _23761_/CLK _22049_/X VGND VGND VPWR VPWR _23505_/Q sky130_fd_sc_hd__dfxtp_4
X_20717_ _24226_/Q _20636_/X _20716_/Y VGND VGND VPWR VPWR _20718_/A sky130_fd_sc_hd__o21a_4
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24485_ _24127_/CLK _24485_/D HRESETn VGND VGND VPWR VPWR _24485_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21697_ _21587_/X _21691_/X _14534_/B _21695_/X VGND VGND VPWR VPWR _23707_/D sky130_fd_sc_hd__o22a_4
XFILLER_106_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23436_ _23404_/CLK _23436_/D VGND VGND VPWR VPWR _12393_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20648_ _20470_/X _20646_/X _24388_/Q _20647_/X VGND VGND VPWR VPWR _20648_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17117__A1 _15382_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20327__A _20264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16524__B _16521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11949__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23367_ _23303_/CLK _23367_/D VGND VGND VPWR VPWR _13199_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18865__A1 _13567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22661__A2 _22658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20579_ _20579_/A _20617_/B VGND VGND VPWR VPWR _20579_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__14325__A _14325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13120_ _12762_/A _23656_/Q VGND VGND VPWR VPWR _13120_/X sky130_fd_sc_hd__or2_4
XFILLER_124_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22318_ _22163_/X _22315_/X _23352_/Q _22312_/X VGND VGND VPWR VPWR _23352_/D sky130_fd_sc_hd__o22a_4
X_23298_ _23523_/CLK _23298_/D VGND VGND VPWR VPWR _15466_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_152_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13051_ _13051_/A VGND VGND VPWR VPWR _13103_/A sky130_fd_sc_hd__buf_2
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22249_ _22129_/X _22244_/X _23398_/Q _22248_/X VGND VGND VPWR VPWR _22249_/X sky130_fd_sc_hd__o22a_4
XFILLER_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19814__B1 _16672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12002_ _12105_/A _11841_/B VGND VGND VPWR VPWR _12006_/B sky130_fd_sc_hd__or2_4
XFILLER_133_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16810_ _16791_/A _23505_/Q VGND VGND VPWR VPWR _16810_/X sky130_fd_sc_hd__or2_4
XANTENNA__19851__A _19848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17790_ _18220_/A VGND VGND VPWR VPWR _18150_/A sky130_fd_sc_hd__buf_2
XANTENNA__14060__A _13705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16741_ _16741_/A _23121_/Q VGND VGND VPWR VPWR _16743_/B sky130_fd_sc_hd__or2_4
XFILLER_115_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13953_ _13953_/A _23520_/Q VGND VGND VPWR VPWR _13954_/C sky130_fd_sc_hd__or2_4
XANTENNA__14995__A _14171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21924__B2 _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12904_ _12904_/A _12904_/B _12903_/X VGND VGND VPWR VPWR _12904_/X sky130_fd_sc_hd__or3_4
X_19460_ _19442_/X VGND VGND VPWR VPWR _19461_/A sky130_fd_sc_hd__buf_2
X_16672_ _16672_/A _23730_/Q VGND VGND VPWR VPWR _16674_/B sky130_fd_sc_hd__or2_4
XFILLER_59_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13884_ _13884_/A _13807_/B VGND VGND VPWR VPWR _13886_/B sky130_fd_sc_hd__or2_4
X_18411_ _18411_/A _18411_/B VGND VGND VPWR VPWR _18411_/X sky130_fd_sc_hd__and2_4
X_15623_ _15642_/A _24065_/Q VGND VGND VPWR VPWR _15624_/C sky130_fd_sc_hd__or2_4
X_12835_ _13349_/A _12835_/B _12834_/X VGND VGND VPWR VPWR _12839_/B sky130_fd_sc_hd__and3_4
X_19391_ _19389_/X _17910_/X _19389_/X _24241_/Q VGND VGND VPWR VPWR _24241_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13404__A _13378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18342_ _17976_/X _17220_/X _17882_/X VGND VGND VPWR VPWR _18343_/B sky130_fd_sc_hd__o21ai_4
X_15554_ _12236_/A _15552_/X _15554_/C VGND VGND VPWR VPWR _15558_/B sky130_fd_sc_hd__and3_4
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _13058_/A VGND VGND VPWR VPWR _12766_/X sky130_fd_sc_hd__buf_2
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14219__B _23551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14505_ _14522_/A _14505_/B _14504_/X VGND VGND VPWR VPWR _14505_/X sky130_fd_sc_hd__or3_4
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _18187_/X _18254_/X _18219_/X _18272_/X VGND VGND VPWR VPWR _18273_/X sky130_fd_sc_hd__o22a_4
X_11717_ _16079_/A VGND VGND VPWR VPWR _11717_/X sky130_fd_sc_hd__buf_2
X_12697_ _12721_/A _12785_/B VGND VGND VPWR VPWR _12697_/X sky130_fd_sc_hd__or2_4
X_15485_ _13229_/A _15485_/B _15485_/C VGND VGND VPWR VPWR _15485_/X sky130_fd_sc_hd__or3_4
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16715__A _11941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17224_ _18265_/A VGND VGND VPWR VPWR _17224_/X sky130_fd_sc_hd__buf_2
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14436_ _12531_/A _14436_/B VGND VGND VPWR VPWR _14438_/B sky130_fd_sc_hd__or2_4
XFILLER_35_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11648_ _11643_/A _11590_/X VGND VGND VPWR VPWR _11648_/X sky130_fd_sc_hd__or2_4
XFILLER_30_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11859__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15119__B1 _15117_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17155_ _12842_/X VGND VGND VPWR VPWR _17156_/A sky130_fd_sc_hd__buf_2
XANTENNA__22652__A2 _22651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14367_ _14367_/A _23996_/Q VGND VGND VPWR VPWR _14367_/X sky130_fd_sc_hd__or2_4
X_11579_ _11576_/X _20142_/A VGND VGND VPWR VPWR _20119_/A sky130_fd_sc_hd__or2_4
X_16106_ _15969_/A _16178_/B VGND VGND VPWR VPWR _16107_/C sky130_fd_sc_hd__or2_4
XFILLER_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13318_ _13318_/A _13316_/X _13317_/X VGND VGND VPWR VPWR _13318_/X sky130_fd_sc_hd__and3_4
X_17086_ _17054_/B VGND VGND VPWR VPWR _17089_/A sky130_fd_sc_hd__inv_2
X_14298_ _13617_/A _14362_/B VGND VGND VPWR VPWR _14298_/X sky130_fd_sc_hd__or2_4
XFILLER_143_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22452__A _20692_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16037_ _16187_/A _16026_/X _16037_/C VGND VGND VPWR VPWR _16053_/B sky130_fd_sc_hd__and3_4
X_13249_ _13256_/A _23879_/Q VGND VGND VPWR VPWR _13250_/C sky130_fd_sc_hd__or2_4
XFILLER_131_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19805__B1 _16659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15066__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17988_ _17823_/X VGND VGND VPWR VPWR _17988_/X sky130_fd_sc_hd__buf_2
XANTENNA__24464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22168__B2 _22106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19727_ _19725_/A _19890_/B _19879_/D _19797_/A VGND VGND VPWR VPWR _19727_/X sky130_fd_sc_hd__a2bb2o_4
X_16939_ _17070_/A VGND VGND VPWR VPWR _16939_/X sky130_fd_sc_hd__buf_2
XANTENNA__21915__A1 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21915__B2 _21913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19658_ _19571_/X _19639_/X _19657_/X _11611_/B _19607_/X VGND VGND VPWR VPWR _19658_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_65_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18609_ _18095_/A _18134_/X VGND VGND VPWR VPWR _18609_/Y sky130_fd_sc_hd__nor2_4
XFILLER_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19589_ _19589_/A VGND VGND VPWR VPWR _19589_/X sky130_fd_sc_hd__buf_2
XFILLER_129_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13314__A _13318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21620_ _21620_/A VGND VGND VPWR VPWR _21620_/X sky130_fd_sc_hd__buf_2
XANTENNA__17347__A1 _17339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21143__A2 _21141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21551_ _20531_/A VGND VGND VPWR VPWR _21551_/X sky130_fd_sc_hd__buf_2
XANTENNA__16625__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20502_ _18210_/X _20446_/X _20638_/A _20501_/Y VGND VGND VPWR VPWR _20502_/X sky130_fd_sc_hd__a211o_4
XFILLER_166_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24270_ _24271_/CLK _24270_/D HRESETn VGND VGND VPWR VPWR _20436_/A sky130_fd_sc_hd__dfrtp_4
X_21482_ _21482_/A VGND VGND VPWR VPWR _21482_/X sky130_fd_sc_hd__buf_2
XANTENNA__13968__B _24000_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24393__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23221_ _23392_/CLK _23221_/D VGND VGND VPWR VPWR _15033_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__11769__A _11768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20433_ _20343_/X _20432_/X _19155_/A _20352_/X VGND VGND VPWR VPWR _20433_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18847__A1 _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14145__A _11898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23152_ _24080_/CLK _23152_/D VGND VGND VPWR VPWR _16428_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_101_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20364_ _20380_/A _20364_/B VGND VGND VPWR VPWR _20364_/X sky130_fd_sc_hd__and2_4
XFILLER_162_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22362__A _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22103_ _20377_/A VGND VGND VPWR VPWR _22103_/X sky130_fd_sc_hd__buf_2
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14333__A1 _14450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17456__A _17455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23083_ _22798_/A _11647_/B _16936_/X _23083_/D VGND VGND VPWR VPWR _23084_/A sky130_fd_sc_hd__or4_4
XANTENNA__16360__A _13407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20295_ _20235_/X _20252_/X _20255_/X _20294_/Y VGND VGND VPWR VPWR _20295_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21893__A2_N _21892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14799__B _14731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22034_ _21879_/X _22031_/X _23512_/Q _22028_/X VGND VGND VPWR VPWR _23512_/D sky130_fd_sc_hd__o22a_4
XFILLER_103_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19671__A HRDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23985_ _23761_/CLK _21194_/X VGND VGND VPWR VPWR _23985_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20610__A _20438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22936_ _22910_/X VGND VGND VPWR VPWR _23079_/B sky130_fd_sc_hd__buf_2
XFILLER_95_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21382__A2 _21377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15423__B _15487_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22867_ _12753_/Y _22846_/X _22853_/X _22866_/X VGND VGND VPWR VPWR _22868_/A sky130_fd_sc_hd__a211o_4
XANTENNA__13224__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12620_ _12670_/A _12618_/X _12619_/X VGND VGND VPWR VPWR _12620_/X sky130_fd_sc_hd__and3_4
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21818_ _21817_/X _21815_/X _23634_/Q _21810_/X VGND VGND VPWR VPWR _21818_/X sky130_fd_sc_hd__o22a_4
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22798_ _22798_/A _17039_/X _20218_/A VGND VGND VPWR VPWR _22799_/A sky130_fd_sc_hd__or3_4
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18734__B _18734_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12551_ _12511_/A _12655_/B VGND VGND VPWR VPWR _12551_/X sky130_fd_sc_hd__or2_4
XANTENNA__21441__A _21441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21749_ _21589_/X _21748_/X _14567_/B _21745_/X VGND VGND VPWR VPWR _21749_/X sky130_fd_sc_hd__o22a_4
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20893__B2 _20861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15270_ _14267_/A _22350_/A VGND VGND VPWR VPWR _15270_/X sky130_fd_sc_hd__or2_4
X_12482_ _13606_/A VGND VGND VPWR VPWR _13964_/A sky130_fd_sc_hd__buf_2
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24468_ _23379_/CLK _24468_/D HRESETn VGND VGND VPWR VPWR _24468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11679__A _15377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14221_ _13865_/A _14221_/B _14220_/X VGND VGND VPWR VPWR _14221_/X sky130_fd_sc_hd__or3_4
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23419_ _23772_/CLK _22214_/X VGND VGND VPWR VPWR _14463_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22634__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24399_ _24397_/CLK _24399_/D HRESETn VGND VGND VPWR VPWR _18983_/A sky130_fd_sc_hd__dfstp_4
X_14152_ _13955_/A VGND VGND VPWR VPWR _14171_/A sky130_fd_sc_hd__buf_2
XFILLER_4_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17510__A1 _11815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24330__CLK _24342_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13103_ _13103_/A _13101_/X _13102_/X VGND VGND VPWR VPWR _13107_/B sky130_fd_sc_hd__and3_4
XANTENNA__13894__A _13894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18960_ _11544_/X VGND VGND VPWR VPWR _18960_/X sky130_fd_sc_hd__buf_2
X_14083_ _15649_/A _14066_/X _14082_/X VGND VGND VPWR VPWR _14084_/C sky130_fd_sc_hd__or3_4
XFILLER_98_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13034_ _12570_/A _13034_/B _13033_/X VGND VGND VPWR VPWR _13038_/B sky130_fd_sc_hd__and3_4
X_17911_ _18220_/A _17911_/B VGND VGND VPWR VPWR _17911_/X sky130_fd_sc_hd__or2_4
XANTENNA__22398__B2 _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18891_ _20447_/A VGND VGND VPWR VPWR _18891_/X sky130_fd_sc_hd__buf_2
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14502__B _14502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17842_ _17233_/A _17177_/X _17817_/A _17204_/X VGND VGND VPWR VPWR _17842_/X sky130_fd_sc_hd__o22a_4
XFILLER_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24480__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17773_ _17905_/A _17493_/X _17694_/X VGND VGND VPWR VPWR _17773_/X sky130_fd_sc_hd__a21bo_4
X_14985_ _14169_/A _23253_/Q VGND VGND VPWR VPWR _14985_/X sky130_fd_sc_hd__or2_4
XANTENNA__12022__B _12021_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19512_ _19512_/A VGND VGND VPWR VPWR _19512_/X sky130_fd_sc_hd__buf_2
XANTENNA__15614__A _13885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16724_ _16724_/A _24081_/Q VGND VGND VPWR VPWR _16725_/C sky130_fd_sc_hd__or2_4
X_13936_ _14390_/A _13845_/B VGND VGND VPWR VPWR _13936_/X sky130_fd_sc_hd__or2_4
XANTENNA__17577__A1 _17574_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22570__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19443_ _19442_/X VGND VGND VPWR VPWR _19480_/A sky130_fd_sc_hd__inv_2
XFILLER_62_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16655_ _16662_/A _23986_/Q VGND VGND VPWR VPWR _16655_/X sky130_fd_sc_hd__or2_4
XFILLER_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13867_ _13884_/A _13796_/B VGND VGND VPWR VPWR _13867_/X sky130_fd_sc_hd__or2_4
XFILLER_90_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13134__A _12696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15606_ _15606_/A VGND VGND VPWR VPWR _15642_/A sky130_fd_sc_hd__buf_2
X_12818_ _13562_/A _12816_/X _12817_/X VGND VGND VPWR VPWR _12818_/X sky130_fd_sc_hd__and3_4
X_19374_ _19372_/X _18671_/X _19372_/X _24249_/Q VGND VGND VPWR VPWR _24249_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16586_ _16586_/A _23506_/Q VGND VGND VPWR VPWR _16588_/B sky130_fd_sc_hd__or2_4
XANTENNA__17329__A1 _11935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22447__A _20632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13798_ _13953_/A VGND VGND VPWR VPWR _13799_/A sky130_fd_sc_hd__buf_2
X_18325_ _18310_/X _18315_/Y _18321_/X _18323_/X _18324_/Y VGND VGND VPWR VPWR _18325_/X
+ sky130_fd_sc_hd__a32o_4
X_15537_ _11900_/A _24001_/Q VGND VGND VPWR VPWR _15537_/X sky130_fd_sc_hd__or2_4
X_12749_ _11872_/A _12745_/X _12749_/C VGND VGND VPWR VPWR _12749_/X sky130_fd_sc_hd__or3_4
XFILLER_163_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18256_ _17094_/Y VGND VGND VPWR VPWR _18314_/A sky130_fd_sc_hd__buf_2
X_15468_ _12597_/A _15464_/X _15467_/X VGND VGND VPWR VPWR _15468_/X sky130_fd_sc_hd__or3_4
XANTENNA__24403__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11589__A _16901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17207_ _17165_/Y _17192_/X _15653_/X _17193_/X VGND VGND VPWR VPWR _17207_/X sky130_fd_sc_hd__o22a_4
X_14419_ _12213_/A VGND VGND VPWR VPWR _14420_/A sky130_fd_sc_hd__buf_2
XANTENNA__18829__A1 _15380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18187_ _16941_/X VGND VGND VPWR VPWR _18187_/X sky130_fd_sc_hd__buf_2
XANTENNA__19756__A HRDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15399_ _14307_/A _15399_/B VGND VGND VPWR VPWR _15399_/X sky130_fd_sc_hd__or2_4
XFILLER_116_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17138_ _14701_/Y _17115_/X _16383_/X _17116_/X VGND VGND VPWR VPWR _17138_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17069_ _16936_/X _17067_/X _22798_/A _11647_/B VGND VGND VPWR VPWR _17069_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16180__A _13413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22389__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20080_ _24479_/Q VGND VGND VPWR VPWR _20080_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21061__B2 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15524__A _12300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23770_ _23770_/CLK _21591_/X VGND VGND VPWR VPWR _14633_/B sky130_fd_sc_hd__dfxtp_4
X_20982_ _20865_/A HRDATA[17] VGND VGND VPWR VPWR _20982_/X sky130_fd_sc_hd__or2_4
XANTENNA__21364__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22561__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22721_ _20770_/A _22715_/X _23104_/Q _22719_/X VGND VGND VPWR VPWR _23104_/D sky130_fd_sc_hd__o22a_4
XPHY_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22652_ _22425_/X _22651_/X _15988_/B _22648_/X VGND VGND VPWR VPWR _23150_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21116__A2 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22357__A _22357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22313__B2 _22312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21261__A _20486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21603_ _21603_/A VGND VGND VPWR VPWR _21706_/A sky130_fd_sc_hd__buf_2
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13979__A _12467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22583_ _22480_/X _22579_/X _15129_/B _22548_/A VGND VGND VPWR VPWR _22583_/X sky130_fd_sc_hd__o22a_4
XFILLER_21_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21534_ _21534_/A VGND VGND VPWR VPWR _21534_/X sky130_fd_sc_hd__buf_2
X_24322_ _24292_/CLK _24322_/D HRESETn VGND VGND VPWR VPWR _24322_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24353__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24253_ _24248_/CLK _19368_/X HRESETn VGND VGND VPWR VPWR _24253_/Q sky130_fd_sc_hd__dfrtp_4
X_21465_ _21309_/X _21462_/X _23832_/Q _21459_/X VGND VGND VPWR VPWR _23832_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23204_ _23204_/CLK _22566_/X VGND VGND VPWR VPWR _15726_/B sky130_fd_sc_hd__dfxtp_4
X_20416_ _21824_/A VGND VGND VPWR VPWR _20416_/X sky130_fd_sc_hd__buf_2
X_24184_ _24184_/CLK _19897_/X HRESETn VGND VGND VPWR VPWR _11646_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_174_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21396_ _21275_/X _21391_/X _13405_/B _21395_/X VGND VGND VPWR VPWR _21396_/X sky130_fd_sc_hd__o22a_4
XFILLER_146_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22092__A _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23135_ _23229_/CLK _22673_/X VGND VGND VPWR VPWR _23135_/Q sky130_fd_sc_hd__dfxtp_4
X_20347_ _20270_/X VGND VGND VPWR VPWR _20347_/X sky130_fd_sc_hd__buf_2
XANTENNA__16090__A _15967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14603__A _11933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23066_ _22908_/X _23064_/X _17780_/A _23065_/X VGND VGND VPWR VPWR _23067_/B sky130_fd_sc_hd__o22a_4
XFILLER_161_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20278_ _18835_/X VGND VGND VPWR VPWR _20279_/B sky130_fd_sc_hd__inv_2
XANTENNA__24315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22017_ _22010_/A VGND VGND VPWR VPWR _22017_/X sky130_fd_sc_hd__buf_2
XANTENNA__12123__A _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11665__C _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_1_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_56_0_HCLK clkbuf_7_57_0_HCLK/A VGND VGND VPWR VPWR _23500_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_63_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14770_ _13694_/A VGND VGND VPWR VPWR _14771_/A sky130_fd_sc_hd__buf_2
X_23968_ _23523_/CLK _21218_/X VGND VGND VPWR VPWR _23968_/Q sky130_fd_sc_hd__dfxtp_4
X_11982_ _11973_/X _11982_/B VGND VGND VPWR VPWR _11982_/X sky130_fd_sc_hd__and2_4
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22552__B2 _22548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13721_ _14541_/A _13721_/B VGND VGND VPWR VPWR _13721_/X sky130_fd_sc_hd__or2_4
XFILLER_112_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22919_ _22908_/X _22918_/X _18628_/X _22914_/X VGND VGND VPWR VPWR _22920_/B sky130_fd_sc_hd__o22a_4
XFILLER_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20563__B1 _24456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18745__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23899_ _23772_/CLK _23899_/D VGND VGND VPWR VPWR _14452_/B sky130_fd_sc_hd__dfxtp_4
X_16440_ _16155_/A _16440_/B _16440_/C VGND VGND VPWR VPWR _16440_/X sky130_fd_sc_hd__and3_4
X_13652_ _13652_/A VGND VGND VPWR VPWR _15402_/A sky130_fd_sc_hd__buf_2
XANTENNA__21107__A2 _21104_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14992__B _15059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22304__B2 _22298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12603_ _12950_/A _12599_/X _12603_/C VGND VGND VPWR VPWR _12603_/X sky130_fd_sc_hd__and3_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13889__A _13916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16371_ _16333_/A _16293_/B VGND VGND VPWR VPWR _16371_/X sky130_fd_sc_hd__or2_4
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13583_ _13583_/A VGND VGND VPWR VPWR _13583_/X sky130_fd_sc_hd__buf_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18110_ _17906_/C VGND VGND VPWR VPWR _18148_/B sky130_fd_sc_hd__buf_2
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15322_ _11708_/A _15260_/B VGND VGND VPWR VPWR _15324_/B sky130_fd_sc_hd__or2_4
X_12534_ _12487_/A VGND VGND VPWR VPWR _12864_/A sky130_fd_sc_hd__buf_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19090_ _19090_/A VGND VGND VPWR VPWR _19090_/Y sky130_fd_sc_hd__inv_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18041_ _18545_/A _18041_/B VGND VGND VPWR VPWR _18042_/D sky130_fd_sc_hd__and2_4
X_15253_ _14137_/A _15253_/B VGND VGND VPWR VPWR _15253_/X sky130_fd_sc_hd__or2_4
X_12465_ _12536_/A _12465_/B _12465_/C VGND VGND VPWR VPWR _12465_/X sky130_fd_sc_hd__and3_4
XANTENNA__22607__A2 _22601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14204_ _14199_/A _23935_/Q VGND VGND VPWR VPWR _14206_/B sky130_fd_sc_hd__or2_4
XFILLER_153_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12396_ _13092_/A _12396_/B _12395_/X VGND VGND VPWR VPWR _12396_/X sky130_fd_sc_hd__and3_4
XFILLER_126_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15184_ _14302_/A _15161_/X _15168_/X _15175_/X _15183_/X VGND VGND VPWR VPWR _15184_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12020__A2 _11632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20515__A _20343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14135_ _13586_/A _14100_/X _14107_/X _14123_/X _14134_/X VGND VGND VPWR VPWR _14135_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15609__A _15625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19992_ _18670_/A VGND VGND VPWR VPWR _19992_/X sky130_fd_sc_hd__buf_2
XANTENNA__21291__B2 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18943_ _11544_/C VGND VGND VPWR VPWR _18953_/B sky130_fd_sc_hd__inv_2
X_14066_ _11780_/A _14058_/X _14065_/X VGND VGND VPWR VPWR _14066_/X sky130_fd_sc_hd__and3_4
XANTENNA__23870__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13017_ _12912_/A _12994_/X _13001_/X _13008_/X _13016_/X VGND VGND VPWR VPWR _13017_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21043__B2 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18874_ _17153_/A _18870_/X _24414_/Q _18871_/X VGND VGND VPWR VPWR _18874_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12033__A _11905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17825_ _17825_/A VGND VGND VPWR VPWR _17825_/X sky130_fd_sc_hd__buf_2
XFILLER_95_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12968__A _12944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11872__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15344__A _11735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24226__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17756_ _17748_/A _17321_/X _17748_/X _17755_/X VGND VGND VPWR VPWR _17756_/X sky130_fd_sc_hd__o22a_4
X_14968_ _14925_/X _14966_/X _14968_/C VGND VGND VPWR VPWR _14968_/X sky130_fd_sc_hd__and3_4
XANTENNA__21346__A2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18747__B1 _17820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16707_ _12051_/A _16782_/B VGND VGND VPWR VPWR _16707_/X sky130_fd_sc_hd__or2_4
X_13919_ _14385_/A _13916_/X _13919_/C VGND VGND VPWR VPWR _13920_/C sky130_fd_sc_hd__and3_4
XANTENNA__15063__B _23285_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20554__B1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17687_ _16987_/A VGND VGND VPWR VPWR _17688_/A sky130_fd_sc_hd__buf_2
X_14899_ _14170_/A _23638_/Q VGND VGND VPWR VPWR _14900_/C sky130_fd_sc_hd__or2_4
XANTENNA__18655__A _18654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19426_ _19425_/X _18618_/X _19425_/X _24220_/Q VGND VGND VPWR VPWR _24220_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16638_ _16672_/A _16638_/B VGND VGND VPWR VPWR _16638_/X sky130_fd_sc_hd__or2_4
XFILLER_23_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22177__A _22184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21081__A _21081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24376__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23250__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19357_ _19324_/A VGND VGND VPWR VPWR _19372_/A sky130_fd_sc_hd__buf_2
XANTENNA__13799__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16569_ _11973_/X _16568_/X VGND VGND VPWR VPWR _16569_/X sky130_fd_sc_hd__and2_4
X_18308_ _17688_/A _16986_/X _16988_/B VGND VGND VPWR VPWR _23009_/B sky130_fd_sc_hd__a21bo_4
XFILLER_31_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19288_ _19242_/A _19289_/A _19287_/Y VGND VGND VPWR VPWR _24293_/D sky130_fd_sc_hd__o21a_4
XFILLER_31_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22905__A _22904_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19486__A _19823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18239_ _18187_/X _19404_/A _18219_/X _18238_/X VGND VGND VPWR VPWR _18239_/X sky130_fd_sc_hd__o22a_4
XFILLER_148_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12208__A _12571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21250_ _21249_/X _21245_/X _23953_/Q _21240_/X VGND VGND VPWR VPWR _23953_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19475__A1 _20246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19475__B2 HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17718__B _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20201_ _19906_/X _18718_/X _20200_/X VGND VGND VPWR VPWR _24133_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__20085__A2 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21282__B2 _21276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21181_ _21004_/X _21176_/X _23990_/Q _21137_/X VGND VGND VPWR VPWR _23990_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15519__A _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14423__A _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20132_ _11583_/X VGND VGND VPWR VPWR _20132_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20063_ _20062_/X VGND VGND VPWR VPWR _20063_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20160__A IRQ[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12878__A _12878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11782__A _12354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15254__A _14138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23822_ _23438_/CLK _21486_/X VGND VGND VPWR VPWR _23822_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21337__A2 _21334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22534__B2 _22498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23753_ _23241_/CLK _23753_/D VGND VGND VPWR VPWR _12919_/B sky130_fd_sc_hd__dfxtp_4
X_20965_ HRDATA[2] VGND VGND VPWR VPWR _20965_/Y sky130_fd_sc_hd__inv_2
XPHY_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22704_ _20486_/A _22701_/X _12398_/B _22698_/X VGND VGND VPWR VPWR _23116_/D sky130_fd_sc_hd__o22a_4
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23684_ _23908_/CLK _23684_/D VGND VGND VPWR VPWR _23684_/Q sky130_fd_sc_hd__dfxtp_4
X_20896_ _20940_/A _20512_/B VGND VGND VPWR VPWR _20896_/X sky130_fd_sc_hd__or2_4
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17961__A1 _16935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22635_ _22484_/X _22608_/A _23157_/Q _22598_/A VGND VGND VPWR VPWR _23157_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16085__A _11671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13502__A _12402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22566_ _22449_/X _22565_/X _15726_/B _22562_/X VGND VGND VPWR VPWR _22566_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24305_ _24306_/CLK _24305_/D HRESETn VGND VGND VPWR VPWR _24305_/Q sky130_fd_sc_hd__dfrtp_4
X_21517_ _21311_/X _21513_/X _15177_/B _21482_/A VGND VGND VPWR VPWR _23799_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19396__A _19377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22497_ _22418_/X _22494_/X _16813_/B _22491_/X VGND VGND VPWR VPWR _22497_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12118__A _16079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12250_ _12250_/A VGND VGND VPWR VPWR _12251_/A sky130_fd_sc_hd__buf_2
X_21448_ _21441_/A VGND VGND VPWR VPWR _21448_/X sky130_fd_sc_hd__buf_2
XFILLER_119_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24236_ _24495_/CLK _19398_/X HRESETn VGND VGND VPWR VPWR _24236_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11957__A _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23893__CLK _23456_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15429__A _15406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24167_ _23991_/CLK _24167_/D HRESETn VGND VGND VPWR VPWR _24167_/Q sky130_fd_sc_hd__dfrtp_4
X_12181_ _12180_/X VGND VGND VPWR VPWR _12182_/B sky130_fd_sc_hd__inv_2
XANTENNA__22470__B1 _14337_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21379_ _21247_/X _21377_/X _23890_/Q _21374_/X VGND VGND VPWR VPWR _23890_/D sky130_fd_sc_hd__o22a_4
X_23118_ _23438_/CLK _22702_/X VGND VGND VPWR VPWR _23118_/Q sky130_fd_sc_hd__dfxtp_4
X_24098_ _23587_/CLK _24098_/D VGND VGND VPWR VPWR _15509_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21025__A1 _20533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15940_ _15982_/A _15940_/B VGND VGND VPWR VPWR _15940_/X sky130_fd_sc_hd__or2_4
XFILLER_135_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23049_ _22931_/A _23049_/B VGND VGND VPWR VPWR _23051_/B sky130_fd_sc_hd__nand2_4
XANTENNA__21025__B2 _20396_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24249__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21576__A2 _21566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21166__A _21152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15871_ _13520_/A _15867_/X _15871_/C VGND VGND VPWR VPWR _15879_/B sky130_fd_sc_hd__or3_4
XFILLER_62_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20070__A _19956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11692__A _13407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17610_ _17423_/A VGND VGND VPWR VPWR _17615_/A sky130_fd_sc_hd__inv_2
XFILLER_95_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14822_ _14834_/A _23385_/Q VGND VGND VPWR VPWR _14824_/B sky130_fd_sc_hd__or2_4
X_18590_ _18506_/A _18582_/X _18583_/Y _18585_/X _18589_/Y VGND VGND VPWR VPWR _18590_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21328__A2 _21327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22525__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23273__CLK _23241_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17541_ _12678_/X _17487_/B VGND VGND VPWR VPWR _17541_/Y sky130_fd_sc_hd__nand2_4
X_14753_ _15446_/A _14753_/B VGND VGND VPWR VPWR _14755_/B sky130_fd_sc_hd__or2_4
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11965_ _11965_/A VGND VGND VPWR VPWR _13981_/A sky130_fd_sc_hd__inv_2
XFILLER_17_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20000__A2 _19983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13704_ _13704_/A VGND VGND VPWR VPWR _13705_/A sky130_fd_sc_hd__buf_2
X_17472_ _17047_/A _17471_/X _17050_/X VGND VGND VPWR VPWR _17473_/A sky130_fd_sc_hd__o21a_4
X_14684_ _14684_/A _14684_/B VGND VGND VPWR VPWR _14685_/C sky130_fd_sc_hd__or2_4
X_11896_ _11895_/X VGND VGND VPWR VPWR _14110_/A sky130_fd_sc_hd__buf_2
X_19211_ _19211_/A VGND VGND VPWR VPWR _19211_/Y sky130_fd_sc_hd__inv_2
X_16423_ _16094_/A _16421_/X _16422_/X VGND VGND VPWR VPWR _16423_/X sky130_fd_sc_hd__and3_4
X_13635_ _15446_/A VGND VGND VPWR VPWR _13675_/A sky130_fd_sc_hd__buf_2
XANTENNA__14766__A1 _13951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13412__A _13379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19142_ _24321_/Q _19142_/B VGND VGND VPWR VPWR _19142_/X sky130_fd_sc_hd__and2_4
X_16354_ _16192_/A _16286_/B VGND VGND VPWR VPWR _16356_/B sky130_fd_sc_hd__or2_4
X_13566_ _13566_/A _13566_/B _13565_/X VGND VGND VPWR VPWR _13566_/X sky130_fd_sc_hd__and3_4
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21500__A2 _21499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14227__B _23967_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15305_ _14994_/A _15305_/B VGND VGND VPWR VPWR _15305_/X sky130_fd_sc_hd__or2_4
X_12517_ _12878_/A _12618_/B VGND VGND VPWR VPWR _12517_/X sky130_fd_sc_hd__or2_4
X_19073_ _19068_/X _19072_/X _19068_/X _24352_/Q VGND VGND VPWR VPWR _24352_/D sky130_fd_sc_hd__a2bb2o_4
X_16285_ _16003_/A _16281_/X _16284_/X VGND VGND VPWR VPWR _16285_/X sky130_fd_sc_hd__or3_4
X_13497_ _13547_/A _13497_/B _13496_/X VGND VGND VPWR VPWR _13497_/X sky130_fd_sc_hd__and3_4
XANTENNA__12028__A _11868_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18024_ _18070_/A _17009_/B VGND VGND VPWR VPWR _18024_/X sky130_fd_sc_hd__or2_4
X_15236_ _14201_/A _15234_/X _15235_/X VGND VGND VPWR VPWR _15236_/X sky130_fd_sc_hd__and3_4
X_12448_ _12852_/A VGND VGND VPWR VPWR _12863_/A sky130_fd_sc_hd__buf_2
XFILLER_8_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15167_ _12444_/A _15165_/X _15166_/X VGND VGND VPWR VPWR _15168_/C sky130_fd_sc_hd__and3_4
X_12379_ _13529_/A _12366_/X _12379_/C VGND VGND VPWR VPWR _12379_/X sky130_fd_sc_hd__and3_4
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14243__A _14663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14118_ _12194_/A VGND VGND VPWR VPWR _14155_/A sky130_fd_sc_hd__buf_2
X_19975_ _19962_/X _19967_/Y _19969_/X _19973_/X _19974_/Y VGND VGND VPWR VPWR _19975_/X
+ sky130_fd_sc_hd__a32o_4
X_15098_ _15106_/A _15094_/X _15098_/C VGND VGND VPWR VPWR _15098_/X sky130_fd_sc_hd__or3_4
XANTENNA__21016__A1 _20343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18926_ _15651_/X _18920_/X _19066_/A _18921_/X VGND VGND VPWR VPWR _24385_/D sky130_fd_sc_hd__o22a_4
X_14049_ _11780_/A _14041_/X _14048_/X VGND VGND VPWR VPWR _14050_/C sky130_fd_sc_hd__and3_4
XFILLER_140_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21567__A2 _21566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22764__A1 SYSTICKCLKDIV[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18857_ _18843_/A VGND VGND VPWR VPWR _18857_/X sky130_fd_sc_hd__buf_2
XFILLER_94_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15074__A _15091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17808_ _11610_/X VGND VGND VPWR VPWR _17809_/A sky130_fd_sc_hd__buf_2
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18788_ _18786_/A VGND VGND VPWR VPWR _18789_/A sky130_fd_sc_hd__inv_2
XANTENNA__22516__B2 _22512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17739_ _17738_/X _17280_/X _17734_/X VGND VGND VPWR VPWR _17739_/X sky130_fd_sc_hd__a21bo_4
XFILLER_165_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12210__B _23788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15802__A _12866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20750_ _20380_/B _20844_/B VGND VGND VPWR VPWR _20750_/X sky130_fd_sc_hd__or2_4
XFILLER_51_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19409_ _19407_/X _18278_/X _19407_/X _24232_/Q VGND VGND VPWR VPWR _19409_/X sky130_fd_sc_hd__a2bb2o_4
X_20681_ _20681_/A VGND VGND VPWR VPWR _20681_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14418__A _12299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13322__A _12516_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22420_ _22420_/A VGND VGND VPWR VPWR _22420_/X sky130_fd_sc_hd__buf_2
XFILLER_91_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22351_ _15213_/B VGND VGND VPWR VPWR _23319_/D sky130_fd_sc_hd__buf_2
XFILLER_164_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21302_ _20892_/A VGND VGND VPWR VPWR _21302_/X sky130_fd_sc_hd__buf_2
XFILLER_117_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19448__A1 HRDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22282_ _22101_/X _22280_/X _16615_/B _22277_/X VGND VGND VPWR VPWR _23378_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17448__B _17448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24021_ _23203_/CLK _21131_/X VGND VGND VPWR VPWR _24021_/Q sky130_fd_sc_hd__dfxtp_4
X_21233_ _23956_/Q VGND VGND VPWR VPWR _21233_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11777__A _11686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21255__B2 _21252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15249__A _11812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14153__A _14171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21164_ _20693_/X _21162_/X _15804_/B _21159_/X VGND VGND VPWR VPWR _24003_/D sky130_fd_sc_hd__o22a_4
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20115_ _24474_/Q VGND VGND VPWR VPWR _20115_/Y sky130_fd_sc_hd__inv_2
X_21095_ _20395_/X _21090_/X _16397_/B _21094_/X VGND VGND VPWR VPWR _21095_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20046_ _19956_/A VGND VGND VPWR VPWR _20046_/X sky130_fd_sc_hd__buf_2
XFILLER_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14600__B _14600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12401__A _12401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22507__B2 _22505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23805_ _23101_/CLK _23805_/D VGND VGND VPWR VPWR _13930_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_27_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _21813_/X _21996_/X _23539_/Q _21993_/X VGND VGND VPWR VPWR _21997_/X sky130_fd_sc_hd__o22a_4
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15712__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11750_ _11750_/A VGND VGND VPWR VPWR _15330_/A sky130_fd_sc_hd__inv_2
XFILLER_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23736_ _23098_/CLK _21651_/X VGND VGND VPWR VPWR _23736_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20470_/A _20947_/X _24376_/Q _18893_/A VGND VGND VPWR VPWR _20948_/X sky130_fd_sc_hd__o22a_4
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21730__A2 _21727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11681_/A VGND VGND VPWR VPWR _11682_/A sky130_fd_sc_hd__buf_2
X_23667_ _23760_/CLK _23667_/D VGND VGND VPWR VPWR _23667_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14328__A _13666_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20879_ _20676_/X _20876_/Y _20878_/X _19101_/Y _20731_/X VGND VGND VPWR VPWR _20880_/A
+ sky130_fd_sc_hd__a32o_4
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13427_/A _13420_/B VGND VGND VPWR VPWR _13421_/C sky130_fd_sc_hd__or2_4
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22618_ _22454_/X _22615_/X _15473_/B _22612_/X VGND VGND VPWR VPWR _23170_/D sky130_fd_sc_hd__o22a_4
X_23598_ _23918_/CLK _21903_/X VGND VGND VPWR VPWR _16039_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_139_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13351_ _13374_/A _23366_/Q VGND VGND VPWR VPWR _13354_/B sky130_fd_sc_hd__or2_4
XANTENNA__21494__B2 _21489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22549_ _22420_/X _22544_/X _16394_/B _22548_/X VGND VGND VPWR VPWR _23216_/D sky130_fd_sc_hd__o22a_4
XFILLER_128_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12302_ _11887_/A VGND VGND VPWR VPWR _13332_/A sky130_fd_sc_hd__buf_2
XFILLER_127_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16070_ _16046_/A _23822_/Q VGND VGND VPWR VPWR _16070_/X sky130_fd_sc_hd__or2_4
X_13282_ _12516_/A _13275_/X _13281_/X VGND VGND VPWR VPWR _13282_/X sky130_fd_sc_hd__or3_4
XANTENNA__24330__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15021_ _13965_/A _15019_/X _15020_/X VGND VGND VPWR VPWR _15022_/C sky130_fd_sc_hd__and3_4
XANTENNA__11687__A _13865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21246__B2 _21240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24219_ _24182_/CLK _24219_/D HRESETn VGND VGND VPWR VPWR _24219_/Q sky130_fd_sc_hd__dfrtp_4
X_12233_ _12233_/A VGND VGND VPWR VPWR _12250_/A sky130_fd_sc_hd__buf_2
XFILLER_68_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14063__A _12581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21797__A2 _21791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12164_ _12164_/A _23827_/Q VGND VGND VPWR VPWR _12165_/C sky130_fd_sc_hd__or2_4
XANTENNA__22280__A _22294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14998__A _13954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19760_ _19441_/X _19759_/X _17816_/X _19700_/X VGND VGND VPWR VPWR _19760_/X sky130_fd_sc_hd__o22a_4
X_16972_ _24135_/Q VGND VGND VPWR VPWR _17743_/A sky130_fd_sc_hd__inv_2
X_12095_ _12064_/X _24115_/Q VGND VGND VPWR VPWR _12095_/X sky130_fd_sc_hd__or2_4
XANTENNA__20512__B _20512_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22746__A1 _19519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18711_ _17974_/X _18711_/B VGND VGND VPWR VPWR _18711_/X sky130_fd_sc_hd__and2_4
X_15923_ _14086_/X _14264_/Y _14085_/X _15922_/Y VGND VGND VPWR VPWR _15923_/X sky130_fd_sc_hd__a211o_4
X_19691_ _19691_/A VGND VGND VPWR VPWR _19691_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13407__A _13407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18642_ _18641_/X VGND VGND VPWR VPWR _18642_/Y sky130_fd_sc_hd__inv_2
X_15854_ _13540_/X _15854_/B VGND VGND VPWR VPWR _15855_/C sky130_fd_sc_hd__or2_4
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_26_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14805_ _14676_/A _14802_/X _14805_/C VGND VGND VPWR VPWR _14809_/B sky130_fd_sc_hd__and3_4
XFILLER_91_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21624__A _21624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18573_ _18531_/X _18572_/X _24478_/Q _18531_/X VGND VGND VPWR VPWR _18573_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13126__B _13125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15785_ _15785_/A _15784_/X VGND VGND VPWR VPWR _15788_/A sky130_fd_sc_hd__and2_4
X_12997_ _12877_/A _12995_/X _12997_/C VGND VGND VPWR VPWR _12997_/X sky130_fd_sc_hd__and3_4
XFILLER_18_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16718__A _11973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17524_ _13270_/X _17522_/B VGND VGND VPWR VPWR _17524_/X sky130_fd_sc_hd__and2_4
X_14736_ _13617_/A _14736_/B VGND VGND VPWR VPWR _14736_/X sky130_fd_sc_hd__or2_4
X_11948_ _11939_/X _11948_/B _11947_/X VGND VGND VPWR VPWR _11948_/X sky130_fd_sc_hd__or3_4
XANTENNA__17925__A1 _17813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21182__B1 _23989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21721__A2 _21720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17455_ _17046_/A _17454_/X _17418_/A VGND VGND VPWR VPWR _17455_/X sky130_fd_sc_hd__o21a_4
X_14667_ _14667_/A _14667_/B _14667_/C VGND VGND VPWR VPWR _14667_/X sky130_fd_sc_hd__and3_4
XFILLER_162_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11879_ _11879_/A VGND VGND VPWR VPWR _11880_/A sky130_fd_sc_hd__buf_2
XANTENNA__24489__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16406_ _16409_/A _16406_/B VGND VGND VPWR VPWR _16406_/X sky130_fd_sc_hd__or2_4
XANTENNA__13142__A _13045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13618_ _15395_/A _13721_/B VGND VGND VPWR VPWR _13618_/X sky130_fd_sc_hd__or2_4
X_17386_ _17384_/X _17385_/X VGND VGND VPWR VPWR _17387_/A sky130_fd_sc_hd__or2_4
XANTENNA__24418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14598_ _13656_/A _14598_/B VGND VGND VPWR VPWR _14598_/X sky130_fd_sc_hd__or2_4
XFILLER_146_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19125_ _18959_/A _19123_/Y _24342_/Q _19124_/X VGND VGND VPWR VPWR _24342_/D sky130_fd_sc_hd__a2bb2o_4
X_16337_ _13414_/A _16331_/X _16336_/X VGND VGND VPWR VPWR _16337_/X sky130_fd_sc_hd__or3_4
X_13549_ _13529_/A _13549_/B _13548_/X VGND VGND VPWR VPWR _13565_/B sky130_fd_sc_hd__and3_4
XANTENNA__22682__B1 _23128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23169__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12981__A _12980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24414__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19056_ _24387_/Q VGND VGND VPWR VPWR _19056_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16268_ _15952_/A _16266_/X _16267_/X VGND VGND VPWR VPWR _16268_/X sky130_fd_sc_hd__and3_4
XANTENNA__13796__B _13796_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18007_ _17583_/A _18007_/B VGND VGND VPWR VPWR _18007_/X sky130_fd_sc_hd__or2_4
XANTENNA__22434__B1 _12579_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11597__A _11646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15219_ _14225_/A _15155_/B VGND VGND VPWR VPWR _15221_/B sky130_fd_sc_hd__or2_4
XANTENNA__15069__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19764__A _19823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16199_ _16181_/X _16199_/B VGND VGND VPWR VPWR _16199_/X sky130_fd_sc_hd__or2_4
XFILLER_126_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18102__B2 _18101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17284__A _14613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20460__A2 _20443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_108_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR _23111_/CLK sky130_fd_sc_hd__clkbuf_1
X_19958_ _19957_/X VGND VGND VPWR VPWR _19959_/A sky130_fd_sc_hd__buf_2
XANTENNA__14701__A _14700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20422__B _20422_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18909_ _17139_/X _18906_/X _24398_/Q _18907_/X VGND VGND VPWR VPWR _24398_/D sky130_fd_sc_hd__o22a_4
X_19889_ _19889_/A _19857_/B _19889_/C _19741_/B VGND VGND VPWR VPWR _19889_/X sky130_fd_sc_hd__and4_4
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21920_ _21906_/A VGND VGND VPWR VPWR _21920_/X sky130_fd_sc_hd__buf_2
XANTENNA__12221__A _13676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21851_ _21839_/A VGND VGND VPWR VPWR _21851_/X sky130_fd_sc_hd__buf_2
XFILLER_35_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16628__A _16646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20802_ _20772_/X _20801_/X _24095_/Q _20746_/X VGND VGND VPWR VPWR _20802_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15532__A _11886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19905__A2 _19904_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21782_ _21560_/X _21777_/X _23654_/Q _21781_/X VGND VGND VPWR VPWR _21782_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23521_ _23617_/CLK _23521_/D VGND VGND VPWR VPWR _15523_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19939__A _22745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20733_ _20732_/X VGND VGND VPWR VPWR _20733_/Y sky130_fd_sc_hd__inv_2
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20920__B1 _20917_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13052__A _13052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20664_ _20664_/A VGND VGND VPWR VPWR _20845_/A sky130_fd_sc_hd__buf_2
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23452_ _23515_/CLK _22155_/X VGND VGND VPWR VPWR _14363_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13987__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22403_ _22169_/X _22376_/A _23285_/Q _22366_/A VGND VGND VPWR VPWR _23285_/D sky130_fd_sc_hd__o22a_4
XFILLER_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21476__B2 _21475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23383_ _23383_/CLK _22269_/X VGND VGND VPWR VPWR _15165_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22673__B1 _23135_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12891__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20595_ _20595_/A VGND VGND VPWR VPWR _20596_/A sky130_fd_sc_hd__buf_2
X_22334_ _23336_/Q VGND VGND VPWR VPWR _22334_/X sky130_fd_sc_hd__buf_2
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22265_ _22258_/A VGND VGND VPWR VPWR _22265_/X sky130_fd_sc_hd__buf_2
XANTENNA__21228__B2 _21223_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21779__A2 _21777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21216_ _21202_/A VGND VGND VPWR VPWR _21216_/X sky130_fd_sc_hd__buf_2
X_24004_ _23908_/CLK _24004_/D VGND VGND VPWR VPWR _15744_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21709__A _21724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22196_ _22125_/X _22194_/X _13105_/B _22191_/X VGND VGND VPWR VPWR _22196_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18644__A2 _18633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21147_ _20416_/X _21141_/X _16339_/B _21145_/X VGND VGND VPWR VPWR _24015_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14611__A _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22728__A1 _20892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22728__B2 _22726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21078_ _21004_/X _21073_/X _14884_/B _21042_/A VGND VGND VPWR VPWR _21078_/X sky130_fd_sc_hd__o22a_4
XFILLER_76_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20203__A2 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12920_ _12972_/A _12918_/X _12919_/X VGND VGND VPWR VPWR _12921_/C sky130_fd_sc_hd__and3_4
XANTENNA__13227__A _13251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20029_ _20016_/X _16954_/Y _20022_/X _20028_/X VGND VGND VPWR VPWR _20029_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21400__B2 _21395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12131__A _11686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21951__A2 _21946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17080__A1 _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12851_ _12851_/A VGND VGND VPWR VPWR _12886_/A sky130_fd_sc_hd__buf_2
XANTENNA__11970__A _11970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15442__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11802_ _12129_/A _11802_/B _11802_/C VGND VGND VPWR VPWR _11807_/B sky130_fd_sc_hd__and3_4
X_15570_ _14430_/A _23649_/Q VGND VGND VPWR VPWR _15571_/C sky130_fd_sc_hd__or2_4
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12782_ _12800_/A _24042_/Q VGND VGND VPWR VPWR _12782_/X sky130_fd_sc_hd__or2_4
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14509_/A _14521_/B _14521_/C VGND VGND VPWR VPWR _14522_/C sky130_fd_sc_hd__and3_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23719_ _23750_/CLK _21680_/X VGND VGND VPWR VPWR _23719_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ _11653_/A VGND VGND VPWR VPWR _13717_/A sky130_fd_sc_hd__inv_2
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14058__A _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _17823_/A _17240_/B VGND VGND VPWR VPWR _17240_/X sky130_fd_sc_hd__or2_4
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _12435_/A _14452_/B VGND VGND VPWR VPWR _14452_/X sky130_fd_sc_hd__or2_4
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A _15377_/A VGND VGND VPWR VPWR _11665_/D sky130_fd_sc_hd__or2_4
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22275__A _22275_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _13376_/A _13403_/B _13402_/X VGND VGND VPWR VPWR _13407_/B sky130_fd_sc_hd__and3_4
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21467__B2 _21431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17171_ _17170_/Y _17144_/X _13270_/X _17146_/X VGND VGND VPWR VPWR _17171_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13897__A _14507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14383_ _14383_/A _14383_/B _14383_/C VGND VGND VPWR VPWR _14383_/X sky130_fd_sc_hd__and3_4
XFILLER_155_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11595_ _11595_/A VGND VGND VPWR VPWR _11596_/A sky130_fd_sc_hd__inv_2
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16122_ _16101_/A _16189_/B VGND VGND VPWR VPWR _16123_/C sky130_fd_sc_hd__or2_4
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _13290_/A _13332_/X _13333_/X VGND VGND VPWR VPWR _13334_/X sky130_fd_sc_hd__and3_4
XFILLER_155_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16053_ _16053_/A _16053_/B _16053_/C VGND VGND VPWR VPWR _16085_/B sky130_fd_sc_hd__or3_4
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19584__A _19705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13265_ _13264_/X VGND VGND VPWR VPWR _13265_/Y sky130_fd_sc_hd__inv_2
X_15004_ _13964_/A _23541_/Q VGND VGND VPWR VPWR _15005_/C sky130_fd_sc_hd__or2_4
X_12216_ _12696_/A _24044_/Q VGND VGND VPWR VPWR _12216_/X sky130_fd_sc_hd__or2_4
X_13196_ _13205_/A _23527_/Q VGND VGND VPWR VPWR _13196_/X sky130_fd_sc_hd__or2_4
X_19812_ _19687_/D _19810_/X _19507_/B _19811_/X VGND VGND VPWR VPWR _19812_/X sky130_fd_sc_hd__a211o_4
XANTENNA_clkbuf_0_HCLK_A HCLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12147_ _16053_/A _12147_/B _12146_/X VGND VGND VPWR VPWR _12147_/X sky130_fd_sc_hd__or3_4
XFILLER_2_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15617__A _13928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19743_ _19742_/X VGND VGND VPWR VPWR _19743_/Y sky130_fd_sc_hd__inv_2
X_16955_ _24151_/Q VGND VGND VPWR VPWR _16989_/A sky130_fd_sc_hd__inv_2
XFILLER_38_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12078_ _16568_/A VGND VGND VPWR VPWR _12078_/X sky130_fd_sc_hd__buf_2
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22195__A2 _22194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15906_ _13515_/X _15836_/B VGND VGND VPWR VPWR _15906_/X sky130_fd_sc_hd__or2_4
X_19674_ _19469_/X _19673_/X _17285_/Y _19515_/X VGND VGND VPWR VPWR _19674_/Y sky130_fd_sc_hd__a22oi_4
X_16886_ _12683_/X _16833_/X _12683_/X _16833_/X VGND VGND VPWR VPWR _16887_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12683__A2 _12680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15837_ _12872_/A _15837_/B VGND VGND VPWR VPWR _15838_/C sky130_fd_sc_hd__or2_4
X_18625_ _11642_/A VGND VGND VPWR VPWR _18625_/X sky130_fd_sc_hd__buf_2
XANTENNA__12976__A _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16448__A _13468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11880__A _11880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15768_ _15743_/X _23812_/Q VGND VGND VPWR VPWR _15768_/X sky130_fd_sc_hd__or2_4
X_18556_ _18555_/X VGND VGND VPWR VPWR _18556_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17507_ _18335_/B VGND VGND VPWR VPWR _17508_/B sky130_fd_sc_hd__inv_2
X_14719_ _14301_/A _14715_/X _14719_/C VGND VGND VPWR VPWR _14719_/X sky130_fd_sc_hd__or3_4
XFILLER_33_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18487_ _18314_/A _18484_/Y _18487_/C _18486_/X VGND VGND VPWR VPWR _18487_/X sky130_fd_sc_hd__or4_4
X_15699_ _12298_/A _15697_/X _15699_/C VGND VGND VPWR VPWR _15699_/X sky130_fd_sc_hd__and3_4
XANTENNA__20902__B1 _20262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17438_ _13947_/X _17438_/B VGND VGND VPWR VPWR _17438_/X sky130_fd_sc_hd__or2_4
XFILLER_162_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15385__A1 _15185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17369_ _15453_/Y _17354_/X _17027_/X _17368_/X VGND VGND VPWR VPWR _17372_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21458__B2 _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16183__A _13379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19520__B1 _19519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19108_ _19096_/X _19107_/X _19096_/X _11520_/A VGND VGND VPWR VPWR _24346_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13600__A _14296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20380_ _20380_/A _20380_/B VGND VGND VPWR VPWR _20380_/X sky130_fd_sc_hd__and2_4
XANTENNA__22913__A _22912_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19039_ _19024_/X _19037_/X _19038_/X _24358_/Q VGND VGND VPWR VPWR _19039_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12216__A _12696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22050_ _22042_/X VGND VGND VPWR VPWR _22050_/X sky130_fd_sc_hd__buf_2
XANTENNA__21529__A _21523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17726__B _17407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21001_ _20935_/A _21001_/B VGND VGND VPWR VPWR _21001_/X sky130_fd_sc_hd__or2_4
XANTENNA__15527__A _12236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21630__B2 _21624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14431__A _14431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22186__A2 _22180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22952_ _22946_/X _17006_/A _22909_/X _22951_/X VGND VGND VPWR VPWR _22952_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24353__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21933__A2 _21930_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21903_ _21826_/X _21902_/X _16039_/B _21899_/X VGND VGND VPWR VPWR _21903_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21264__A _21264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12886__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22883_ _22845_/A _22882_/X VGND VGND VPWR VPWR HWDATA[25] sky130_fd_sc_hd__nor2_4
X_21834_ _21834_/A VGND VGND VPWR VPWR _21834_/X sky130_fd_sc_hd__buf_2
XFILLER_70_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21697__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21765_ _21532_/X _21763_/X _23666_/Q _21760_/X VGND VGND VPWR VPWR _23666_/D sky130_fd_sc_hd__o22a_4
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23504_ _23533_/CLK _23504_/D VGND VGND VPWR VPWR _16435_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20716_ _20857_/A _20716_/B VGND VGND VPWR VPWR _20716_/Y sky130_fd_sc_hd__nand2_4
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24484_ _24134_/CLK _24484_/D HRESETn VGND VGND VPWR VPWR _24484_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21696_ _21584_/X _21691_/X _14399_/B _21695_/X VGND VGND VPWR VPWR _21696_/X sky130_fd_sc_hd__o22a_4
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22095__A _20298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23435_ _23558_/CLK _22192_/X VGND VGND VPWR VPWR _12657_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21449__B2 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20647_ _18891_/X VGND VGND VPWR VPWR _20647_/X sky130_fd_sc_hd__buf_2
XANTENNA__16093__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14606__A _13593_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13510__A _13564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23366_ _24102_/CLK _22299_/X VGND VGND VPWR VPWR _23366_/Q sky130_fd_sc_hd__dfxtp_4
X_20578_ _20316_/X VGND VGND VPWR VPWR _20617_/B sky130_fd_sc_hd__buf_2
XFILLER_165_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22317_ _22161_/X _22315_/X _14779_/B _22312_/X VGND VGND VPWR VPWR _22317_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12126__A _11762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23297_ _23617_/CLK _23297_/D VGND VGND VPWR VPWR _15533_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13050_ _12630_/A VGND VGND VPWR VPWR _13091_/A sky130_fd_sc_hd__buf_2
XFILLER_106_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22248_ _22226_/A VGND VGND VPWR VPWR _22248_/X sky130_fd_sc_hd__buf_2
XANTENNA__20343__A _20343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12001_ _12001_/A VGND VGND VPWR VPWR _12001_/X sky130_fd_sc_hd__buf_2
XANTENNA__11965__A _11965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21621__B2 _21617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22179_ _22208_/A VGND VGND VPWR VPWR _22194_/A sky130_fd_sc_hd__buf_2
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14341__A _13720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15156__B _15156_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16740_ _12078_/X _16740_/B _16739_/X VGND VGND VPWR VPWR _16740_/X sky130_fd_sc_hd__or3_4
X_13952_ _13952_/A _23264_/Q VGND VGND VPWR VPWR _13952_/X sky130_fd_sc_hd__or2_4
XANTENNA__13862__A1 _11969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17053__A1 _12112_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21924__A2 _21923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12903_ _12903_/A _12903_/B _12903_/C VGND VGND VPWR VPWR _12903_/X sky130_fd_sc_hd__and3_4
X_16671_ _16659_/A _16671_/B _16670_/X VGND VGND VPWR VPWR _16671_/X sky130_fd_sc_hd__and3_4
X_13883_ _12336_/A VGND VGND VPWR VPWR _13886_/A sky130_fd_sc_hd__buf_2
XANTENNA__12796__A _15778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15172__A _13617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18410_ _18409_/X VGND VGND VPWR VPWR _18410_/Y sky130_fd_sc_hd__inv_2
X_15622_ _15641_/A _15555_/B VGND VGND VPWR VPWR _15624_/B sky130_fd_sc_hd__or2_4
X_12834_ _12834_/A _24106_/Q VGND VGND VPWR VPWR _12834_/X sky130_fd_sc_hd__or2_4
X_19390_ _19389_/X _17789_/X _19389_/X _24242_/Q VGND VGND VPWR VPWR _19390_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18341_ _18341_/A VGND VGND VPWR VPWR _18443_/B sky130_fd_sc_hd__inv_2
XANTENNA__13404__B _23718_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21902__A _21909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15553_ _12304_/A _23969_/Q VGND VGND VPWR VPWR _15554_/C sky130_fd_sc_hd__or2_4
XFILLER_15_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12634_/A VGND VGND VPWR VPWR _13058_/A sky130_fd_sc_hd__buf_2
XANTENNA__18483__A _18483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14383_/A _14502_/X _14503_/X VGND VGND VPWR VPWR _14504_/X sky130_fd_sc_hd__and3_4
X_11716_ _16031_/A VGND VGND VPWR VPWR _16079_/A sky130_fd_sc_hd__buf_2
XANTENNA__15900__A _13546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _18255_/X _18261_/Y _18268_/X _18270_/X _18271_/Y VGND VGND VPWR VPWR _18272_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _12354_/A _15476_/X _15483_/X VGND VGND VPWR VPWR _15485_/C sky130_fd_sc_hd__and3_4
X_12696_ _12696_/A _24042_/Q VGND VGND VPWR VPWR _12698_/B sky130_fd_sc_hd__or2_4
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17223_ _18772_/A _17090_/X VGND VGND VPWR VPWR _18265_/A sky130_fd_sc_hd__nand2_4
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ _12461_/A _14431_/X _14435_/C VGND VGND VPWR VPWR _14435_/X sky130_fd_sc_hd__or3_4
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _11592_/X _11647_/B _17017_/A _16936_/A VGND VGND VPWR VPWR _16926_/B sky130_fd_sc_hd__or4_4
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13420__A _13427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17154_ _17153_/Y _17131_/X _12680_/X _17133_/X VGND VGND VPWR VPWR _17154_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14366_ _14366_/A _14366_/B VGND VGND VPWR VPWR _14368_/B sky130_fd_sc_hd__or2_4
XFILLER_11_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15119__B2 _15118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11578_ _24464_/Q IRQ[27] _20186_/A VGND VGND VPWR VPWR _20142_/A sky130_fd_sc_hd__a21o_4
XANTENNA__14235__B _23135_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16105_ _15967_/A _16177_/B VGND VGND VPWR VPWR _16107_/B sky130_fd_sc_hd__or2_4
XFILLER_156_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16867__A1 _15048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13317_ _13313_/A _23846_/Q VGND VGND VPWR VPWR _13317_/X sky130_fd_sc_hd__or2_4
X_17085_ _17085_/A _18220_/A VGND VGND VPWR VPWR _17085_/X sky130_fd_sc_hd__or2_4
XFILLER_115_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14297_ _14297_/A _14297_/B _14297_/C VGND VGND VPWR VPWR _14297_/X sky130_fd_sc_hd__and3_4
XANTENNA__12036__A _16702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16036_ _11759_/X _16029_/X _16036_/C VGND VGND VPWR VPWR _16037_/C sky130_fd_sc_hd__or3_4
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13248_ _13248_/A _23719_/Q VGND VGND VPWR VPWR _13250_/B sky130_fd_sc_hd__or2_4
XANTENNA__11875__A _16159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15347__A _11673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13179_ _11888_/A _13179_/B VGND VGND VPWR VPWR _13181_/B sky130_fd_sc_hd__or2_4
XFILLER_123_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17987_ _17819_/X _17839_/X _17945_/X _17841_/X VGND VGND VPWR VPWR _17987_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22168__A2 _22159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19726_ _19684_/X _19725_/X _19899_/A VGND VGND VPWR VPWR _19726_/Y sky130_fd_sc_hd__a21oi_4
X_16938_ _17038_/A _16937_/X VGND VGND VPWR VPWR _17070_/A sky130_fd_sc_hd__or2_4
XANTENNA__20179__A1 _24456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21915__A2 _21909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19657_ _19781_/A _19657_/B _19657_/C _19656_/X VGND VGND VPWR VPWR _19657_/X sky130_fd_sc_hd__or4_4
X_16869_ _14705_/X _16868_/X _14705_/X _16868_/X VGND VGND VPWR VPWR _16869_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18792__A1 _12180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15082__A _15106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18608_ _18519_/X _18607_/Y _17308_/X VGND VGND VPWR VPWR _18608_/X sky130_fd_sc_hd__o21a_4
XFILLER_164_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19588_ _19539_/A _19533_/B _19588_/C VGND VGND VPWR VPWR _19589_/A sky130_fd_sc_hd__or3_4
XANTENNA__22908__A _22908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21679__B2 _21674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19489__A _19539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18539_ _18538_/X _18510_/X _18538_/X _18507_/X VGND VGND VPWR VPWR _18539_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21550_ _21548_/X _21542_/X _23787_/Q _21549_/X VGND VGND VPWR VPWR _21550_/X sky130_fd_sc_hd__o22a_4
X_20501_ _20501_/A _20501_/B VGND VGND VPWR VPWR _20501_/Y sky130_fd_sc_hd__nor2_4
X_21481_ _21249_/X _21478_/X _23825_/Q _21475_/X VGND VGND VPWR VPWR _23825_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22628__B1 _14502_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14426__A _14430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13330__A _13330_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20432_ _20344_/X _20431_/X _24366_/Q _20269_/X VGND VGND VPWR VPWR _20432_/X sky130_fd_sc_hd__o22a_4
X_23220_ _23476_/CLK _23220_/D VGND VGND VPWR VPWR _11763_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22643__A _22672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23151_ _23119_/CLK _23151_/D VGND VGND VPWR VPWR _16286_/B sky130_fd_sc_hd__dfxtp_4
X_20363_ _18779_/X VGND VGND VPWR VPWR _20380_/A sky130_fd_sc_hd__buf_2
XFILLER_173_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16641__A _16659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_0_0_HCLK clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_134_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22102_ _22101_/X _22099_/X _16640_/B _22094_/X VGND VGND VPWR VPWR _22102_/X sky130_fd_sc_hd__o22a_4
X_23082_ _23081_/X VGND VGND VPWR VPWR HADDR[31] sky130_fd_sc_hd__inv_2
X_20294_ _20293_/X VGND VGND VPWR VPWR _20294_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24132__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11785__A _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22033_ _21877_/X _22031_/X _23513_/Q _22028_/X VGND VGND VPWR VPWR _23513_/D sky130_fd_sc_hd__o22a_4
XFILLER_103_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19952__A _19951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15257__A _15257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14161__A _14267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24282__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23984_ _24080_/CLK _23984_/D VGND VGND VPWR VPWR _16422_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22935_ _23078_/A _22935_/B _22934_/X VGND VGND VPWR VPWR _22939_/B sky130_fd_sc_hd__or3_4
XFILLER_17_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15046__B1 _11603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21119__B1 _24031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22866_ _17284_/Y _22800_/Y _22815_/X VGND VGND VPWR VPWR _22866_/X sky130_fd_sc_hd__o21a_4
XFILLER_25_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13224__B _13148_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21817_ _21532_/A VGND VGND VPWR VPWR _21817_/X sky130_fd_sc_hd__buf_2
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19399__A _19428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22797_ _22796_/X VGND VGND VPWR VPWR _24125_/D sky130_fd_sc_hd__inv_2
XANTENNA__16816__A _16682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15720__A _12762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _12869_/A _12548_/X _12549_/X VGND VGND VPWR VPWR _12550_/X sky130_fd_sc_hd__and3_4
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21748_ _21741_/A VGND VGND VPWR VPWR _21748_/X sky130_fd_sc_hd__buf_2
XFILLER_106_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _12194_/A VGND VGND VPWR VPWR _13606_/A sky130_fd_sc_hd__buf_2
X_24467_ _23379_/CLK _24467_/D HRESETn VGND VGND VPWR VPWR _24467_/Q sky130_fd_sc_hd__dfrtp_4
X_21679_ _21556_/X _21677_/X _23720_/Q _21674_/X VGND VGND VPWR VPWR _21679_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14336__A _13884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_16_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR _24495_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ _12336_/A _14218_/X _14220_/C VGND VGND VPWR VPWR _14220_/X sky130_fd_sc_hd__and3_4
XFILLER_32_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23418_ _23772_/CLK _22216_/X VGND VGND VPWR VPWR _23418_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24398_ _24398_/CLK _24398_/D HRESETn VGND VGND VPWR VPWR _24398_/Q sky130_fd_sc_hd__dfstp_4
Xclkbuf_7_79_0_HCLK clkbuf_7_79_0_HCLK/A VGND VGND VPWR VPWR _23101_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_165_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21842__A1 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14151_ _14133_/A VGND VGND VPWR VPWR _14277_/A sky130_fd_sc_hd__buf_2
XANTENNA__21842__B2 _21834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23349_ _23617_/CLK _23349_/D VGND VGND VPWR VPWR _23349_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16551__A _11891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13102_ _13095_/A _23848_/Q VGND VGND VPWR VPWR _13102_/X sky130_fd_sc_hd__or2_4
XANTENNA__21169__A _21136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14082_ _11680_/A _14074_/X _14082_/C VGND VGND VPWR VPWR _14082_/X sky130_fd_sc_hd__and3_4
XFILLER_140_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22398__A2 _22397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13033_ _12569_/A _24104_/Q VGND VGND VPWR VPWR _13033_/X sky130_fd_sc_hd__or2_4
X_17910_ _17780_/A _17909_/A _24159_/Q _17909_/Y VGND VGND VPWR VPWR _17910_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15167__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18890_ _20274_/A VGND VGND VPWR VPWR _20447_/A sky130_fd_sc_hd__buf_2
XFILLER_26_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17841_ _17233_/A _17174_/X _17817_/A _17176_/X VGND VGND VPWR VPWR _17841_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20801__A _20801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17772_ _17772_/A _17771_/Y VGND VGND VPWR VPWR _18301_/A sky130_fd_sc_hd__or2_4
XFILLER_47_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14984_ _14984_/A VGND VGND VPWR VPWR _17339_/A sky130_fd_sc_hd__buf_2
X_19511_ _19558_/A _19503_/X _19510_/X VGND VGND VPWR VPWR _19511_/Y sky130_fd_sc_hd__o21ai_4
X_13935_ _12367_/A _13931_/X _13934_/X VGND VGND VPWR VPWR _13935_/X sky130_fd_sc_hd__or3_4
X_16723_ _16700_/A _23633_/Q VGND VGND VPWR VPWR _16725_/B sky130_fd_sc_hd__or2_4
XFILLER_75_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16654_ _16654_/A _23922_/Q VGND VGND VPWR VPWR _16654_/X sky130_fd_sc_hd__or2_4
X_19442_ _18576_/B _24128_/Q VGND VGND VPWR VPWR _19442_/X sky130_fd_sc_hd__or2_4
XFILLER_170_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13866_ _13866_/A VGND VGND VPWR VPWR _13884_/A sky130_fd_sc_hd__buf_2
X_15605_ _15641_/A _15546_/B VGND VGND VPWR VPWR _15605_/X sky130_fd_sc_hd__or2_4
X_12817_ _12775_/A _12817_/B VGND VGND VPWR VPWR _12817_/X sky130_fd_sc_hd__or2_4
X_16585_ _16593_/A VGND VGND VPWR VPWR _16586_/A sky130_fd_sc_hd__buf_2
X_19373_ _19369_/X _18665_/X _19372_/X _24250_/Q VGND VGND VPWR VPWR _24250_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13797_ _12450_/X VGND VGND VPWR VPWR _13953_/A sky130_fd_sc_hd__buf_2
XANTENNA__16726__A _16592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19723__B1 _20866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18526__B2 _18525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15536_ _14420_/A _23681_/Q VGND VGND VPWR VPWR _15536_/X sky130_fd_sc_hd__or2_4
X_18324_ _17527_/D _18322_/X _18060_/X VGND VGND VPWR VPWR _18324_/Y sky130_fd_sc_hd__a21oi_4
X_12748_ _12748_/A _12746_/X _12747_/X VGND VGND VPWR VPWR _12749_/C sky130_fd_sc_hd__and3_4
X_18255_ _18310_/A _17461_/X VGND VGND VPWR VPWR _18255_/X sky130_fd_sc_hd__or2_4
XFILLER_72_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15467_ _12650_/A _15465_/X _15467_/C VGND VGND VPWR VPWR _15467_/X sky130_fd_sc_hd__and3_4
X_12679_ _12678_/X VGND VGND VPWR VPWR _12679_/Y sky130_fd_sc_hd__inv_2
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14246__A _14201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13150__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17206_ _17160_/A _17204_/X _17164_/A _17205_/X VGND VGND VPWR VPWR _17206_/X sky130_fd_sc_hd__o22a_4
X_14418_ _12299_/A VGND VGND VPWR VPWR _14418_/X sky130_fd_sc_hd__buf_2
XFILLER_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18186_ _18145_/X _18185_/X _20017_/A _18145_/X VGND VGND VPWR VPWR _24492_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22086__B2 _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15398_ _15398_/A _15398_/B _15398_/C VGND VGND VPWR VPWR _15398_/X sky130_fd_sc_hd__or3_4
XANTENNA__24155__CLK _24306_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12574__A1 _11857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12574__B2 _12573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17137_ _16710_/A VGND VGND VPWR VPWR _17137_/X sky130_fd_sc_hd__buf_2
XANTENNA__17557__A _11611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14349_ _14516_/A _14349_/B VGND VGND VPWR VPWR _14349_/X sky130_fd_sc_hd__or2_4
XFILLER_156_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17068_ _17016_/C VGND VGND VPWR VPWR _22798_/A sky130_fd_sc_hd__buf_2
XFILLER_170_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22389__A2 _22383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16019_ _16047_/A _16017_/X _16018_/X VGND VGND VPWR VPWR _16019_/X sky130_fd_sc_hd__and3_4
XFILLER_112_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21061__A2 _21059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15805__A _12889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17292__A _17290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19709_ _19742_/A _19889_/C VGND VGND VPWR VPWR _19709_/X sky130_fd_sc_hd__or2_4
X_20981_ _20894_/X _20980_/X _15170_/B _20396_/A VGND VGND VPWR VPWR _24087_/D sky130_fd_sc_hd__o22a_4
XFILLER_65_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_0_0_HCLK_A clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22561__A2 _22558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22720_ _20745_/A _22715_/X _15634_/B _22719_/X VGND VGND VPWR VPWR _23105_/D sky130_fd_sc_hd__o22a_4
XPHY_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21542__A _21542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22651_ _22658_/A VGND VGND VPWR VPWR _22651_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16636__A _11768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22313__A2 _22308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21602_ _23764_/Q VGND VGND VPWR VPWR _21602_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22582_ _22478_/X _22579_/X _15260_/B _22576_/X VGND VGND VPWR VPWR _23192_/D sky130_fd_sc_hd__o22a_4
XFILLER_159_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20158__A IRQ[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24321_ _24292_/CLK _24321_/D HRESETn VGND VGND VPWR VPWR _24321_/Q sky130_fd_sc_hd__dfrtp_4
X_21533_ _21532_/X _21530_/X _23794_/Q _21525_/X VGND VGND VPWR VPWR _23794_/D sky130_fd_sc_hd__o22a_4
XFILLER_166_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19947__A _22908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14156__A _14170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24252_ _24248_/CLK _19370_/X HRESETn VGND VGND VPWR VPWR _24252_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22077__B2 _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21464_ _21307_/X _21462_/X _14744_/B _21459_/X VGND VGND VPWR VPWR _21464_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22373__A _22358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23203_ _23203_/CLK _22567_/X VGND VGND VPWR VPWR _15796_/B sky130_fd_sc_hd__dfxtp_4
X_20415_ _20415_/A VGND VGND VPWR VPWR _21824_/A sky130_fd_sc_hd__buf_2
XANTENNA__17467__A _12842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21395_ _21388_/A VGND VGND VPWR VPWR _21395_/X sky130_fd_sc_hd__buf_2
X_24183_ _23671_/CLK _19901_/Y HRESETn VGND VGND VPWR VPWR _11593_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23134_ _23229_/CLK _22674_/X VGND VGND VPWR VPWR _13757_/B sky130_fd_sc_hd__dfxtp_4
X_20346_ _20277_/X _20345_/X _24402_/Q _18894_/B VGND VGND VPWR VPWR _20346_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23065_ _19924_/A _17902_/Y _22929_/A VGND VGND VPWR VPWR _23065_/X sky130_fd_sc_hd__o21a_4
X_20277_ _20470_/A VGND VGND VPWR VPWR _20277_/X sky130_fd_sc_hd__buf_2
XANTENNA__12404__A _15851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22820__B _15048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22016_ _21848_/X _22010_/X _13420_/B _22014_/X VGND VGND VPWR VPWR _23525_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21717__A _21717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11665__D _11665_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15715__A _11864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22001__B2 _22000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23967_ _23323_/CLK _23967_/D VGND VGND VPWR VPWR _23967_/Q sky130_fd_sc_hd__dfxtp_4
X_11981_ _16568_/A _11977_/X _11980_/X VGND VGND VPWR VPWR _11982_/B sky130_fd_sc_hd__or3_4
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22552__A2 _22551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13235__A _13235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24028__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13720_ _13720_/A VGND VGND VPWR VPWR _13752_/A sky130_fd_sc_hd__buf_2
X_22918_ _19924_/A _16970_/A _18718_/X _18696_/X _22930_/A VGND VGND VPWR VPWR _22918_/X
+ sky130_fd_sc_hd__o32a_4
X_23898_ _24090_/CLK _21363_/X VGND VGND VPWR VPWR _14583_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22548__A _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21452__A _21438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13651_ _14480_/A _13611_/X _13626_/X _13641_/X _13650_/X VGND VGND VPWR VPWR _13651_/X
+ sky130_fd_sc_hd__a32o_4
X_22849_ _22801_/X VGND VGND VPWR VPWR _22849_/X sky130_fd_sc_hd__buf_2
XANTENNA__16546__A _11951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22304__A2 _22301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12602_ _12644_/A _23787_/Q VGND VGND VPWR VPWR _12603_/C sky130_fd_sc_hd__or2_4
XANTENNA__15450__A _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16370_ _13392_/A VGND VGND VPWR VPWR _16370_/X sky130_fd_sc_hd__buf_2
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13582_ _13582_/A _13582_/B VGND VGND VPWR VPWR _16831_/A sky130_fd_sc_hd__or2_4
XANTENNA__13889__B _24029_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24178__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ _15321_/A _15317_/X _15321_/C VGND VGND VPWR VPWR _15331_/B sky130_fd_sc_hd__or3_4
X_12533_ _12891_/A _12533_/B VGND VGND VPWR VPWR _12536_/B sky130_fd_sc_hd__or2_4
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14066__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17731__A2 _17399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18040_ _18440_/A VGND VGND VPWR VPWR _18545_/A sky130_fd_sc_hd__buf_2
X_15252_ _15252_/A VGND VGND VPWR VPWR _15252_/X sky130_fd_sc_hd__buf_2
X_12464_ _12885_/A _23787_/Q VGND VGND VPWR VPWR _12465_/C sky130_fd_sc_hd__or2_4
XANTENNA__22068__B2 _22064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14203_ _14614_/A _14192_/X _14203_/C VGND VGND VPWR VPWR _14223_/B sky130_fd_sc_hd__and3_4
XANTENNA__17377__A _17360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15183_ _13853_/A _15182_/X VGND VGND VPWR VPWR _15183_/X sky130_fd_sc_hd__and2_4
XFILLER_137_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12395_ _15894_/A _12391_/X _12394_/X VGND VGND VPWR VPWR _12395_/X sky130_fd_sc_hd__or3_4
XANTENNA_clkbuf_4_11_0_HCLK_A clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12020__A3 _11983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14134_ _15281_/A _14133_/X VGND VGND VPWR VPWR _14134_/X sky130_fd_sc_hd__and2_4
XFILLER_126_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18692__B1 _18335_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21291__A2 _21281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19991_ _19991_/A VGND VGND VPWR VPWR _24160_/D sky130_fd_sc_hd__inv_2
X_18942_ _16866_/X _18897_/A _24373_/Q _18900_/A VGND VGND VPWR VPWR _24373_/D sky130_fd_sc_hd__o22a_4
X_14065_ _14074_/A _14065_/B _14065_/C VGND VGND VPWR VPWR _14065_/X sky130_fd_sc_hd__or3_4
XANTENNA__12314__A _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_9_0_HCLK clkbuf_6_4_0_HCLK/X VGND VGND VPWR VPWR _24419_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21579__B1 _23775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13016_ _13016_/A _13016_/B VGND VGND VPWR VPWR _13016_/X sky130_fd_sc_hd__and2_4
XANTENNA__21627__A _21620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21043__A2 _21038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22240__B2 _22234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18873_ _14261_/A _18870_/X _24415_/Q _18871_/X VGND VGND VPWR VPWR _18873_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20531__A _20531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17824_ _17823_/X VGND VGND VPWR VPWR _17824_/X sky130_fd_sc_hd__buf_2
XANTENNA__15625__A _15625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17755_ _17749_/A _17329_/X _17749_/X _18721_/A VGND VGND VPWR VPWR _17755_/X sky130_fd_sc_hd__o22a_4
X_14967_ _14967_/A _14967_/B VGND VGND VPWR VPWR _14968_/C sky130_fd_sc_hd__or2_4
XFILLER_94_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14481__A1 _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13145__A _13145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16706_ _16725_/A _16706_/B _16706_/C VGND VGND VPWR VPWR _16710_/B sky130_fd_sc_hd__and3_4
X_13918_ _13937_/A _24061_/Q VGND VGND VPWR VPWR _13919_/C sky130_fd_sc_hd__or2_4
XFILLER_81_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17686_ _17686_/A _17511_/X VGND VGND VPWR VPWR _17691_/A sky130_fd_sc_hd__and2_4
X_14898_ _14165_/A _23222_/Q VGND VGND VPWR VPWR _14898_/X sky130_fd_sc_hd__or2_4
XFILLER_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19425_ _19428_/A VGND VGND VPWR VPWR _19425_/X sky130_fd_sc_hd__buf_2
XFILLER_39_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21362__A _21322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13849_ _13676_/A _23645_/Q VGND VGND VPWR VPWR _13849_/X sky130_fd_sc_hd__or2_4
X_16637_ _16788_/A VGND VGND VPWR VPWR _16672_/A sky130_fd_sc_hd__buf_2
XANTENNA__16456__A _13377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15360__A _11735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19356_ _19354_/X _18397_/X _19354_/X _24261_/Q VGND VGND VPWR VPWR _24261_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21081__B _22039_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16568_ _16568_/A _16568_/B _16568_/C VGND VGND VPWR VPWR _16568_/X sky130_fd_sc_hd__or3_4
XFILLER_128_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18307_ _17900_/A VGND VGND VPWR VPWR _18307_/X sky130_fd_sc_hd__buf_2
X_15519_ _15453_/Y _15517_/X VGND VGND VPWR VPWR _15519_/X sky130_fd_sc_hd__or2_4
X_16499_ _16507_/A _16497_/X _16498_/X VGND VGND VPWR VPWR _16499_/X sky130_fd_sc_hd__and3_4
X_19287_ _19243_/B VGND VGND VPWR VPWR _19287_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17183__B1 _15252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22059__B2 _22057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18238_ _18221_/X _18226_/Y _18232_/X _18236_/X _18237_/Y VGND VGND VPWR VPWR _18238_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_15_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20609__A2 _20599_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16191__A _11714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18169_ _17452_/X VGND VGND VPWR VPWR _18169_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14704__A _14613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_62_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR _24074_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20200_ _20200_/A _20200_/B VGND VGND VPWR VPWR _20200_/X sky130_fd_sc_hd__or2_4
XFILLER_143_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21282__A2 _21281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21180_ _20980_/X _21176_/X _15211_/B _21137_/X VGND VGND VPWR VPWR _23991_/D sky130_fd_sc_hd__o22a_4
XFILLER_85_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15519__B _15517_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22921__A _22912_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20131_ _19956_/X _20130_/X _19402_/X _24135_/Q VGND VGND VPWR VPWR _24135_/D sky130_fd_sc_hd__o22a_4
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21537__A _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18435__B1 _18027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20062_ _20040_/X _18368_/A _20046_/X _20061_/X VGND VGND VPWR VPWR _20062_/X sky130_fd_sc_hd__o22a_4
XFILLER_98_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22231__B2 _22227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15535__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23821_ _24077_/CLK _23821_/D VGND VGND VPWR VPWR _16224_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13055__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23752_ _23496_/CLK _23752_/D VGND VGND VPWR VPWR _23752_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20964_ _20943_/A _20963_/X VGND VGND VPWR VPWR _20964_/X sky130_fd_sc_hd__and2_4
XPHY_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21742__B1 _23679_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22703_ _20464_/A _22701_/X _23117_/Q _22698_/X VGND VGND VPWR VPWR _22703_/X sky130_fd_sc_hd__o22a_4
XPHY_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23683_ _23656_/CLK _21736_/X VGND VGND VPWR VPWR _15803_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24320__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ _20895_/A VGND VGND VPWR VPWR _20895_/X sky130_fd_sc_hd__buf_2
XANTENNA__15270__A _14267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22634_ _22482_/X _22629_/X _23158_/Q _22598_/A VGND VGND VPWR VPWR _23158_/D sky130_fd_sc_hd__o22a_4
XFILLER_110_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22565_ _22558_/A VGND VGND VPWR VPWR _22565_/X sky130_fd_sc_hd__buf_2
XANTENNA__18910__A1 _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24304_ _24306_/CLK _24304_/D HRESETn VGND VGND VPWR VPWR _19253_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_142_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24470__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21516_ _21309_/X _21513_/X _15305_/B _21510_/X VGND VGND VPWR VPWR _23800_/D sky130_fd_sc_hd__o22a_4
XFILLER_10_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22496_ _22416_/X _22494_/X _16679_/B _22491_/X VGND VGND VPWR VPWR _22496_/X sky130_fd_sc_hd__o22a_4
X_24235_ _24240_/CLK _24235_/D HRESETn VGND VGND VPWR VPWR _24235_/Q sky130_fd_sc_hd__dfrtp_4
X_21447_ _21278_/X _21441_/X _23845_/Q _21445_/X VGND VGND VPWR VPWR _23845_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24166_ _23991_/CLK _19943_/X HRESETn VGND VGND VPWR VPWR _24166_/Q sky130_fd_sc_hd__dfrtp_4
X_12180_ _12180_/A VGND VGND VPWR VPWR _12180_/X sky130_fd_sc_hd__buf_2
XANTENNA__15429__B _15493_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21378_ _21243_/X _21377_/X _23891_/Q _21374_/X VGND VGND VPWR VPWR _21378_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22470__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23117_ _24077_/CLK _22703_/X VGND VGND VPWR VPWR _23117_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20329_ _20313_/X _20329_/B VGND VGND VPWR VPWR _20329_/Y sky130_fd_sc_hd__nor2_4
XFILLER_123_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24097_ _23523_/CLK _20747_/X VGND VGND VPWR VPWR _24097_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_110_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23048_ _23048_/A VGND VGND VPWR VPWR _23048_/X sky130_fd_sc_hd__buf_2
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11973__A _16130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15445__A _11878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15870_ _13503_/X _15868_/X _15870_/C VGND VGND VPWR VPWR _15871_/C sky130_fd_sc_hd__and3_4
XFILLER_23_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14821_ _15112_/A _14821_/B _14821_/C VGND VGND VPWR VPWR _14821_/X sky130_fd_sc_hd__and3_4
XFILLER_92_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18756__A _18413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19926__B1 _20246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17540_ _17490_/B _17538_/Y _17539_/X VGND VGND VPWR VPWR _17540_/X sky130_fd_sc_hd__o21a_4
X_14752_ _12251_/A _14752_/B _14751_/X VGND VGND VPWR VPWR _14756_/B sky130_fd_sc_hd__and3_4
X_11964_ _12108_/A _11964_/B _11964_/C VGND VGND VPWR VPWR _11964_/X sky130_fd_sc_hd__or3_4
XFILLER_17_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13703_ _12327_/A VGND VGND VPWR VPWR _13704_/A sky130_fd_sc_hd__buf_2
X_17471_ _11867_/X _17035_/A VGND VGND VPWR VPWR _17471_/X sky130_fd_sc_hd__and2_4
X_14683_ _14653_/A _14604_/B VGND VGND VPWR VPWR _14683_/X sky130_fd_sc_hd__or2_4
X_11895_ _12194_/A VGND VGND VPWR VPWR _11895_/X sky130_fd_sc_hd__buf_2
X_19210_ _19137_/A _19211_/A _19209_/Y VGND VGND VPWR VPWR _24316_/D sky130_fd_sc_hd__o21a_4
XANTENNA__15180__A _13953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22289__A1 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16422_ _16009_/X _16422_/B VGND VGND VPWR VPWR _16422_/X sky130_fd_sc_hd__or2_4
X_13634_ _11623_/A VGND VGND VPWR VPWR _15446_/A sky130_fd_sc_hd__buf_2
XANTENNA__22289__B2 _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16353_ _13414_/A _16349_/X _16352_/X VGND VGND VPWR VPWR _16353_/X sky130_fd_sc_hd__or3_4
X_19141_ _19141_/A _19141_/B VGND VGND VPWR VPWR _19142_/B sky130_fd_sc_hd__and2_4
X_13565_ _13416_/A _13565_/B _13565_/C VGND VGND VPWR VPWR _13565_/X sky130_fd_sc_hd__or3_4
XFILLER_158_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12309__A _12300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18901__A1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15304_ _14169_/A _15304_/B VGND VGND VPWR VPWR _15306_/B sky130_fd_sc_hd__or2_4
X_12516_ _12516_/A _12508_/X _12516_/C VGND VGND VPWR VPWR _12516_/X sky130_fd_sc_hd__or3_4
X_19072_ _19046_/X _19070_/Y _19071_/Y _19049_/X VGND VGND VPWR VPWR _19072_/X sky130_fd_sc_hd__o22a_4
X_16284_ _15936_/X _16282_/X _16283_/X VGND VGND VPWR VPWR _16284_/X sky130_fd_sc_hd__and3_4
XFILLER_118_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13496_ _13496_/A _23749_/Q VGND VGND VPWR VPWR _13496_/X sky130_fd_sc_hd__or2_4
XFILLER_146_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18023_ _16950_/Y VGND VGND VPWR VPWR _18070_/A sky130_fd_sc_hd__buf_2
X_15235_ _15198_/X _15177_/B VGND VGND VPWR VPWR _15235_/X sky130_fd_sc_hd__or2_4
X_12447_ _12877_/A VGND VGND VPWR VPWR _12536_/A sky130_fd_sc_hd__buf_2
XFILLER_126_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20245__B HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_49_0_HCLK clkbuf_6_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15166_ _12453_/A _15166_/B VGND VGND VPWR VPWR _15166_/X sky130_fd_sc_hd__or2_4
X_12378_ _15894_/A _12371_/X _12378_/C VGND VGND VPWR VPWR _12379_/C sky130_fd_sc_hd__or3_4
XFILLER_158_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22741__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14117_ _14154_/A _14117_/B VGND VGND VPWR VPWR _14117_/X sky130_fd_sc_hd__or2_4
XANTENNA__20472__B1 _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19974_ _19973_/A _19972_/X _18009_/X VGND VGND VPWR VPWR _19974_/Y sky130_fd_sc_hd__a21oi_4
X_15097_ _15081_/A _15095_/X _15097_/C VGND VGND VPWR VPWR _15098_/C sky130_fd_sc_hd__and3_4
XANTENNA__12044__A _16568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18925_ _17169_/X _18920_/X _24386_/Q _18921_/X VGND VGND VPWR VPWR _24386_/D sky130_fd_sc_hd__o22a_4
X_14048_ _14074_/A _14044_/X _14048_/C VGND VGND VPWR VPWR _14048_/X sky130_fd_sc_hd__or3_4
XANTENNA__22213__B2 _22212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12979__A _12979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20261__A _20233_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11883__A _11882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18856_ _18840_/A VGND VGND VPWR VPWR _18856_/X sky130_fd_sc_hd__buf_2
XFILLER_95_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17807_ _17807_/A VGND VGND VPWR VPWR _17807_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_4_0_HCLK clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_8_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24343__CLK _24342_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18787_ _18796_/A VGND VGND VPWR VPWR _18787_/X sky130_fd_sc_hd__buf_2
X_15999_ _15998_/X VGND VGND VPWR VPWR _16110_/A sky130_fd_sc_hd__buf_2
XANTENNA__19917__B1 _22904_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17570__A _16085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17738_ _17734_/A VGND VGND VPWR VPWR _17738_/X sky130_fd_sc_hd__buf_2
X_17669_ _17669_/A _17567_/X VGND VGND VPWR VPWR _17669_/X sky130_fd_sc_hd__or2_4
XFILLER_91_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15090__A _15112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19408_ _19396_/X _18254_/X _19407_/X _24233_/Q VGND VGND VPWR VPWR _19408_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24493__CLK _24306_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20680_ _20676_/X _20677_/Y _20679_/X _19056_/Y _20495_/X VGND VGND VPWR VPWR _20681_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_52_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19339_ _19324_/A VGND VGND VPWR VPWR _19340_/A sky130_fd_sc_hd__buf_2
XFILLER_52_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22350_ _22350_/A VGND VGND VPWR VPWR _23320_/D sky130_fd_sc_hd__buf_2
XFILLER_148_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21301_ _21299_/X _21293_/X _14359_/B _21300_/X VGND VGND VPWR VPWR _23932_/D sky130_fd_sc_hd__o22a_4
X_22281_ _22097_/X _22280_/X _12119_/B _22277_/X VGND VGND VPWR VPWR _22281_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14434__A _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19448__A2 _18576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24020_ _23668_/CLK _24020_/D VGND VGND VPWR VPWR _24020_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21255__A2 _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21232_ _21024_/X _21198_/A _23957_/Q _21195_/A VGND VGND VPWR VPWR _23957_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22651__A _22658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16131__A1 _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21163_ _20659_/X _21162_/X _15744_/B _21159_/X VGND VGND VPWR VPWR _24004_/D sky130_fd_sc_hd__o22a_4
XFILLER_172_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20114_ _20098_/X _20113_/Y _11642_/A _18624_/X _18666_/X VGND VGND VPWR VPWR _20114_/X
+ sky130_fd_sc_hd__o32a_4
X_21094_ _21086_/X VGND VGND VPWR VPWR _21094_/X sky130_fd_sc_hd__buf_2
XANTENNA__22204__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12889__A _12889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11793__A _11792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20045_ _20045_/A VGND VGND VPWR VPWR _24149_/D sky130_fd_sc_hd__inv_2
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18576__A _24212_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22507__A2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23804_ _23515_/CLK _23804_/D VGND VGND VPWR VPWR _14397_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17480__A _12574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21996_ _22010_/A VGND VGND VPWR VPWR _21996_/X sky130_fd_sc_hd__buf_2
XFILLER_2_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22098__A _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23735_ _23770_/CLK _23735_/D VGND VGND VPWR VPWR _23735_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _24408_/Q _20427_/A _24440_/Q _20282_/A VGND VGND VPWR VPWR _20947_/X sky130_fd_sc_hd__o22a_4
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14609__A _15415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23666_ _23852_/CLK _23666_/D VGND VGND VPWR VPWR _23666_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11680_/A VGND VGND VPWR VPWR _11681_/A sky130_fd_sc_hd__buf_2
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _20878_/A _20730_/B VGND VGND VPWR VPWR _20878_/X sky130_fd_sc_hd__or2_4
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22617_ _22452_/X _22615_/X _15868_/B _22612_/X VGND VGND VPWR VPWR _22617_/X sky130_fd_sc_hd__o22a_4
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17147__B1 _17145_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23597_ _23533_/CLK _21904_/X VGND VGND VPWR VPWR _16189_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22140__B1 _15474_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13350_ _13387_/A VGND VGND VPWR VPWR _13374_/A sky130_fd_sc_hd__buf_2
XANTENNA__21494__A2 _21492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22548_ _22548_/A VGND VGND VPWR VPWR _22548_/X sky130_fd_sc_hd__buf_2
XFILLER_6_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12301_ _12301_/A VGND VGND VPWR VPWR _12741_/A sky130_fd_sc_hd__buf_2
XFILLER_139_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11968__A _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13281_ _13321_/A _13281_/B _13280_/X VGND VGND VPWR VPWR _13281_/X sky130_fd_sc_hd__and3_4
X_22479_ _22478_/X _22474_/X _15253_/B _22469_/X VGND VGND VPWR VPWR _23256_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24216__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15020_ _13957_/A _24053_/Q VGND VGND VPWR VPWR _15020_/X sky130_fd_sc_hd__or2_4
X_12232_ _12704_/A _12229_/X _12232_/C VGND VGND VPWR VPWR _12247_/B sky130_fd_sc_hd__and3_4
XFILLER_108_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24218_ _24182_/CLK _24218_/D HRESETn VGND VGND VPWR VPWR _24218_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21246__A2 _21245_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22443__B2 _22433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12163_ _12127_/A _23123_/Q VGND VGND VPWR VPWR _12163_/X sky130_fd_sc_hd__or2_4
X_24149_ _24306_/CLK _24149_/D HRESETn VGND VGND VPWR VPWR _18250_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_155_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16971_ _16971_/A VGND VGND VPWR VPWR _17749_/A sky130_fd_sc_hd__inv_2
X_12094_ _12058_/A _23507_/Q VGND VGND VPWR VPWR _12094_/X sky130_fd_sc_hd__or2_4
XANTENNA__12799__A _13563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18710_ _18709_/A _18709_/B VGND VGND VPWR VPWR _18710_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15175__A _14301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15922_ _15391_/C _15921_/Y VGND VGND VPWR VPWR _15922_/Y sky130_fd_sc_hd__nor2_4
X_19690_ _19687_/A _19690_/B VGND VGND VPWR VPWR _19691_/A sky130_fd_sc_hd__or2_4
XFILLER_65_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18641_ _17621_/B _18639_/X _17792_/X _18640_/X VGND VGND VPWR VPWR _18641_/X sky130_fd_sc_hd__a211o_4
X_15853_ _13539_/A _15853_/B VGND VGND VPWR VPWR _15855_/B sky130_fd_sc_hd__or2_4
XFILLER_76_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14804_ _14823_/A _14721_/B VGND VGND VPWR VPWR _14805_/C sky130_fd_sc_hd__or2_4
X_18572_ _18499_/X _18569_/X _18527_/X _18571_/X VGND VGND VPWR VPWR _18572_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12996_ _12876_/A _23784_/Q VGND VGND VPWR VPWR _12997_/C sky130_fd_sc_hd__or2_4
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15784_ _15783_/X VGND VGND VPWR VPWR _15784_/X sky130_fd_sc_hd__buf_2
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17523_ _17522_/X VGND VGND VPWR VPWR _17523_/Y sky130_fd_sc_hd__inv_2
X_14735_ _15450_/A _14712_/X _14719_/X _14726_/X _14734_/X VGND VGND VPWR VPWR _14735_/X
+ sky130_fd_sc_hd__a32o_4
X_11947_ _11943_/X _11947_/B _11946_/X VGND VGND VPWR VPWR _11947_/X sky130_fd_sc_hd__and3_4
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14519__A _14519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21182__B2 _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13423__A _13427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17454_ _12097_/X _17481_/B VGND VGND VPWR VPWR _17454_/X sky130_fd_sc_hd__and2_4
X_14666_ _14675_/A _14584_/B VGND VGND VPWR VPWR _14667_/C sky130_fd_sc_hd__or2_4
X_11878_ _11878_/A VGND VGND VPWR VPWR _11879_/A sky130_fd_sc_hd__buf_2
XFILLER_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22736__A _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16405_ _16413_/A VGND VGND VPWR VPWR _16409_/A sky130_fd_sc_hd__buf_2
X_13617_ _13617_/A VGND VGND VPWR VPWR _15395_/A sky130_fd_sc_hd__buf_2
XFILLER_158_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17385_ _15786_/Y _17383_/A VGND VGND VPWR VPWR _17385_/X sky130_fd_sc_hd__and2_4
XANTENNA__17138__B1 _16383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14597_ _12477_/A _14597_/B VGND VGND VPWR VPWR _14597_/X sky130_fd_sc_hd__or2_4
X_19124_ _19126_/A _19021_/A _18957_/X VGND VGND VPWR VPWR _19124_/X sky130_fd_sc_hd__a21o_4
X_13548_ _13528_/A _13542_/X _13548_/C VGND VGND VPWR VPWR _13548_/X sky130_fd_sc_hd__or3_4
X_16336_ _11702_/X _16333_/X _16335_/X VGND VGND VPWR VPWR _16336_/X sky130_fd_sc_hd__and3_4
XFILLER_146_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22682__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11878__A _11878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16267_ _11904_/X _16267_/B VGND VGND VPWR VPWR _16267_/X sky130_fd_sc_hd__or2_4
X_19055_ _19053_/Y _19054_/Y _11530_/B VGND VGND VPWR VPWR _19055_/X sky130_fd_sc_hd__o21a_4
X_13479_ _12511_/A _23717_/Q VGND VGND VPWR VPWR _13481_/B sky130_fd_sc_hd__or2_4
XFILLER_145_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15218_ _11673_/A _15202_/X _15218_/C VGND VGND VPWR VPWR _15218_/X sky130_fd_sc_hd__or3_4
X_18006_ _17974_/X _17562_/A _18002_/X _17919_/X _18005_/Y VGND VGND VPWR VPWR _18007_/B
+ sky130_fd_sc_hd__a32o_4
X_16198_ _16214_/A _16190_/X _16197_/X VGND VGND VPWR VPWR _16198_/X sky130_fd_sc_hd__or3_4
XANTENNA__22434__B2 _22433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22471__A _22471_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15149_ _14988_/A _15149_/B VGND VGND VPWR VPWR _15151_/B sky130_fd_sc_hd__or2_4
XFILLER_5_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21087__A _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19957_ _19957_/A _19949_/X VGND VGND VPWR VPWR _19957_/X sky130_fd_sc_hd__or2_4
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18908_ _16381_/X _18906_/X _18983_/A _18907_/X VGND VGND VPWR VPWR _24399_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15085__A _12322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19888_ _19806_/A _19888_/B VGND VGND VPWR VPWR _19888_/X sky130_fd_sc_hd__or2_4
XANTENNA__23733__CLK _23904_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21815__A _21839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18839_ _18838_/X VGND VGND VPWR VPWR _18840_/A sky130_fd_sc_hd__buf_2
XFILLER_110_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18396__A _18064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15813__A _12875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21850_ _21280_/A VGND VGND VPWR VPWR _21850_/X sky130_fd_sc_hd__buf_2
X_20801_ _20801_/A VGND VGND VPWR VPWR _20801_/X sky130_fd_sc_hd__buf_2
XFILLER_24_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21781_ _21774_/A VGND VGND VPWR VPWR _21781_/X sky130_fd_sc_hd__buf_2
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14429__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23520_ _23649_/CLK _23520_/D VGND VGND VPWR VPWR _23520_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20732_ _20676_/X _20727_/Y _20730_/X _19066_/Y _20731_/X VGND VGND VPWR VPWR _20732_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23451_ _23772_/CLK _23451_/D VGND VGND VPWR VPWR _14503_/B sky130_fd_sc_hd__dfxtp_4
X_20663_ _11590_/X VGND VGND VPWR VPWR _20664_/A sky130_fd_sc_hd__buf_2
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22402_ _22167_/X _22397_/X _14929_/B _22366_/A VGND VGND VPWR VPWR _23286_/D sky130_fd_sc_hd__o22a_4
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23382_ _23095_/CLK _23382_/D VGND VGND VPWR VPWR _14961_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13987__B _24064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20594_ _24231_/Q _20534_/X _20593_/X VGND VGND VPWR VPWR _20595_/A sky130_fd_sc_hd__o21a_4
XFILLER_52_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20166__A IRQ[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22673__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22333_ _23337_/Q VGND VGND VPWR VPWR _22333_/X sky130_fd_sc_hd__buf_2
XFILLER_109_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17568__A1_N _16016_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19955__A _23083_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24376__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14164__A _14277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24199__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21228__A2 _21226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22264_ _22156_/X _22258_/X _14462_/B _22262_/X VGND VGND VPWR VPWR _23387_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24128__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12913__A1 _13453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24003_ _23939_/CLK _24003_/D VGND VGND VPWR VPWR _15804_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_151_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21215_ _20719_/X _21212_/X _15487_/B _21209_/X VGND VGND VPWR VPWR _21215_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_6_32_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_65_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17475__A _17145_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22195_ _22122_/X _22194_/X _23433_/Q _22191_/X VGND VGND VPWR VPWR _22195_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17906__C _17906_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21146_ _20395_/X _21141_/X _16406_/B _21145_/X VGND VGND VPWR VPWR _21146_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22728__A2 _22722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12412__A _12373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21077_ _20980_/X _21073_/X _15223_/B _21042_/A VGND VGND VPWR VPWR _21077_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21936__B1 _23573_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21400__A2 _21398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20028_ _18243_/X _20007_/X _20027_/Y _20018_/X VGND VGND VPWR VPWR _20028_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18801__B1 _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16819__A _11671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12850_ _12236_/A VGND VGND VPWR VPWR _12851_/A sky130_fd_sc_hd__buf_2
XANTENNA__15723__A _12783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11801_ _11833_/A _24020_/Q VGND VGND VPWR VPWR _11802_/C sky130_fd_sc_hd__or2_4
X_12781_ _12780_/X VGND VGND VPWR VPWR _12800_/A sky130_fd_sc_hd__buf_2
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _21869_/X _21974_/X _23548_/Q _21978_/X VGND VGND VPWR VPWR _21979_/X sky130_fd_sc_hd__o22a_4
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21164__B2 _21159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13243__A _13251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14520_ _14520_/A _24059_/Q VGND VGND VPWR VPWR _14521_/C sky130_fd_sc_hd__or2_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23718_ _23397_/CLK _21682_/X VGND VGND VPWR VPWR _23718_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11732_ _11705_/X _11718_/X _11731_/X VGND VGND VPWR VPWR _11732_/X sky130_fd_sc_hd__and3_4
XFILLER_109_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21661__A2_N _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _13046_/A _14428_/X _14435_/X _14442_/X _14450_/X VGND VGND VPWR VPWR _14451_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23649_ _23649_/CLK _23649_/D VGND VGND VPWR VPWR _23649_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11663_ _11663_/A VGND VGND VPWR VPWR _15377_/A sky130_fd_sc_hd__buf_2
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16554__A _12015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13375_/A _23814_/Q VGND VGND VPWR VPWR _13402_/X sky130_fd_sc_hd__or2_4
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ _17169_/X VGND VGND VPWR VPWR _17170_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14382_ _14511_/A _24060_/Q VGND VGND VPWR VPWR _14383_/C sky130_fd_sc_hd__or2_4
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21467__A2 _21462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22664__B2 _22662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11594_ _17038_/A _17038_/B VGND VGND VPWR VPWR _11647_/B sky130_fd_sc_hd__or2_4
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16121_ _16112_/A _23949_/Q VGND VGND VPWR VPWR _16123_/B sky130_fd_sc_hd__or2_4
Xclkbuf_7_114_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR _23650_/CLK sky130_fd_sc_hd__clkbuf_1
X_13333_ _13333_/A _23814_/Q VGND VGND VPWR VPWR _13333_/X sky130_fd_sc_hd__or2_4
XANTENNA__11698__A _11698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14074__A _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16052_ _16222_/A _16044_/X _16052_/C VGND VGND VPWR VPWR _16053_/C sky130_fd_sc_hd__and3_4
X_13264_ _13192_/X _13270_/A VGND VGND VPWR VPWR _13264_/X sky130_fd_sc_hd__or2_4
XFILLER_155_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22291__A _22291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20804__A _20422_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12306__B _23660_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15003_ _13990_/A _15003_/B VGND VGND VPWR VPWR _15005_/B sky130_fd_sc_hd__or2_4
X_12215_ _12228_/A VGND VGND VPWR VPWR _12696_/A sky130_fd_sc_hd__buf_2
XFILLER_124_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13195_ _13230_/A _23271_/Q VGND VGND VPWR VPWR _13195_/X sky130_fd_sc_hd__or2_4
XFILLER_124_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19811_ _19811_/A _19811_/B VGND VGND VPWR VPWR _19811_/X sky130_fd_sc_hd__and2_4
X_12146_ _11786_/X _12138_/X _12146_/C VGND VGND VPWR VPWR _12146_/X sky130_fd_sc_hd__and3_4
XFILLER_9_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19742_ _19742_/A _19777_/A VGND VGND VPWR VPWR _19742_/X sky130_fd_sc_hd__or2_4
XANTENNA__13418__A _13342_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16954_ _18190_/A VGND VGND VPWR VPWR _16954_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12077_ _11984_/X VGND VGND VPWR VPWR _12077_/X sky130_fd_sc_hd__buf_2
XANTENNA__12322__A _12322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15905_ _13514_/A _15905_/B _15904_/X VGND VGND VPWR VPWR _15909_/B sky130_fd_sc_hd__and3_4
X_19673_ _19576_/X _19666_/Y _19670_/Y _19467_/X _19672_/Y VGND VGND VPWR VPWR _19673_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_42_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16885_ _16527_/A _16836_/X _16527_/A _16836_/X VGND VGND VPWR VPWR _16885_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16729__A _16702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18624_ _18623_/Y VGND VGND VPWR VPWR _18624_/X sky130_fd_sc_hd__buf_2
XANTENNA__15633__A _13928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15836_ _12871_/A _15836_/B VGND VGND VPWR VPWR _15838_/B sky130_fd_sc_hd__or2_4
XFILLER_65_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18555_ _18111_/A _18533_/B _18553_/Y _18026_/X _18554_/Y VGND VGND VPWR VPWR _18555_/X
+ sky130_fd_sc_hd__a32o_4
X_12979_ _12979_/A _12979_/B _12979_/C VGND VGND VPWR VPWR _12979_/X sky130_fd_sc_hd__and3_4
X_15767_ _15741_/X _23108_/Q VGND VGND VPWR VPWR _15767_/X sky130_fd_sc_hd__or2_4
XANTENNA__17359__B1 _17358_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14249__A _12336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13153__A _12702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17506_ _17172_/X _18334_/B VGND VGND VPWR VPWR _18335_/B sky130_fd_sc_hd__or2_4
X_14718_ _12469_/A _14718_/B _14718_/C VGND VGND VPWR VPWR _14719_/C sky130_fd_sc_hd__and3_4
XFILLER_162_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18486_ _18440_/A _17365_/A VGND VGND VPWR VPWR _18486_/X sky130_fd_sc_hd__and2_4
X_15698_ _13145_/A _15698_/B VGND VGND VPWR VPWR _15699_/C sky130_fd_sc_hd__or2_4
XANTENNA__22466__A _20840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17437_ _17437_/A _17437_/B VGND VGND VPWR VPWR _17437_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__12992__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15385__A2 _15252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14649_ _14657_/A _14649_/B VGND VGND VPWR VPWR _14649_/X sky130_fd_sc_hd__or2_4
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21458__A2 _21455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17368_ _17360_/A _17367_/X VGND VGND VPWR VPWR _17368_/X sky130_fd_sc_hd__or2_4
XFILLER_158_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19520__A1 _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19520__B2 HRDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19107_ _18987_/A _19104_/Y _19105_/Y _19106_/X VGND VGND VPWR VPWR _19107_/X sky130_fd_sc_hd__o22a_4
X_16319_ _16314_/X _16316_/X _16319_/C VGND VGND VPWR VPWR _16319_/X sky130_fd_sc_hd__and3_4
X_17299_ _14767_/Y _17018_/X _17025_/Y _17298_/X VGND VGND VPWR VPWR _17300_/B sky130_fd_sc_hd__o22a_4
XANTENNA__24292__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19038_ _19024_/A VGND VGND VPWR VPWR _19038_/X sky130_fd_sc_hd__buf_2
XANTENNA__19494__B _19705_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12216__B _24044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20714__A _20714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_19_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14712__A _13589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21000_ _24246_/Q _20231_/A _20999_/X VGND VGND VPWR VPWR _21001_/B sky130_fd_sc_hd__o21a_4
XFILLER_138_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21630__A2 _21627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14431__B _14431_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12232__A _12704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22951_ _22947_/X _22949_/X _22951_/C VGND VGND VPWR VPWR _22951_/X sky130_fd_sc_hd__and3_4
XFILLER_28_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21394__B2 _21388_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21902_ _21909_/A VGND VGND VPWR VPWR _21902_/X sky130_fd_sc_hd__buf_2
X_22882_ _16016_/Y _22836_/X _22875_/X _22881_/X VGND VGND VPWR VPWR _22882_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21833_ _20509_/A VGND VGND VPWR VPWR _21833_/X sky130_fd_sc_hd__buf_2
XANTENNA__21146__B2 _21145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21764_ _21528_/X _21763_/X _23667_/Q _21760_/X VGND VGND VPWR VPWR _23667_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21697__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22376__A _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23503_ _23918_/CLK _22052_/X VGND VGND VPWR VPWR _16293_/B sky130_fd_sc_hd__dfxtp_4
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20715_ _20695_/X _20701_/Y _20712_/X _20713_/Y _20714_/X VGND VGND VPWR VPWR _20716_/B
+ sky130_fd_sc_hd__a32o_4
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24483_ _24134_/CLK _18452_/X HRESETn VGND VGND VPWR VPWR _24483_/Q sky130_fd_sc_hd__dfrtp_4
X_21695_ _21674_/A VGND VGND VPWR VPWR _21695_/X sky130_fd_sc_hd__buf_2
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21449__A2 _21448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23434_ _23404_/CLK _23434_/D VGND VGND VPWR VPWR _12731_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20646_ _24420_/Q _20645_/X _20159_/A _20471_/X VGND VGND VPWR VPWR _20646_/X sky130_fd_sc_hd__o22a_4
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22646__B2 _22641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23365_ _23397_/CLK _22300_/X VGND VGND VPWR VPWR _23365_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20577_ _20444_/X _19773_/X _20308_/A VGND VGND VPWR VPWR _20577_/X sky130_fd_sc_hd__a21o_4
XANTENNA__22823__B _15117_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22316_ _22158_/X _22315_/X _23354_/Q _22312_/X VGND VGND VPWR VPWR _22316_/X sky130_fd_sc_hd__o22a_4
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23296_ _23617_/CLK _23296_/D VGND VGND VPWR VPWR _23296_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20409__B1 _20638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16821__B _16821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23000__A _19438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22247_ _22127_/X _22244_/X _13240_/B _22241_/X VGND VGND VPWR VPWR _23399_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23071__A1 _19953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15718__A _15717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14622__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12000_ _16148_/A VGND VGND VPWR VPWR _12001_/A sky130_fd_sc_hd__buf_2
XFILLER_65_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21621__A2 _21620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22178_ _22171_/Y _22177_/X _22095_/X _22177_/X VGND VGND VPWR VPWR _22178_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21129_ _20980_/X _21125_/X _15134_/B _21086_/X VGND VGND VPWR VPWR _24023_/D sky130_fd_sc_hd__o22a_4
XFILLER_87_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21455__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13951_ _11853_/A VGND VGND VPWR VPWR _13951_/X sky130_fd_sc_hd__buf_2
XANTENNA__21385__B2 _21381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22582__B1 _15260_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11981__A _16568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12902_ _12514_/A _12902_/B VGND VGND VPWR VPWR _12903_/C sky130_fd_sc_hd__or2_4
Xclkbuf_7_39_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR _24080_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_86_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16670_ _16658_/A _23826_/Q VGND VGND VPWR VPWR _16670_/X sky130_fd_sc_hd__or2_4
X_13882_ _13882_/A VGND VGND VPWR VPWR _14348_/A sky130_fd_sc_hd__buf_2
XANTENNA__24404__CLK _23409_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12833_ _12833_/A _12833_/B VGND VGND VPWR VPWR _12835_/B sky130_fd_sc_hd__or2_4
X_15621_ _12337_/A _15619_/X _15621_/C VGND VGND VPWR VPWR _15625_/B sky130_fd_sc_hd__and3_4
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18764__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14069__A _11698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18340_ _17873_/X _18339_/X _17847_/A _17243_/X VGND VGND VPWR VPWR _18341_/A sky130_fd_sc_hd__o22a_4
X_12764_ _13562_/A _12759_/X _12764_/C VGND VGND VPWR VPWR _12764_/X sky130_fd_sc_hd__and3_4
X_15552_ _12239_/A _15552_/B VGND VGND VPWR VPWR _15552_/X sky130_fd_sc_hd__or2_4
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21190__A _21219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11715_ _11715_/A VGND VGND VPWR VPWR _16031_/A sky130_fd_sc_hd__buf_2
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _14511_/A _14503_/B VGND VGND VPWR VPWR _14503_/X sky130_fd_sc_hd__or2_4
X_15483_ _12630_/A _15479_/X _15482_/X VGND VGND VPWR VPWR _15483_/X sky130_fd_sc_hd__or3_4
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18271_ _17490_/A _18269_/X _18060_/X VGND VGND VPWR VPWR _18271_/Y sky130_fd_sc_hd__a21oi_4
X_12695_ _12691_/A _12693_/X _12695_/C VGND VGND VPWR VPWR _12699_/B sky130_fd_sc_hd__and3_4
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17222_ _17222_/A VGND VGND VPWR VPWR _18734_/B sky130_fd_sc_hd__inv_2
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14434_ _12428_/A _14432_/X _14433_/X VGND VGND VPWR VPWR _14435_/C sky130_fd_sc_hd__and3_4
X_11646_ _11646_/A VGND VGND VPWR VPWR _16936_/A sky130_fd_sc_hd__buf_2
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14516__B _14452_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ _13756_/A _14361_/X _14364_/X VGND VGND VPWR VPWR _14365_/X sky130_fd_sc_hd__or3_4
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17153_ _17153_/A VGND VGND VPWR VPWR _17153_/Y sky130_fd_sc_hd__inv_2
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11577_ _24463_/Q IRQ[26] VGND VGND VPWR VPWR _20186_/A sky130_fd_sc_hd__and2_4
XANTENNA__12317__A _11864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13316_ _13309_/A _13316_/B VGND VGND VPWR VPWR _13316_/X sky130_fd_sc_hd__or2_4
X_16104_ _15971_/A _16092_/X _16104_/C VGND VGND VPWR VPWR _16104_/X sky130_fd_sc_hd__or3_4
X_17084_ _18517_/A VGND VGND VPWR VPWR _18220_/A sky130_fd_sc_hd__buf_2
XANTENNA__16867__A2 _16866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14296_ _14296_/A _14360_/B VGND VGND VPWR VPWR _14297_/C sky130_fd_sc_hd__or2_4
XANTENNA__20534__A _20895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16035_ _16035_/A _16032_/X _16034_/X VGND VGND VPWR VPWR _16036_/C sky130_fd_sc_hd__and3_4
X_13247_ _13235_/A _13247_/B _13246_/X VGND VGND VPWR VPWR _13247_/X sky130_fd_sc_hd__and3_4
XANTENNA__19409__A2_N _18278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13178_ _13324_/A _13176_/X _13177_/X VGND VGND VPWR VPWR _13182_/B sky130_fd_sc_hd__and3_4
XFILLER_69_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14251__B _23487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13148__A _13303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20820__B1 _24094_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12129_ _12129_/A _12129_/B _12128_/X VGND VGND VPWR VPWR _12130_/C sky130_fd_sc_hd__and3_4
X_17986_ _17229_/X VGND VGND VPWR VPWR _17986_/X sky130_fd_sc_hd__buf_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19725_ _19725_/A _19712_/X VGND VGND VPWR VPWR _19725_/X sky130_fd_sc_hd__or2_4
X_16937_ _17017_/A _16936_/X _11592_/X _17087_/A VGND VGND VPWR VPWR _16937_/X sky130_fd_sc_hd__or4_4
XANTENNA__20179__A2 IRQ[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16459__A _11727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22573__B1 _23199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19656_ _19509_/X _19655_/X VGND VGND VPWR VPWR _19656_/X sky130_fd_sc_hd__and2_4
XFILLER_38_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16868_ _15386_/X _14848_/Y _15387_/B VGND VGND VPWR VPWR _16868_/X sky130_fd_sc_hd__o21a_4
X_18607_ _18483_/A _17307_/X VGND VGND VPWR VPWR _18607_/Y sky130_fd_sc_hd__nor2_4
X_15819_ _12847_/A _15819_/B VGND VGND VPWR VPWR _15819_/X sky130_fd_sc_hd__or2_4
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19587_ _19493_/A _19581_/A _19643_/A VGND VGND VPWR VPWR _19588_/C sky130_fd_sc_hd__or3_4
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21128__B2 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16799_ _16811_/A _16799_/B VGND VGND VPWR VPWR _16799_/X sky130_fd_sc_hd__or2_4
X_18538_ _18538_/A VGND VGND VPWR VPWR _18538_/X sky130_fd_sc_hd__buf_2
XANTENNA__21679__A2 _21677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18469_ _18413_/X _17362_/X _18466_/X _18467_/X _18468_/Y VGND VGND VPWR VPWR _18469_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16194__A _11727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14707__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13611__A _14292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20500_ _20754_/A _20499_/X _24331_/Q _20761_/A VGND VGND VPWR VPWR _20501_/B sky130_fd_sc_hd__o22a_4
X_21480_ _21247_/X _21478_/X _23826_/Q _21475_/X VGND VGND VPWR VPWR _23826_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23921__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22628__B2 _22626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22924__A _23078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20431_ _20425_/X _20430_/X _24302_/Q _20349_/X VGND VGND VPWR VPWR _20431_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12227__A _11880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16922__A _16915_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23150_ _23918_/CLK _23150_/D VGND VGND VPWR VPWR _15988_/B sky130_fd_sc_hd__dfxtp_4
X_20362_ _20302_/X _20361_/X _24114_/Q _20225_/X VGND VGND VPWR VPWR _24114_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20444__A _18779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22101_ _20360_/A VGND VGND VPWR VPWR _22101_/X sky130_fd_sc_hd__buf_2
XANTENNA__15538__A _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23081_ _19953_/A _19328_/Y _22742_/A _23080_/X VGND VGND VPWR VPWR _23081_/X sky130_fd_sc_hd__a211o_4
XANTENNA__14442__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20293_ _19975_/X _20260_/X _20262_/X _20292_/X VGND VGND VPWR VPWR _20293_/X sky130_fd_sc_hd__a211o_4
X_22032_ _21874_/X _22031_/X _23514_/Q _22028_/X VGND VGND VPWR VPWR _23514_/D sky130_fd_sc_hd__o22a_4
XFILLER_87_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14161__B _23231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23983_ _23983_/CLK _23983_/D VGND VGND VPWR VPWR _16280_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12897__A _12874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16369__A _16362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21367__B2 _21331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15273__A _13788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22934_ _17741_/A _16973_/X _17738_/X VGND VGND VPWR VPWR _22934_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19980__A1 _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22865_ _22865_/A VGND VGND VPWR VPWR HWDATA[20] sky130_fd_sc_hd__inv_2
XANTENNA__21119__B2 _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21816_ _21813_/X _21815_/X _23635_/Q _21810_/X VGND VGND VPWR VPWR _23635_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22867__A1 _12753_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22796_ _22794_/Y _22791_/X _24117_/D _22795_/Y VGND VGND VPWR VPWR _22796_/X sky130_fd_sc_hd__a211o_4
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21747_ _21587_/X _21741_/X _14436_/B _21745_/X VGND VGND VPWR VPWR _23675_/D sky130_fd_sc_hd__o22a_4
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _12867_/A _12608_/B VGND VGND VPWR VPWR _12489_/B sky130_fd_sc_hd__or2_4
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24466_ _23379_/CLK _18793_/X HRESETn VGND VGND VPWR VPWR _24466_/Q sky130_fd_sc_hd__dfrtp_4
X_21678_ _21553_/X _21677_/X _23721_/Q _21674_/X VGND VGND VPWR VPWR _21678_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24143__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23417_ _23772_/CLK _23417_/D VGND VGND VPWR VPWR _23417_/Q sky130_fd_sc_hd__dfxtp_4
X_20629_ _24261_/Q _20443_/X _20628_/X VGND VGND VPWR VPWR _20629_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19496__B1 HRDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24397_ _24397_/CLK _24397_/D HRESETn VGND VGND VPWR VPWR _24397_/Q sky130_fd_sc_hd__dfstp_4
X_14150_ _11869_/A _14150_/B _14149_/X VGND VGND VPWR VPWR _14150_/X sky130_fd_sc_hd__or3_4
XFILLER_138_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23348_ _23668_/CLK _23348_/D VGND VGND VPWR VPWR _11804_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21842__A2 _21839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13101_ _13094_/A _13025_/B VGND VGND VPWR VPWR _13101_/X sky130_fd_sc_hd__or2_4
XFILLER_125_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15448__A _12251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19380__A2_N _18741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14081_ _11753_/A _14081_/B _14080_/X VGND VGND VPWR VPWR _14082_/C sky130_fd_sc_hd__or3_4
X_23279_ _23760_/CLK _22424_/X VGND VGND VPWR VPWR _16247_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14352__A _13697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13032_ _12510_/A _23496_/Q VGND VGND VPWR VPWR _13034_/B sky130_fd_sc_hd__or2_4
XFILLER_65_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14071__B _23712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20802__B1 _24095_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17840_ _17922_/A _17835_/X _17836_/X _17839_/X VGND VGND VPWR VPWR _17840_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17771_ _17693_/X VGND VGND VPWR VPWR _17771_/Y sky130_fd_sc_hd__inv_2
X_14983_ _14983_/A VGND VGND VPWR VPWR _14984_/A sky130_fd_sc_hd__inv_2
XFILLER_75_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21358__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19510_ _19509_/X VGND VGND VPWR VPWR _19510_/X sky130_fd_sc_hd__buf_2
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15183__A _13853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16722_ _16695_/A _16722_/B _16722_/C VGND VGND VPWR VPWR _16726_/B sky130_fd_sc_hd__and3_4
X_13934_ _13720_/A _13932_/X _13933_/X VGND VGND VPWR VPWR _13934_/X sky130_fd_sc_hd__and3_4
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21913__A _21906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19441_ _19719_/A VGND VGND VPWR VPWR _19441_/X sky130_fd_sc_hd__buf_2
XANTENNA__13048__B1 _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16653_ _16053_/A _16630_/X _16652_/X VGND VGND VPWR VPWR _16685_/B sky130_fd_sc_hd__or3_4
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13865_ _13865_/A VGND VGND VPWR VPWR _14335_/A sky130_fd_sc_hd__buf_2
XFILLER_16_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15911__A _12676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15604_ _13866_/A VGND VGND VPWR VPWR _15641_/A sky130_fd_sc_hd__buf_2
X_12816_ _12759_/A _12816_/B VGND VGND VPWR VPWR _12816_/X sky130_fd_sc_hd__or2_4
X_19372_ _19372_/A VGND VGND VPWR VPWR _19372_/X sky130_fd_sc_hd__buf_2
XANTENNA__22858__A1 _17518_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23944__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16584_ _16561_/A _16580_/X _16584_/C VGND VGND VPWR VPWR _16584_/X sky130_fd_sc_hd__or3_4
X_13796_ _14304_/A _13796_/B VGND VGND VPWR VPWR _13801_/B sky130_fd_sc_hd__or2_4
X_18323_ _17527_/D _18322_/X VGND VGND VPWR VPWR _18323_/X sky130_fd_sc_hd__or2_4
XFILLER_128_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15535_ _15442_/A _15535_/B _15534_/X VGND VGND VPWR VPWR _15535_/X sky130_fd_sc_hd__or3_4
XFILLER_31_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12747_ _12747_/A _12747_/B VGND VGND VPWR VPWR _12747_/X sky130_fd_sc_hd__or2_4
XANTENNA__20333__A2 _20305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13431__A _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18254_ _23020_/B _18253_/Y _17681_/A _18253_/A VGND VGND VPWR VPWR _18254_/X sky130_fd_sc_hd__o22a_4
X_15466_ _12592_/A _15466_/B VGND VGND VPWR VPWR _15467_/C sky130_fd_sc_hd__or2_4
X_12678_ _12677_/X VGND VGND VPWR VPWR _12678_/X sky130_fd_sc_hd__buf_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17205_ _13270_/X _17197_/X _17170_/Y _17198_/X VGND VGND VPWR VPWR _17205_/X sky130_fd_sc_hd__o22a_4
X_11629_ _11629_/A VGND VGND VPWR VPWR _11630_/A sky130_fd_sc_hd__buf_2
X_14417_ _14415_/Y _14417_/B VGND VGND VPWR VPWR _14417_/X sky130_fd_sc_hd__or2_4
X_18185_ _18020_/X _18179_/X _18065_/X _18184_/X VGND VGND VPWR VPWR _18185_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19487__B1 HRDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22086__A2 _22081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15397_ _15401_/A _15395_/X _15397_/C VGND VGND VPWR VPWR _15398_/C sky130_fd_sc_hd__and3_4
XANTENNA__16742__A _16742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17136_ _17817_/A _17126_/X _17128_/X _17135_/X VGND VGND VPWR VPWR _17136_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21294__B1 _23935_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14348_ _14348_/A VGND VGND VPWR VPWR _14522_/A sky130_fd_sc_hd__buf_2
XANTENNA__11886__A _11886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17067_ _18782_/B _11595_/A _11648_/X VGND VGND VPWR VPWR _17067_/X sky130_fd_sc_hd__a21o_4
X_14279_ _12454_/A _23772_/Q VGND VGND VPWR VPWR _14280_/C sky130_fd_sc_hd__or2_4
XFILLER_171_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16018_ _16033_/A _15940_/B VGND VGND VPWR VPWR _16018_/X sky130_fd_sc_hd__or2_4
XANTENNA__15077__B _23989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21597__B2 _21524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17969_ _18674_/A VGND VGND VPWR VPWR _18407_/A sky130_fd_sc_hd__buf_2
XFILLER_100_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21349__B2 _21345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19708_ _19546_/X _19883_/A VGND VGND VPWR VPWR _19889_/C sky130_fd_sc_hd__or2_4
XANTENNA__12510__A _12510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20980_ _21311_/A VGND VGND VPWR VPWR _20980_/X sky130_fd_sc_hd__buf_2
XFILLER_38_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19639_ _20776_/A _19573_/X _19637_/X _19638_/X VGND VGND VPWR VPWR _19639_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_22_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR _24471_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_85_0_HCLK clkbuf_6_42_0_HCLK/X VGND VGND VPWR VPWR _23416_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15821__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22650_ _22423_/X _22644_/X _16286_/B _22648_/X VGND VGND VPWR VPWR _23151_/D sky130_fd_sc_hd__o22a_4
XFILLER_129_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21601_ _21600_/X _21542_/A _23765_/Q _21524_/X VGND VGND VPWR VPWR _23765_/D sky130_fd_sc_hd__o22a_4
XFILLER_90_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22581_ _22476_/X _22579_/X _14713_/B _22576_/X VGND VGND VPWR VPWR _23193_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14437__A _13010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24320_ _24292_/CLK _19202_/X HRESETn VGND VGND VPWR VPWR _19141_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21532_ _21532_/A VGND VGND VPWR VPWR _21532_/X sky130_fd_sc_hd__buf_2
XFILLER_166_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24251_ _24248_/CLK _24251_/D HRESETn VGND VGND VPWR VPWR _24251_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22077__A2 _22074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19478__B1 HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21463_ _21304_/X _21462_/X _14591_/B _21459_/X VGND VGND VPWR VPWR _23834_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16652__A _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23202_ _23204_/CLK _23202_/D VGND VGND VPWR VPWR _15399_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20414_ _24239_/Q _20304_/X _20413_/X VGND VGND VPWR VPWR _20415_/A sky130_fd_sc_hd__o21a_4
XFILLER_147_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24182_ _24182_/CLK _19905_/Y HRESETn VGND VGND VPWR VPWR _17038_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_162_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21394_ _21273_/X _21391_/X _23879_/Q _21388_/X VGND VGND VPWR VPWR _23879_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11796__A _16635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23133_ _23229_/CLK _22675_/X VGND VGND VPWR VPWR _13838_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15268__A _14269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20345_ _24434_/Q _18837_/B _24466_/Q _20282_/X VGND VGND VPWR VPWR _20345_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14172__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23064_ _19924_/A _24159_/Q _16997_/B _17957_/X _22930_/A VGND VGND VPWR VPWR _23064_/X
+ sky130_fd_sc_hd__o32a_4
X_20276_ _20275_/X VGND VGND VPWR VPWR _20470_/A sky130_fd_sc_hd__buf_2
XFILLER_115_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12404__B _12314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21588__B2 _21585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22015_ _21845_/X _22010_/X _13274_/B _22014_/X VGND VGND VPWR VPWR _22015_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17483__A _17482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14900__A _14897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16099__A _12561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22001__A2 _21996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12420__A _12320_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11980_ _11951_/A _11978_/X _11979_/X VGND VGND VPWR VPWR _11980_/X sky130_fd_sc_hd__and3_4
X_23966_ _23880_/CLK _21221_/X VGND VGND VPWR VPWR _23966_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22917_ _22916_/X VGND VGND VPWR VPWR HADDR[2] sky130_fd_sc_hd__inv_2
XFILLER_17_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23897_ _23294_/CLK _23897_/D VGND VGND VPWR VPWR _14736_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15731__A _12778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13650_ _15420_/A _13649_/X VGND VGND VPWR VPWR _13650_/X sky130_fd_sc_hd__and2_4
X_22848_ _22800_/Y VGND VGND VPWR VPWR _22848_/X sky130_fd_sc_hd__buf_2
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24324__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _12927_/A VGND VGND VPWR VPWR _12644_/A sky130_fd_sc_hd__buf_2
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13581_ _13581_/A VGND VGND VPWR VPWR _13582_/B sky130_fd_sc_hd__inv_2
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ _22753_/Y _22778_/B VGND VGND VPWR VPWR _22781_/B sky130_fd_sc_hd__or2_4
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13251__A _13251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21512__B2 _21510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12532_ _12875_/A VGND VGND VPWR VPWR _12891_/A sky130_fd_sc_hd__buf_2
X_15320_ _15372_/A _15318_/X _15320_/C VGND VGND VPWR VPWR _15321_/C sky130_fd_sc_hd__and3_4
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12463_ _12863_/A _12599_/B VGND VGND VPWR VPWR _12465_/B sky130_fd_sc_hd__or2_4
XANTENNA__22068__A2 _22067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15251_ _15251_/A VGND VGND VPWR VPWR _15252_/A sky130_fd_sc_hd__inv_2
XFILLER_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24449_ _23475_/CLK _24449_/D HRESETn VGND VGND VPWR VPWR _24449_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16562__A _11960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14202_ _14630_/A _14202_/B _14201_/X VGND VGND VPWR VPWR _14203_/C sky130_fd_sc_hd__or3_4
X_15182_ _15029_/A _15178_/X _15182_/C VGND VGND VPWR VPWR _15182_/X sky130_fd_sc_hd__or3_4
X_12394_ _12339_/X _12394_/B _12394_/C VGND VGND VPWR VPWR _12394_/X sky130_fd_sc_hd__and3_4
X_14133_ _14133_/A _14129_/X _14132_/X VGND VGND VPWR VPWR _14133_/X sky130_fd_sc_hd__or3_4
XANTENNA__15178__A _13954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19990_ _18670_/X _17655_/A _19956_/X _19989_/X VGND VGND VPWR VPWR _19991_/A sky130_fd_sc_hd__o22a_4
XANTENNA__14082__A _11680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18941_ _15118_/X _18897_/A _20990_/A _18900_/A VGND VGND VPWR VPWR _24374_/D sky130_fd_sc_hd__o22a_4
X_14064_ _11736_/A _14062_/X _14063_/X VGND VGND VPWR VPWR _14065_/C sky130_fd_sc_hd__and3_4
XANTENNA__23497__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12314__B _12314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21579__B2 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13015_ _12461_/A _13015_/B _13014_/X VGND VGND VPWR VPWR _13016_/B sky130_fd_sc_hd__or3_4
XANTENNA__22240__A2 _22237_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19641__B1 HRDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18872_ _17161_/X _18870_/X _24416_/Q _18871_/X VGND VGND VPWR VPWR _18872_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14810__A _14682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17823_ _17823_/A VGND VGND VPWR VPWR _17823_/X sky130_fd_sc_hd__buf_2
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22528__B1 _14469_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13426__A _13455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17754_ _17005_/A _17336_/X _17752_/X _17753_/X VGND VGND VPWR VPWR _18721_/A sky130_fd_sc_hd__o22a_4
X_14966_ _14973_/A _14902_/B VGND VGND VPWR VPWR _14966_/X sky130_fd_sc_hd__or2_4
XFILLER_48_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16705_ _16724_/A _24017_/Q VGND VGND VPWR VPWR _16706_/C sky130_fd_sc_hd__or2_4
XFILLER_130_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19944__B2 _20598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13917_ _13877_/A VGND VGND VPWR VPWR _13937_/A sky130_fd_sc_hd__buf_2
X_17685_ _16988_/A VGND VGND VPWR VPWR _17686_/A sky130_fd_sc_hd__buf_2
XFILLER_75_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20554__A2 _20536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14897_ _13591_/A VGND VGND VPWR VPWR _14897_/X sky130_fd_sc_hd__buf_2
XANTENNA__21751__A1 _21594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21751__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19424_ _19421_/X _18580_/X _19421_/X _24221_/Q VGND VGND VPWR VPWR _19424_/X sky130_fd_sc_hd__a2bb2o_4
X_16636_ _11768_/X VGND VGND VPWR VPWR _16788_/A sky130_fd_sc_hd__buf_2
X_13848_ _13675_/A _13848_/B VGND VGND VPWR VPWR _13850_/B sky130_fd_sc_hd__or2_4
XFILLER_90_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24122__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19355_ _19354_/X _18353_/X _19354_/X _20608_/A VGND VGND VPWR VPWR _24262_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16567_ _11951_/A _16567_/B _16567_/C VGND VGND VPWR VPWR _16568_/C sky130_fd_sc_hd__and3_4
X_13779_ _12576_/A _13771_/X _13778_/X VGND VGND VPWR VPWR _13779_/X sky130_fd_sc_hd__and3_4
XANTENNA__14257__A _13882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13161__A _13277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18306_ _18244_/X _18305_/X _20036_/A _18244_/X VGND VGND VPWR VPWR _24488_/D sky130_fd_sc_hd__a2bb2o_4
X_15518_ _15453_/Y _15517_/X VGND VGND VPWR VPWR _15518_/X sky130_fd_sc_hd__and2_4
X_19286_ _24294_/Q _19243_/B _19285_/Y VGND VGND VPWR VPWR _24294_/D sky130_fd_sc_hd__o21a_4
X_16498_ _16491_/A _16429_/B VGND VGND VPWR VPWR _16498_/X sky130_fd_sc_hd__or2_4
XANTENNA__22474__A _22462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17183__A1 _17132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18237_ _17490_/B _18235_/X _18176_/X VGND VGND VPWR VPWR _18237_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__22059__A2 _22053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15449_ _15449_/A _15445_/X _15448_/X VGND VGND VPWR VPWR _15449_/X sky130_fd_sc_hd__or3_4
XFILLER_15_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18168_ _18168_/A VGND VGND VPWR VPWR _18168_/X sky130_fd_sc_hd__buf_2
XANTENNA__14704__B _14701_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17119_ _17164_/A VGND VGND VPWR VPWR _17119_/X sky130_fd_sc_hd__buf_2
XFILLER_144_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19783__A HRDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18683__A1 _18032_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18683__B2 _18682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18099_ _18099_/A _18098_/X VGND VGND VPWR VPWR _18099_/X sky130_fd_sc_hd__or2_4
XFILLER_143_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20130_ _19952_/Y _20129_/X _24473_/Q _19979_/X VGND VGND VPWR VPWR _20130_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20722__A _20364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18435__A1 _18022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15816__A _12858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20061_ _18451_/X _20055_/X _20060_/Y _20042_/X VGND VGND VPWR VPWR _20061_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22231__A2 _22230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14720__A _13666_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23820_ _23852_/CLK _23820_/D VGND VGND VPWR VPWR _12399_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23751_ _23750_/CLK _23751_/D VGND VGND VPWR VPWR _23751_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19935__B2 _21007_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20963_ _20864_/X _20961_/X _20962_/X HRDATA[10] _20869_/X VGND VGND VPWR VPWR _20963_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16749__A1 _11984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16647__A _16647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22702_ _20441_/A _22701_/X _23118_/Q _22698_/X VGND VGND VPWR VPWR _22702_/X sky130_fd_sc_hd__o22a_4
XPHY_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21742__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23682_ _23650_/CLK _21737_/X VGND VGND VPWR VPWR _15477_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20894_ _20772_/A VGND VGND VPWR VPWR _20894_/X sky130_fd_sc_hd__buf_2
XPHY_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15421__A1 _14480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22633_ _22480_/X _22629_/X _15149_/B _22598_/A VGND VGND VPWR VPWR _23159_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13071__A _13103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22564_ _22447_/X _22558_/X _13500_/B _22562_/X VGND VGND VPWR VPWR _23205_/D sky130_fd_sc_hd__o22a_4
XFILLER_16_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24303_ _24306_/CLK _24303_/D HRESETn VGND VGND VPWR VPWR _19252_/A sky130_fd_sc_hd__dfrtp_4
X_21515_ _21307_/X _21513_/X _14758_/B _21510_/X VGND VGND VPWR VPWR _21515_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16382__A _16381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22495_ _22412_/X _22494_/X _12173_/B _22491_/X VGND VGND VPWR VPWR _23251_/D sky130_fd_sc_hd__o22a_4
X_24234_ _24271_/CLK _24234_/D HRESETn VGND VGND VPWR VPWR _24234_/Q sky130_fd_sc_hd__dfrtp_4
X_21446_ _21275_/X _21441_/X _23846_/Q _21445_/X VGND VGND VPWR VPWR _21446_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24165_ _23991_/CLK _24165_/D HRESETn VGND VGND VPWR VPWR _24165_/Q sky130_fd_sc_hd__dfrtp_4
X_21377_ _21391_/A VGND VGND VPWR VPWR _21377_/X sky130_fd_sc_hd__buf_2
XANTENNA__19871__B1 _21081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12415__A _15887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23116_ _23852_/CLK _23116_/D VGND VGND VPWR VPWR _12398_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20328_ _20754_/A _20326_/X _24339_/Q _20761_/A VGND VGND VPWR VPWR _20329_/B sky130_fd_sc_hd__o22a_4
X_24096_ _24096_/CLK _24096_/D VGND VGND VPWR VPWR _24096_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20632__A _20632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15726__A _12758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23047_ _23047_/A VGND VGND VPWR VPWR HADDR[24] sky130_fd_sc_hd__inv_2
X_20259_ _20259_/A VGND VGND VPWR VPWR _20260_/A sky130_fd_sc_hd__buf_2
XFILLER_7_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14820_ _14820_/A _14744_/B VGND VGND VPWR VPWR _14821_/C sky130_fd_sc_hd__or2_4
XANTENNA__12150__A _11762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24145__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14751_ _15447_/A _14751_/B VGND VGND VPWR VPWR _14751_/X sky130_fd_sc_hd__or2_4
X_23949_ _24077_/CLK _21260_/X VGND VGND VPWR VPWR _23949_/Q sky130_fd_sc_hd__dfxtp_4
X_11963_ _11963_/A _11961_/X _11962_/X VGND VGND VPWR VPWR _11964_/C sky130_fd_sc_hd__and3_4
XANTENNA__16557__A _12001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20536__A2 _20917_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21733__B2 _21731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13702_ _14541_/A _13702_/B VGND VGND VPWR VPWR _13702_/X sky130_fd_sc_hd__or2_4
X_17470_ _18165_/B VGND VGND VPWR VPWR _17490_/B sky130_fd_sc_hd__inv_2
X_11894_ _13792_/A VGND VGND VPWR VPWR _12194_/A sky130_fd_sc_hd__inv_2
X_14682_ _14682_/A _14682_/B _14682_/C VGND VGND VPWR VPWR _14699_/B sky130_fd_sc_hd__and3_4
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16421_ _16007_/X _16421_/B VGND VGND VPWR VPWR _16421_/X sky130_fd_sc_hd__or2_4
X_13633_ _11879_/A _13629_/X _13633_/C VGND VGND VPWR VPWR _13641_/B sky130_fd_sc_hd__and3_4
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22289__A2 _22287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14077__A _11736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24295__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19140_ _24319_/Q _19205_/A VGND VGND VPWR VPWR _19141_/B sky130_fd_sc_hd__and2_4
X_16352_ _11702_/X _16350_/X _16351_/X VGND VGND VPWR VPWR _16352_/X sky130_fd_sc_hd__and3_4
X_13564_ _13564_/A _13564_/B _13564_/C VGND VGND VPWR VPWR _13565_/C sky130_fd_sc_hd__and3_4
XFILLER_9_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22294__A _22294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15303_ _14301_/A _15303_/B _15302_/X VGND VGND VPWR VPWR _15303_/X sky130_fd_sc_hd__or3_4
X_12515_ _12515_/A _12515_/B _12515_/C VGND VGND VPWR VPWR _12516_/C sky130_fd_sc_hd__and3_4
X_19071_ _24384_/Q VGND VGND VPWR VPWR _19071_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13495_ _12949_/A VGND VGND VPWR VPWR _13496_/A sky130_fd_sc_hd__buf_2
X_16283_ _16287_/A _16283_/B VGND VGND VPWR VPWR _16283_/X sky130_fd_sc_hd__or2_4
XANTENNA__16292__A _16159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18022_ _18148_/A VGND VGND VPWR VPWR _18022_/X sky130_fd_sc_hd__buf_2
X_12446_ _13011_/A VGND VGND VPWR VPWR _12877_/A sky130_fd_sc_hd__buf_2
X_15234_ _15196_/X _15176_/B VGND VGND VPWR VPWR _15234_/X sky130_fd_sc_hd__or2_4
XANTENNA__14524__B _14460_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12377_ _12339_/X _12377_/B _12377_/C VGND VGND VPWR VPWR _12378_/C sky130_fd_sc_hd__and3_4
X_15165_ _14574_/A _15165_/B VGND VGND VPWR VPWR _15165_/X sky130_fd_sc_hd__or2_4
XANTENNA__19862__B1 _19788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14116_ _14165_/A VGND VGND VPWR VPWR _14154_/A sky130_fd_sc_hd__buf_2
XANTENNA__21638__A _21624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19973_ _19973_/A _19972_/X VGND VGND VPWR VPWR _19973_/X sky130_fd_sc_hd__or2_4
X_15096_ _15096_/A _23413_/Q VGND VGND VPWR VPWR _15097_/C sky130_fd_sc_hd__or2_4
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18924_ _15916_/X _18920_/X _24387_/Q _18921_/X VGND VGND VPWR VPWR _18924_/X sky130_fd_sc_hd__o22a_4
X_14047_ _11736_/A _14045_/X _14047_/C VGND VGND VPWR VPWR _14048_/C sky130_fd_sc_hd__and3_4
XANTENNA__22213__A2 _22208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15355__B _23128_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18855_ _12678_/X _18849_/X _24427_/Q _18850_/X VGND VGND VPWR VPWR _24427_/D sky130_fd_sc_hd__o22a_4
XFILLER_95_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13156__A _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17806_ _17805_/X VGND VGND VPWR VPWR _17807_/A sky130_fd_sc_hd__buf_2
XANTENNA__21972__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18786_ _18786_/A VGND VGND VPWR VPWR _18796_/A sky130_fd_sc_hd__buf_2
X_15998_ _13474_/A VGND VGND VPWR VPWR _15998_/X sky130_fd_sc_hd__buf_2
XANTENNA__19917__A1 _19906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22469__A _22433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21373__A _21388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17737_ _17737_/A _17735_/A VGND VGND VPWR VPWR _17737_/X sky130_fd_sc_hd__or2_4
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14949_ _14663_/A _14941_/X _14948_/X VGND VGND VPWR VPWR _14949_/X sky130_fd_sc_hd__and3_4
XANTENNA__12995__A _12875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20527__A2 _20513_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15371__A _13704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17668_ _17667_/X VGND VGND VPWR VPWR _17668_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19407_ _19406_/X VGND VGND VPWR VPWR _19407_/X sky130_fd_sc_hd__buf_2
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16619_ _16675_/A _16612_/X _16618_/X VGND VGND VPWR VPWR _16619_/X sky130_fd_sc_hd__or3_4
XFILLER_91_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17599_ _17485_/X _17598_/Y _17478_/B _17487_/X VGND VGND VPWR VPWR _17599_/X sky130_fd_sc_hd__a211o_4
X_19338_ _19335_/X _17960_/X _19335_/X _20373_/A VGND VGND VPWR VPWR _24273_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19269_ _19252_/B VGND VGND VPWR VPWR _19269_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14715__A _14297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21300_ _21264_/A VGND VGND VPWR VPWR _21300_/X sky130_fd_sc_hd__buf_2
X_22280_ _22294_/A VGND VGND VPWR VPWR _22280_/X sky130_fd_sc_hd__buf_2
XFILLER_116_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21231_ _21004_/X _21226_/X _23958_/Q _21195_/A VGND VGND VPWR VPWR _21231_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12235__A _13687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21162_ _21155_/A VGND VGND VPWR VPWR _21162_/X sky130_fd_sc_hd__buf_2
XFILLER_137_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20113_ _20112_/X VGND VGND VPWR VPWR _20113_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22204__A2 _22201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15546__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21093_ _20378_/X _21090_/X _24049_/Q _21087_/X VGND VGND VPWR VPWR _24049_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14450__A _14450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20044_ _20040_/X _17688_/A _20022_/X _20043_/X VGND VGND VPWR VPWR _20045_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24168__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21963__B2 _21957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18576__B _18576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23803_ _23515_/CLK _23803_/D VGND VGND VPWR VPWR _14474_/B sky130_fd_sc_hd__dfxtp_4
X_21995_ _21991_/A VGND VGND VPWR VPWR _22010_/A sky130_fd_sc_hd__buf_2
XANTENNA__16377__A _16370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24399__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21715__B2 _21710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15281__A _15281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _20943_/X _20945_/X _20262_/X VGND VGND VPWR VPWR _20946_/Y sky130_fd_sc_hd__o21ai_4
X_23734_ _23194_/CLK _23734_/D VGND VGND VPWR VPWR _23734_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_55_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23665_ _23761_/CLK _23665_/D VGND VGND VPWR VPWR _23665_/Q sky130_fd_sc_hd__dfxtp_4
X_20877_ _24443_/Q VGND VGND VPWR VPWR _20878_/A sky130_fd_sc_hd__inv_2
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22826__B _17327_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22616_ _22449_/X _22615_/X _15737_/B _22612_/X VGND VGND VPWR VPWR _22616_/X sky130_fd_sc_hd__o22a_4
X_23596_ _23500_/CLK _23596_/D VGND VGND VPWR VPWR _23596_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17147__A1 _13947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22140__B2 _22130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23003__A _18350_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22547_ _22418_/X _22544_/X _16761_/B _22541_/X VGND VGND VPWR VPWR _23217_/D sky130_fd_sc_hd__o22a_4
X_12300_ _12300_/A VGND VGND VPWR VPWR _12301_/A sky130_fd_sc_hd__buf_2
XFILLER_33_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13280_ _13313_/A _13280_/B VGND VGND VPWR VPWR _13280_/X sky130_fd_sc_hd__or2_4
X_22478_ _20958_/A VGND VGND VPWR VPWR _22478_/X sky130_fd_sc_hd__buf_2
X_12231_ _12273_/A _24012_/Q VGND VGND VPWR VPWR _12232_/C sky130_fd_sc_hd__or2_4
XFILLER_136_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21429_ _21247_/X _21427_/X _23858_/Q _21424_/X VGND VGND VPWR VPWR _23858_/D sky130_fd_sc_hd__o22a_4
X_24217_ _24182_/CLK _24217_/D HRESETn VGND VGND VPWR VPWR _24217_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22443__A2 _22438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12162_ _11786_/X _12162_/B _12161_/X VGND VGND VPWR VPWR _12178_/B sky130_fd_sc_hd__and3_4
XFILLER_2_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24148_ _24271_/CLK _20050_/Y HRESETn VGND VGND VPWR VPWR _16958_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11984__A _11973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24079_ _23983_/CLK _24079_/D VGND VGND VPWR VPWR _16283_/B sky130_fd_sc_hd__dfxtp_4
X_16970_ _16970_/A VGND VGND VPWR VPWR _17748_/A sky130_fd_sc_hd__inv_2
X_12093_ _12001_/X VGND VGND VPWR VPWR _12093_/X sky130_fd_sc_hd__buf_2
XFILLER_7_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15921_ _13782_/X _13949_/Y _13784_/A VGND VGND VPWR VPWR _15921_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_162_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21954__B2 _21950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18640_ _18545_/A _17618_/Y VGND VGND VPWR VPWR _18640_/X sky130_fd_sc_hd__and2_4
XANTENNA__23535__CLK _23246_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15852_ _13542_/A _15850_/X _15851_/X VGND VGND VPWR VPWR _15852_/X sky130_fd_sc_hd__and3_4
XFILLER_49_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14803_ _14669_/A VGND VGND VPWR VPWR _14823_/A sky130_fd_sc_hd__buf_2
X_18571_ _17730_/X _18570_/X _17730_/X _18570_/X VGND VGND VPWR VPWR _18571_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15903__B _15833_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15783_ _12979_/A _15783_/B _15783_/C VGND VGND VPWR VPWR _15783_/X sky130_fd_sc_hd__and3_4
X_12995_ _12875_/A _12995_/B VGND VGND VPWR VPWR _12995_/X sky130_fd_sc_hd__or2_4
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17522_ _13270_/X _17522_/B VGND VGND VPWR VPWR _17522_/X sky130_fd_sc_hd__or2_4
XANTENNA__13704__A _13704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14734_ _11967_/A _14733_/X VGND VGND VPWR VPWR _14734_/X sky130_fd_sc_hd__and2_4
X_11946_ _16742_/A _11774_/B VGND VGND VPWR VPWR _11946_/X sky130_fd_sc_hd__or2_4
XANTENNA__21182__A2 _21155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17453_ _12914_/X VGND VGND VPWR VPWR _17453_/Y sky130_fd_sc_hd__inv_2
X_14665_ _14665_/A VGND VGND VPWR VPWR _14675_/A sky130_fd_sc_hd__buf_2
X_11877_ _11877_/A VGND VGND VPWR VPWR _11878_/A sky130_fd_sc_hd__buf_2
XFILLER_33_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16404_ _12561_/A VGND VGND VPWR VPWR _16413_/A sky130_fd_sc_hd__buf_2
XANTENNA__22736__B HREADY VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13616_ _13990_/A VGND VGND VPWR VPWR _13617_/A sky130_fd_sc_hd__buf_2
X_17384_ _15784_/X _18406_/B VGND VGND VPWR VPWR _17384_/X sky130_fd_sc_hd__and2_4
XANTENNA__17138__A1 _14701_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14596_ _15398_/A _14592_/X _14596_/C VGND VGND VPWR VPWR _14596_/X sky130_fd_sc_hd__or3_4
XANTENNA__22131__B2 _22130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19123_ _20990_/A _18963_/X _11515_/Y _18968_/X VGND VGND VPWR VPWR _19123_/Y sky130_fd_sc_hd__a22oi_4
X_16335_ _16342_/A _16274_/B VGND VGND VPWR VPWR _16335_/X sky130_fd_sc_hd__or2_4
XFILLER_41_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13547_ _13547_/A _13544_/X _13547_/C VGND VGND VPWR VPWR _13548_/C sky130_fd_sc_hd__and3_4
XANTENNA__22682__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20256__B _16918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19054_ _19054_/A VGND VGND VPWR VPWR _19054_/Y sky130_fd_sc_hd__inv_2
X_16266_ _11890_/X _16266_/B VGND VGND VPWR VPWR _16266_/X sky130_fd_sc_hd__or2_4
X_13478_ _12869_/A _13476_/X _13477_/X VGND VGND VPWR VPWR _13478_/X sky130_fd_sc_hd__and3_4
XFILLER_127_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14254__B _23231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18005_ _17583_/B _18004_/X _17588_/Y VGND VGND VPWR VPWR _18005_/Y sky130_fd_sc_hd__o21ai_4
X_15217_ _14663_/A _15217_/B _15216_/X VGND VGND VPWR VPWR _15218_/C sky130_fd_sc_hd__and3_4
XANTENNA__22434__A2 _22426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12429_ _12862_/A VGND VGND VPWR VPWR _12440_/A sky130_fd_sc_hd__buf_2
X_16197_ _16185_/A _16193_/X _16196_/X VGND VGND VPWR VPWR _16197_/X sky130_fd_sc_hd__and3_4
XFILLER_127_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12055__A _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21642__B1 _23743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15148_ _14171_/A _15146_/X _15147_/X VGND VGND VPWR VPWR _15152_/B sky130_fd_sc_hd__and3_4
XANTENNA__24310__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24498__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11894__A _13792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15366__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19956_ _19956_/A VGND VGND VPWR VPWR _19956_/X sky130_fd_sc_hd__buf_2
X_15079_ _15103_/A _15003_/B VGND VGND VPWR VPWR _15081_/B sky130_fd_sc_hd__or2_4
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14270__A _14270_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18907_ _18900_/A VGND VGND VPWR VPWR _18907_/X sky130_fd_sc_hd__buf_2
XANTENNA__15085__B _23893_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19887_ _19553_/X _19886_/X _22798_/A _19553_/X VGND VGND VPWR VPWR _19887_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18838_ _18837_/X VGND VGND VPWR VPWR _18838_/X sky130_fd_sc_hd__buf_2
XFILLER_67_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15813__B _15868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18769_ _17015_/X _17089_/A _17085_/A _18768_/Y VGND VGND VPWR VPWR _18769_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20800_ _22461_/A VGND VGND VPWR VPWR _20801_/A sky130_fd_sc_hd__buf_2
XANTENNA__13614__A _14297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21780_ _21558_/X _21777_/X _23655_/Q _21774_/X VGND VGND VPWR VPWR _23655_/D sky130_fd_sc_hd__o22a_4
XFILLER_24_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22370__B2 _22366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21831__A _20486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20731_ _20495_/A VGND VGND VPWR VPWR _20731_/X sky130_fd_sc_hd__buf_2
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20381__B1 _20235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23450_ _24057_/CLK _22160_/X VGND VGND VPWR VPWR _23450_/Q sky130_fd_sc_hd__dfxtp_4
X_20662_ _20261_/X VGND VGND VPWR VPWR _20662_/X sky130_fd_sc_hd__buf_2
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22401_ _22165_/X _22397_/X _15136_/B _22366_/A VGND VGND VPWR VPWR _22401_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23381_ _23392_/CLK _23381_/D VGND VGND VPWR VPWR _23381_/Q sky130_fd_sc_hd__dfxtp_4
X_20593_ _20535_/X _20592_/X VGND VGND VPWR VPWR _20593_/X sky130_fd_sc_hd__or2_4
XANTENNA__14445__A _12445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22332_ _12803_/B VGND VGND VPWR VPWR _22332_/X sky130_fd_sc_hd__buf_2
X_22263_ _22153_/X _22258_/X _14391_/B _22262_/X VGND VGND VPWR VPWR _22263_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16660__A _16682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24002_ _23587_/CLK _24002_/D VGND VGND VPWR VPWR _15478_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_151_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21214_ _20693_/X _21212_/X _15820_/B _21209_/X VGND VGND VPWR VPWR _21214_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22194_ _22194_/A VGND VGND VPWR VPWR _22194_/X sky130_fd_sc_hd__buf_2
XFILLER_132_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21145_ _21137_/X VGND VGND VPWR VPWR _21145_/X sky130_fd_sc_hd__buf_2
XANTENNA__15276__A _14114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22189__A1 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22189__B2 _22184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21076_ _20959_/X _21073_/X _24056_/Q _21070_/X VGND VGND VPWR VPWR _21076_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18587__A _18545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21936__B2 _21899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20027_ _20027_/A VGND VGND VPWR VPWR _20027_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17491__A _13485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18801__A1 _12419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11800_ _11832_/A _21705_/A VGND VGND VPWR VPWR _11802_/B sky130_fd_sc_hd__or2_4
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _13067_/A VGND VGND VPWR VPWR _12780_/X sky130_fd_sc_hd__buf_2
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21164__A2 _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21978_ _21957_/A VGND VGND VPWR VPWR _21978_/X sky130_fd_sc_hd__buf_2
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21741__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23717_ _23241_/CLK _21683_/X VGND VGND VPWR VPWR _23717_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11731_ _12156_/A _23540_/Q VGND VGND VPWR VPWR _11731_/X sky130_fd_sc_hd__or2_4
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20929_ _20781_/X _20928_/X _19134_/A _20791_/X VGND VGND VPWR VPWR _20929_/X sky130_fd_sc_hd__o22a_4
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14450_/A _14449_/X VGND VGND VPWR VPWR _14450_/X sky130_fd_sc_hd__and2_4
XFILLER_42_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _14369_/A VGND VGND VPWR VPWR _12955_/A sky130_fd_sc_hd__buf_2
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23648_ _24096_/CLK _23648_/D VGND VGND VPWR VPWR _23648_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13374_/A _23110_/Q VGND VGND VPWR VPWR _13403_/B sky130_fd_sc_hd__or2_4
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18868__A1 _17169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14381_ _13937_/A VGND VGND VPWR VPWR _14511_/A sky130_fd_sc_hd__buf_2
X_11593_ _11593_/A VGND VGND VPWR VPWR _17038_/A sky130_fd_sc_hd__buf_2
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22664__A2 _22658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23579_ _23515_/CLK _23579_/D VGND VGND VPWR VPWR _14500_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_167_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16120_ _16145_/A _16116_/X _16120_/C VGND VGND VPWR VPWR _16120_/X sky130_fd_sc_hd__or3_4
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ _13332_/A _23110_/Q VGND VGND VPWR VPWR _13332_/X sky130_fd_sc_hd__or2_4
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22572__A _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24333__CLK _24294_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16051_ _11693_/X _16051_/B _16050_/X VGND VGND VPWR VPWR _16052_/C sky130_fd_sc_hd__or3_4
XFILLER_157_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13263_ _13262_/X VGND VGND VPWR VPWR _13270_/A sky130_fd_sc_hd__inv_2
XFILLER_136_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15002_ _13965_/A _15000_/X _15002_/C VGND VGND VPWR VPWR _15002_/X sky130_fd_sc_hd__and3_4
XFILLER_142_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12214_ _15439_/A VGND VGND VPWR VPWR _12228_/A sky130_fd_sc_hd__buf_2
XANTENNA__21188__A _21195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13194_ _11675_/A VGND VGND VPWR VPWR _13229_/A sky130_fd_sc_hd__buf_2
XFILLER_29_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12145_ _12169_/A _12145_/B _12144_/X VGND VGND VPWR VPWR _12146_/C sky130_fd_sc_hd__or3_4
X_19810_ _19888_/B _19808_/Y _19809_/Y VGND VGND VPWR VPWR _19810_/X sky130_fd_sc_hd__a21o_4
XANTENNA__15186__A _14773_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12603__A _12950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14090__A _12218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24483__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21916__A _21909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16953_ _17676_/A VGND VGND VPWR VPWR _17703_/A sky130_fd_sc_hd__inv_2
XFILLER_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19741_ _19682_/A _19741_/B VGND VGND VPWR VPWR _19777_/A sky130_fd_sc_hd__or2_4
X_12076_ _12028_/X _12043_/X _12054_/X _12067_/X _12075_/X VGND VGND VPWR VPWR _12076_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13418__B _13417_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15904_ _13496_/A _15834_/B VGND VGND VPWR VPWR _15904_/X sky130_fd_sc_hd__or2_4
X_19672_ _19519_/X HRDATA[9] _20422_/B _19518_/X VGND VGND VPWR VPWR _19672_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__15914__A _15849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16884_ _16884_/A _16880_/X _16881_/Y _16884_/D VGND VGND VPWR VPWR _16884_/X sky130_fd_sc_hd__and4_4
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18623_ _20196_/A VGND VGND VPWR VPWR _18623_/Y sky130_fd_sc_hd__inv_2
X_15835_ _12873_/A _15833_/X _15834_/X VGND VGND VPWR VPWR _15835_/X sky130_fd_sc_hd__and3_4
XANTENNA__13434__A _13475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18554_ _18553_/A _16977_/X _18534_/Y VGND VGND VPWR VPWR _18554_/Y sky130_fd_sc_hd__a21oi_4
X_15766_ _13092_/A _15758_/X _15765_/X VGND VGND VPWR VPWR _15782_/B sky130_fd_sc_hd__and3_4
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12978_ _12978_/A _12978_/B _12978_/C VGND VGND VPWR VPWR _12979_/C sky130_fd_sc_hd__or3_4
XFILLER_18_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24382__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17505_ _17503_/B VGND VGND VPWR VPWR _18334_/B sky130_fd_sc_hd__inv_2
X_14717_ _13823_/A _14717_/B VGND VGND VPWR VPWR _14718_/C sky130_fd_sc_hd__or2_4
X_11929_ _11929_/A VGND VGND VPWR VPWR _11930_/A sky130_fd_sc_hd__buf_2
X_18485_ _18485_/A _18466_/A VGND VGND VPWR VPWR _18487_/C sky130_fd_sc_hd__nor2_4
X_15697_ _12735_/A _15762_/B VGND VGND VPWR VPWR _15697_/X sky130_fd_sc_hd__or2_4
XFILLER_60_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16745__A _11990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17436_ _17436_/A _17436_/B _17436_/C _17435_/Y VGND VGND VPWR VPWR _17437_/B sky130_fd_sc_hd__or4_4
XANTENNA__21370__B _21370_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14648_ _13866_/A VGND VGND VPWR VPWR _14657_/A sky130_fd_sc_hd__buf_2
XFILLER_159_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20267__A _18889_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22104__B2 _22094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11889__A _13455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _16918_/A _17378_/A _17358_/Y VGND VGND VPWR VPWR _17367_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18859__A1 _12980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14579_ _13593_/A _14577_/X _14578_/X VGND VGND VPWR VPWR _14579_/X sky130_fd_sc_hd__and3_4
XANTENNA__18960__A _11544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19106_ _19021_/A VGND VGND VPWR VPWR _19106_/X sky130_fd_sc_hd__buf_2
X_16318_ _16318_/A _16253_/B VGND VGND VPWR VPWR _16319_/C sky130_fd_sc_hd__or2_4
X_17298_ _22687_/A _17039_/X _11855_/A _17297_/X VGND VGND VPWR VPWR _17298_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19037_ _19016_/X _19035_/Y _19036_/Y _19021_/X VGND VGND VPWR VPWR _19037_/X sky130_fd_sc_hd__o22a_4
X_16249_ _16155_/A _16247_/X _16248_/X VGND VGND VPWR VPWR _16255_/B sky130_fd_sc_hd__and3_4
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21091__B2 _21087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13609__A _15423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19791__A HRDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12513__A _12513_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19939_ _22745_/A VGND VGND VPWR VPWR _19939_/X sky130_fd_sc_hd__buf_2
XANTENNA__21918__B2 _21913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22950_ _18590_/X _22938_/B VGND VGND VPWR VPWR _22951_/C sky130_fd_sc_hd__or2_4
XANTENNA__21394__A2 _21391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18795__B1 _24464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21901_ _21824_/X _21895_/X _16271_/B _21899_/X VGND VGND VPWR VPWR _23599_/D sky130_fd_sc_hd__o22a_4
XFILLER_83_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22881_ _22876_/X _22823_/X _13692_/Y _22877_/X VGND VGND VPWR VPWR _22881_/X sky130_fd_sc_hd__o22a_4
XFILLER_83_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13344__A _12833_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_120_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR _23656_/CLK sky130_fd_sc_hd__clkbuf_1
X_21832_ _21831_/X _21827_/X _23628_/Q _21822_/X VGND VGND VPWR VPWR _23628_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24206__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21146__A2 _21141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21561__A _21549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21763_ _21770_/A VGND VGND VPWR VPWR _21763_/X sky130_fd_sc_hd__buf_2
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23502_ _24078_/CLK _23502_/D VGND VGND VPWR VPWR _16076_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_19_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20714_ _20714_/A VGND VGND VPWR VPWR _20714_/X sky130_fd_sc_hd__buf_2
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21694_ _21582_/X _21691_/X _23709_/Q _21688_/X VGND VGND VPWR VPWR _23709_/D sky130_fd_sc_hd__o22a_4
X_24482_ _24134_/CLK _24482_/D HRESETn VGND VGND VPWR VPWR _24482_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13998__B _24096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24356__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23433_ _23561_/CLK _22195_/X VGND VGND VPWR VPWR _23433_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19966__A _17793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20645_ _18835_/X VGND VGND VPWR VPWR _20645_/X sky130_fd_sc_hd__buf_2
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22646__A2 _22644_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23364_ _23588_/CLK _22302_/X VGND VGND VPWR VPWR _15660_/B sky130_fd_sc_hd__dfxtp_4
X_20576_ _20533_/X _20575_/X _24104_/Q _20510_/X VGND VGND VPWR VPWR _24104_/D sky130_fd_sc_hd__o22a_4
XFILLER_30_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22315_ _22275_/A VGND VGND VPWR VPWR _22315_/X sky130_fd_sc_hd__buf_2
X_23295_ _23294_/CLK _23295_/D VGND VGND VPWR VPWR _23295_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16390__A _16007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23380__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20409__A1 _18062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22246_ _22125_/X _22244_/X _13028_/B _22241_/X VGND VGND VPWR VPWR _23400_/D sky130_fd_sc_hd__o22a_4
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20300__A2_N _20225_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13519__A _13562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22177_ _22184_/A VGND VGND VPWR VPWR _22177_/X sky130_fd_sc_hd__buf_2
X_21128_ _20959_/X _21125_/X _24024_/Q _21122_/X VGND VGND VPWR VPWR _24024_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20640__A _16899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21059_ _21045_/A VGND VGND VPWR VPWR _21059_/X sky130_fd_sc_hd__buf_2
X_13950_ _13863_/X _13947_/X _13949_/Y VGND VGND VPWR VPWR _13950_/X sky130_fd_sc_hd__a21o_4
XFILLER_59_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18110__A _17906_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21385__A2 _21384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12901_ _12511_/A _23241_/Q VGND VGND VPWR VPWR _12903_/B sky130_fd_sc_hd__or2_4
XANTENNA__22582__B2 _22576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13881_ _15330_/A VGND VGND VPWR VPWR _13882_/A sky130_fd_sc_hd__buf_2
XFILLER_100_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13254__A _12338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15620_ _15620_/A _23969_/Q VGND VGND VPWR VPWR _15621_/C sky130_fd_sc_hd__or2_4
X_12832_ _13556_/A _12826_/X _12831_/X VGND VGND VPWR VPWR _12832_/X sky130_fd_sc_hd__or3_4
XFILLER_43_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15551_ _14480_/A _15528_/X _15535_/X _15542_/X _15550_/X VGND VGND VPWR VPWR _15551_/X
+ sky130_fd_sc_hd__a32o_4
X_12763_ _12775_/A _12763_/B VGND VGND VPWR VPWR _12764_/C sky130_fd_sc_hd__or2_4
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20345__B1 _24466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17210__B1 _12093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14502_ _14510_/A _14502_/B VGND VGND VPWR VPWR _14502_/X sky130_fd_sc_hd__or2_4
X_11714_ _11714_/A VGND VGND VPWR VPWR _11715_/A sky130_fd_sc_hd__buf_2
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18270_ _17490_/A _18269_/X VGND VGND VPWR VPWR _18270_/X sky130_fd_sc_hd__or2_4
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _13058_/A _15482_/B _15481_/X VGND VGND VPWR VPWR _15482_/X sky130_fd_sc_hd__and3_4
X_12694_ _12687_/A _23786_/Q VGND VGND VPWR VPWR _12695_/C sky130_fd_sc_hd__or2_4
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_25_0_HCLK clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _11610_/X _17181_/Y _17847_/A _17220_/X VGND VGND VPWR VPWR _17222_/A sky130_fd_sc_hd__o22a_4
X_14433_ _12455_/A _14495_/B VGND VGND VPWR VPWR _14433_/X sky130_fd_sc_hd__or2_4
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11644_/X _17060_/A VGND VGND VPWR VPWR _11645_/X sky130_fd_sc_hd__and2_4
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18780__A _18779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14085__A _14086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17152_ _13781_/X VGND VGND VPWR VPWR _17153_/A sky130_fd_sc_hd__buf_2
X_14364_ _14543_/A _14362_/X _14363_/X VGND VGND VPWR VPWR _14364_/X sky130_fd_sc_hd__and3_4
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11576_ _24462_/Q IRQ[25] _11575_/X VGND VGND VPWR VPWR _11576_/X sky130_fd_sc_hd__a21o_4
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16103_ _16144_/A _16103_/B _16103_/C VGND VGND VPWR VPWR _16104_/C sky130_fd_sc_hd__and3_4
X_13315_ _12904_/A _13311_/X _13314_/X VGND VGND VPWR VPWR _13315_/X sky130_fd_sc_hd__or3_4
XFILLER_155_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17083_ _17188_/A _17083_/B VGND VGND VPWR VPWR _18517_/A sky130_fd_sc_hd__or2_4
X_14295_ _14295_/A _14359_/B VGND VGND VPWR VPWR _14297_/B sky130_fd_sc_hd__or2_4
XFILLER_170_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16034_ _16046_/A _23310_/Q VGND VGND VPWR VPWR _16034_/X sky130_fd_sc_hd__or2_4
X_13246_ _13253_/A _23815_/Q VGND VGND VPWR VPWR _13246_/X sky130_fd_sc_hd__or2_4
XFILLER_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13429__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13177_ _13333_/A _24103_/Q VGND VGND VPWR VPWR _13177_/X sky130_fd_sc_hd__or2_4
XANTENNA__12333__A _11701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13148__B _13148_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20820__B2 _20746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12128_ _12164_/A _12128_/B VGND VGND VPWR VPWR _12128_/X sky130_fd_sc_hd__or2_4
X_17985_ _17849_/A VGND VGND VPWR VPWR _17985_/X sky130_fd_sc_hd__buf_2
XFILLER_111_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19724_ _19724_/A VGND VGND VPWR VPWR _19725_/A sky130_fd_sc_hd__inv_2
XFILLER_38_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16936_ _16936_/A VGND VGND VPWR VPWR _16936_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12059_ _11990_/A VGND VGND VPWR VPWR _12059_/X sky130_fd_sc_hd__buf_2
XANTENNA__15644__A _13884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24229__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18020__A _18019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22573__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19655_ _19600_/X _19655_/B _19651_/X _19655_/D VGND VGND VPWR VPWR _19655_/X sky130_fd_sc_hd__or4_4
X_16867_ _15048_/X _16866_/X _15120_/Y _15385_/X VGND VGND VPWR VPWR _16867_/X sky130_fd_sc_hd__a211o_4
XFILLER_77_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13164__A _13164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15818_ _13339_/A _15795_/X _15802_/X _15809_/X _15817_/X VGND VGND VPWR VPWR _15818_/X
+ sky130_fd_sc_hd__a32o_4
X_18606_ _17311_/Y _18604_/X VGND VGND VPWR VPWR _18606_/X sky130_fd_sc_hd__or2_4
X_19586_ _19445_/A _19585_/X HRDATA[7] _19461_/A VGND VGND VPWR VPWR _19643_/A sky130_fd_sc_hd__o22a_4
XFILLER_129_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21128__A2 _21125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16798_ _16791_/A _16798_/B VGND VGND VPWR VPWR _16798_/X sky130_fd_sc_hd__or2_4
XFILLER_19_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23253__CLK _23904_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21381__A _21381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18537_ _18536_/X VGND VGND VPWR VPWR _18537_/Y sky130_fd_sc_hd__inv_2
X_15749_ _11689_/X _15745_/X _15748_/X VGND VGND VPWR VPWR _15750_/C sky130_fd_sc_hd__or3_4
XFILLER_18_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17201__B1 _12093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18468_ _18420_/X VGND VGND VPWR VPWR _18468_/Y sky130_fd_sc_hd__inv_2
X_17419_ _14086_/A _17020_/X _17020_/X _17418_/X VGND VGND VPWR VPWR _17421_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18399_ _11642_/A VGND VGND VPWR VPWR _18399_/X sky130_fd_sc_hd__buf_2
X_20430_ _20277_/X _20428_/X _24398_/Q _20429_/X VGND VGND VPWR VPWR _20430_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20725__A _20257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15819__A _12847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20361_ _21532_/A VGND VGND VPWR VPWR _20361_/X sky130_fd_sc_hd__buf_2
XANTENNA__14723__A _12190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22100_ _22097_/X _22099_/X _12136_/B _22094_/X VGND VGND VPWR VPWR _23475_/D sky130_fd_sc_hd__o22a_4
XFILLER_173_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23080_ _23080_/A _23078_/X _23080_/C VGND VGND VPWR VPWR _23080_/X sky130_fd_sc_hd__and3_4
X_20292_ _20292_/A _20266_/X _20292_/C VGND VGND VPWR VPWR _20292_/X sky130_fd_sc_hd__and3_4
XFILLER_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_45_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR _23533_/CLK sky130_fd_sc_hd__clkbuf_1
X_22031_ _21991_/A VGND VGND VPWR VPWR _22031_/X sky130_fd_sc_hd__buf_2
XANTENNA__13339__A _13339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21064__B2 _21063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12243__A _12258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15818__A1 _13339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15554__A _12236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23982_ _24078_/CLK _21199_/X VGND VGND VPWR VPWR _23982_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21367__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22564__B2 _22562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22933_ _22945_/A _22933_/B _22933_/C VGND VGND VPWR VPWR HADDR[5] sky130_fd_sc_hd__and3_4
XFILLER_84_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22864_ _17453_/Y _22847_/X _22853_/X _22863_/X VGND VGND VPWR VPWR _22865_/A sky130_fd_sc_hd__a211o_4
XFILLER_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22387__A _22358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22316__B2 _22312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21815_ _21839_/A VGND VGND VPWR VPWR _21815_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22795_ _22794_/Y _22791_/X VGND VGND VPWR VPWR _22795_/Y sky130_fd_sc_hd__nor2_4
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13802__A _13617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21746_ _21584_/X _21741_/X _14366_/B _21745_/X VGND VGND VPWR VPWR _23676_/D sky130_fd_sc_hd__o22a_4
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24465_ _23379_/CLK _18794_/X HRESETn VGND VGND VPWR VPWR _24465_/Q sky130_fd_sc_hd__dfrtp_4
X_21677_ _21677_/A VGND VGND VPWR VPWR _21677_/X sky130_fd_sc_hd__buf_2
XANTENNA__12418__A _13566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23416_ _23416_/CLK _23416_/D VGND VGND VPWR VPWR _23416_/Q sky130_fd_sc_hd__dfxtp_4
X_20628_ _20234_/X _20616_/X _20537_/X _20627_/Y VGND VGND VPWR VPWR _20628_/X sky130_fd_sc_hd__a211o_4
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20635__A _20533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24396_ _24398_/CLK _24396_/D HRESETn VGND VGND VPWR VPWR _24396_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20559_ _21268_/A VGND VGND VPWR VPWR _20559_/X sky130_fd_sc_hd__buf_2
X_23347_ _23347_/CLK _23347_/D VGND VGND VPWR VPWR _12142_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20354__B _20353_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13100_ _13100_/A _13100_/B _13099_/X VGND VGND VPWR VPWR _13108_/B sky130_fd_sc_hd__or3_4
XANTENNA__24183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14080_ _11698_/A _14080_/B _14080_/C VGND VGND VPWR VPWR _14080_/X sky130_fd_sc_hd__and3_4
X_23278_ _23662_/CLK _23278_/D VGND VGND VPWR VPWR _23278_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21055__B2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13249__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13031_ _12911_/A _13031_/B _13030_/X VGND VGND VPWR VPWR _13031_/X sky130_fd_sc_hd__or3_4
XANTENNA__23126__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22229_ _22258_/A VGND VGND VPWR VPWR _22244_/A sky130_fd_sc_hd__buf_2
XFILLER_156_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20802__B2 _20746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_2_0_HCLK clkbuf_5_1_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11992__A _11939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17770_ _17770_/A _17703_/X VGND VGND VPWR VPWR _17770_/Y sky130_fd_sc_hd__nand2_4
X_14982_ _11665_/X _14950_/X _14981_/X VGND VGND VPWR VPWR _14983_/A sky130_fd_sc_hd__and3_4
XANTENNA__21358__A2 _21355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16721_ _16691_/A _23985_/Q VGND VGND VPWR VPWR _16722_/C sky130_fd_sc_hd__or2_4
X_13933_ _13706_/A _13933_/B VGND VGND VPWR VPWR _13933_/X sky130_fd_sc_hd__or2_4
XFILLER_75_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19440_ _19512_/A VGND VGND VPWR VPWR _19719_/A sky130_fd_sc_hd__buf_2
X_16652_ _16786_/A _16642_/X _16652_/C VGND VGND VPWR VPWR _16652_/X sky130_fd_sc_hd__and3_4
XANTENNA__13048__A1 _11856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13864_ _11680_/A VGND VGND VPWR VPWR _13894_/A sky130_fd_sc_hd__buf_2
XFILLER_90_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22307__B2 _22305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15603_ _12337_/A _15603_/B _15602_/X VGND VGND VPWR VPWR _15603_/X sky130_fd_sc_hd__and3_4
X_12815_ _13563_/A _12811_/X _12815_/C VGND VGND VPWR VPWR _12815_/X sky130_fd_sc_hd__or3_4
X_19371_ _19369_/X _18626_/X _19369_/X _24251_/Q VGND VGND VPWR VPWR _24251_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16583_ _16588_/A _16581_/X _16583_/C VGND VGND VPWR VPWR _16584_/C sky130_fd_sc_hd__and3_4
X_13795_ _14574_/A VGND VGND VPWR VPWR _14304_/A sky130_fd_sc_hd__buf_2
XFILLER_37_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18322_ _18206_/X _18294_/X _18206_/X _18291_/X VGND VGND VPWR VPWR _18322_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15534_ _14418_/X _15532_/X _15533_/X VGND VGND VPWR VPWR _15534_/X sky130_fd_sc_hd__and3_4
X_12746_ _13183_/A _23722_/Q VGND VGND VPWR VPWR _12746_/X sky130_fd_sc_hd__or2_4
XFILLER_31_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14527__B _14463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18253_ _18253_/A VGND VGND VPWR VPWR _18253_/Y sky130_fd_sc_hd__inv_2
X_15465_ _15477_/A _15465_/B VGND VGND VPWR VPWR _15465_/X sky130_fd_sc_hd__or2_4
X_12677_ _12979_/A _12677_/B _12677_/C VGND VGND VPWR VPWR _12677_/X sky130_fd_sc_hd__and3_4
XFILLER_124_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12328__A _12580_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _17173_/Y _17192_/X _15913_/Y _17193_/X VGND VGND VPWR VPWR _17204_/X sky130_fd_sc_hd__o22a_4
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14416_ _14334_/X _14413_/Y VGND VGND VPWR VPWR _14417_/B sky130_fd_sc_hd__and2_4
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18184_ _17769_/X _18183_/X _17769_/X _18183_/X VGND VGND VPWR VPWR _18184_/X sky130_fd_sc_hd__a2bb2o_4
X_11628_ _11628_/A VGND VGND VPWR VPWR _11629_/A sky130_fd_sc_hd__buf_2
X_15396_ _15400_/A _23746_/Q VGND VGND VPWR VPWR _15397_/C sky130_fd_sc_hd__or2_4
XFILLER_129_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17135_ _17130_/X _17134_/X VGND VGND VPWR VPWR _17135_/X sky130_fd_sc_hd__and2_4
XANTENNA__21294__B2 _21288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15639__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14347_ _14513_/A _14340_/X _14346_/X VGND VGND VPWR VPWR _14347_/X sky130_fd_sc_hd__or3_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11559_ _11550_/X _11551_/X _11553_/X _11558_/X VGND VGND VPWR VPWR _11559_/X sky130_fd_sc_hd__or4_4
XFILLER_143_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20264__B _18889_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17066_ _17060_/X _17096_/A _11643_/Y _17017_/B VGND VGND VPWR VPWR _17070_/B sky130_fd_sc_hd__a211o_4
XFILLER_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14278_ _14278_/A _14349_/B VGND VGND VPWR VPWR _14278_/X sky130_fd_sc_hd__or2_4
XANTENNA__22760__A SYSTICKCLKDIV[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16017_ _16031_/A _23278_/Q VGND VGND VPWR VPWR _16017_/X sky130_fd_sc_hd__or2_4
XANTENNA__13159__A _11970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21046__B2 _21042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13229_ _13229_/A _13229_/B _13229_/C VGND VGND VPWR VPWR _13229_/X sky130_fd_sc_hd__or3_4
XFILLER_170_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21376__A _21405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12998__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15374__A _12580_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17968_ _18222_/A _17968_/B VGND VGND VPWR VPWR _17972_/B sky130_fd_sc_hd__and2_4
XANTENNA__21349__A2 _21348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22546__B2 _22541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19707_ _19683_/A VGND VGND VPWR VPWR _19742_/A sky130_fd_sc_hd__buf_2
X_16919_ _16918_/X _17060_/B _16911_/X VGND VGND VPWR VPWR _16919_/X sky130_fd_sc_hd__o21a_4
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17899_ _11642_/A VGND VGND VPWR VPWR _17900_/A sky130_fd_sc_hd__buf_2
XFILLER_81_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19638_ _19465_/A VGND VGND VPWR VPWR _19638_/X sky130_fd_sc_hd__buf_2
XFILLER_81_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22000__A _22000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19569_ _19556_/X _19559_/Y _19565_/X _19467_/X _19568_/Y VGND VGND VPWR VPWR _19569_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14718__A _12469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21600_ _21024_/A VGND VGND VPWR VPWR _21600_/X sky130_fd_sc_hd__buf_2
XANTENNA__13622__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22580_ _22473_/X _22579_/X _14560_/B _22576_/X VGND VGND VPWR VPWR _22580_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22935__A _23078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21531_ _21528_/X _21530_/X _23795_/Q _21525_/X VGND VGND VPWR VPWR _21531_/X sky130_fd_sc_hd__o22a_4
XFILLER_166_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24250_ _24248_/CLK _24250_/D HRESETn VGND VGND VPWR VPWR _24250_/Q sky130_fd_sc_hd__dfrtp_4
X_21462_ _21455_/A VGND VGND VPWR VPWR _21462_/X sky130_fd_sc_hd__buf_2
X_23201_ _23203_/CLK _23201_/D VGND VGND VPWR VPWR _23201_/Q sky130_fd_sc_hd__dfxtp_4
X_20413_ _20334_/A _20412_/X VGND VGND VPWR VPWR _20413_/X sky130_fd_sc_hd__or2_4
XANTENNA__15549__A _12288_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21393_ _21271_/X _21391_/X _23880_/Q _21388_/X VGND VGND VPWR VPWR _23880_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24181_ _24182_/CLK _19911_/Y HRESETn VGND VGND VPWR VPWR _20237_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14453__A _12455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23132_ _24096_/CLK _22677_/X VGND VGND VPWR VPWR _14387_/B sky130_fd_sc_hd__dfxtp_4
X_20344_ _20344_/A VGND VGND VPWR VPWR _20344_/X sky130_fd_sc_hd__buf_2
XFILLER_161_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13069__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23063_ _23063_/A VGND VGND VPWR VPWR HADDR[27] sky130_fd_sc_hd__inv_2
X_20275_ _20495_/A VGND VGND VPWR VPWR _20275_/X sky130_fd_sc_hd__buf_2
XANTENNA__21588__A2 _21578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22014_ _22007_/A VGND VGND VPWR VPWR _22014_/X sky130_fd_sc_hd__buf_2
XFILLER_88_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15284__A _15257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12701__A _13277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23965_ _23323_/CLK _23965_/D VGND VGND VPWR VPWR _23965_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12420__B _12419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22829__B _17319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22916_ _22908_/X _18718_/X _22909_/X _22915_/X VGND VGND VPWR VPWR _22916_/X sky130_fd_sc_hd__a211o_4
XFILLER_95_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23896_ _23098_/CLK _21365_/X VGND VGND VPWR VPWR _23896_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_140_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22847_ _22846_/X VGND VGND VPWR VPWR _22847_/X sky130_fd_sc_hd__buf_2
X_12600_ _12600_/A VGND VGND VPWR VPWR _12927_/A sky130_fd_sc_hd__buf_2
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17004__A _18576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19408__A2_N _18254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A VGND VGND VPWR VPWR _13580_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22778_ _22753_/Y _22778_/B VGND VGND VPWR VPWR _22780_/A sky130_fd_sc_hd__nand2_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21512__A2 _21506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12531_ _12531_/A VGND VGND VPWR VPWR _12875_/A sky130_fd_sc_hd__buf_2
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21729_ _21556_/X _21727_/X _23688_/Q _21724_/X VGND VGND VPWR VPWR _23688_/D sky130_fd_sc_hd__o22a_4
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15250_ _11665_/X _15218_/X _15250_/C VGND VGND VPWR VPWR _15251_/A sky130_fd_sc_hd__and3_4
XFILLER_71_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12462_ _12881_/A VGND VGND VPWR VPWR _12890_/A sky130_fd_sc_hd__buf_2
XFILLER_36_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24448_ _23476_/CLK _18819_/X HRESETn VGND VGND VPWR VPWR _24448_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14201_ _14201_/A _14199_/X _14201_/C VGND VGND VPWR VPWR _14201_/X sky130_fd_sc_hd__and3_4
XFILLER_166_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11987__A _16713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15181_ _15018_/A _15181_/B _15181_/C VGND VGND VPWR VPWR _15182_/C sky130_fd_sc_hd__and3_4
X_12393_ _12363_/X _12393_/B VGND VGND VPWR VPWR _12394_/C sky130_fd_sc_hd__or2_4
XANTENNA__14363__A _12583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24379_ _24382_/CLK _24379_/D HRESETn VGND VGND VPWR VPWR _19101_/A sky130_fd_sc_hd__dfstp_4
XFILLER_153_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18141__B2 _18140_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14132_ _12425_/A _14130_/X _14132_/C VGND VGND VPWR VPWR _14132_/X sky130_fd_sc_hd__and3_4
XFILLER_67_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18940_ _15251_/A _18934_/X _19120_/A _18935_/X VGND VGND VPWR VPWR _24375_/D sky130_fd_sc_hd__o22a_4
X_14063_ _12581_/A _23424_/Q VGND VGND VPWR VPWR _14063_/X sky130_fd_sc_hd__or2_4
XFILLER_153_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21579__A2 _21578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13014_ _12492_/A _13012_/X _13013_/X VGND VGND VPWR VPWR _13014_/X sky130_fd_sc_hd__and3_4
XANTENNA__17393__B _17448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15906__B _15836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18871_ _18842_/A VGND VGND VPWR VPWR _18871_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_91_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR _23518_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17822_ _17815_/X _17818_/X _17820_/X _17821_/X VGND VGND VPWR VPWR _17822_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22528__B2 _22526_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17753_ _17005_/A _17336_/X _17005_/A _17336_/X VGND VGND VPWR VPWR _17753_/X sky130_fd_sc_hd__a2bb2o_4
X_14965_ _15362_/A _14957_/X _14964_/X VGND VGND VPWR VPWR _14965_/X sky130_fd_sc_hd__and3_4
XFILLER_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21200__B2 _21195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16704_ _16704_/A _23697_/Q VGND VGND VPWR VPWR _16706_/B sky130_fd_sc_hd__or2_4
X_13916_ _13916_/A _23613_/Q VGND VGND VPWR VPWR _13916_/X sky130_fd_sc_hd__or2_4
X_17684_ _16988_/A _17511_/X VGND VGND VPWR VPWR _17698_/A sky130_fd_sc_hd__or2_4
X_14896_ _14114_/A _14894_/X _14896_/C VGND VGND VPWR VPWR _14896_/X sky130_fd_sc_hd__and3_4
XANTENNA__21751__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16635_ _16635_/A VGND VGND VPWR VPWR _16659_/A sky130_fd_sc_hd__buf_2
X_19423_ _19421_/X _18556_/Y _19421_/X _24222_/Q VGND VGND VPWR VPWR _19423_/X sky130_fd_sc_hd__a2bb2o_4
X_13847_ _13677_/A _13847_/B _13847_/C VGND VGND VPWR VPWR _13847_/X sky130_fd_sc_hd__and3_4
XFILLER_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14538__A _14519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13442__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19354_ _19340_/A VGND VGND VPWR VPWR _19354_/X sky130_fd_sc_hd__buf_2
X_16566_ _16594_/A _16640_/B VGND VGND VPWR VPWR _16567_/C sky130_fd_sc_hd__or2_4
X_13778_ _12597_/A _13778_/B _13777_/X VGND VGND VPWR VPWR _13778_/X sky130_fd_sc_hd__or3_4
XANTENNA__22755__A SYSTICKCLKDIV[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15517_ _15517_/A _15485_/X _15516_/X VGND VGND VPWR VPWR _15517_/X sky130_fd_sc_hd__and3_4
XANTENNA__22700__B2 _22698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18305_ _18215_/X _18300_/X _18240_/X _18304_/X VGND VGND VPWR VPWR _18305_/X sky130_fd_sc_hd__o22a_4
X_12729_ _12704_/A _12727_/X _12729_/C VGND VGND VPWR VPWR _12729_/X sky130_fd_sc_hd__and3_4
X_19285_ _19244_/B VGND VGND VPWR VPWR _19285_/Y sky130_fd_sc_hd__inv_2
X_16497_ _16490_/A _16428_/B VGND VGND VPWR VPWR _16497_/X sky130_fd_sc_hd__or2_4
XANTENNA__16753__A _16635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18236_ _17490_/B _18235_/X VGND VGND VPWR VPWR _18236_/X sky130_fd_sc_hd__or2_4
X_15448_ _12251_/A _15446_/X _15448_/C VGND VGND VPWR VPWR _15448_/X sky130_fd_sc_hd__and3_4
XFILLER_90_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11897__A _14110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21267__B2 _21264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15369__A _15369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18167_ _17600_/D _18167_/B VGND VGND VPWR VPWR _18167_/X sky130_fd_sc_hd__or2_4
X_15379_ _11665_/X _15347_/X _15378_/X VGND VGND VPWR VPWR _15380_/A sky130_fd_sc_hd__and3_4
XFILLER_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14273__A _14304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17118_ _12064_/X VGND VGND VPWR VPWR _17164_/A sky130_fd_sc_hd__buf_2
XFILLER_85_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18098_ _18095_/X _17578_/X _18096_/X _17919_/X _18097_/Y VGND VGND VPWR VPWR _18098_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15088__B _23605_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22490__A _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18683__A2 _18681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23441__CLK _23409_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17049_ _17049_/A VGND VGND VPWR VPWR _17418_/A sky130_fd_sc_hd__buf_2
XANTENNA__17891__B1 _17890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22767__A1 SYSTICKCLKDIV[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20060_ _24483_/Q VGND VGND VPWR VPWR _20060_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19632__A1 _19797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20242__A2 HRDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13617__A _13617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12521__A _12506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13336__B _13405_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15832__A _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23750_ _23750_/CLK _21632_/X VGND VGND VPWR VPWR _13280_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20962_ _21007_/A _20776_/A VGND VGND VPWR VPWR _20962_/X sky130_fd_sc_hd__or2_4
XANTENNA__21742__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22701_ _22708_/A VGND VGND VPWR VPWR _22701_/X sky130_fd_sc_hd__buf_2
XPHY_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ _23908_/CLK _23681_/D VGND VGND VPWR VPWR _23681_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ _20772_/X _20892_/X _24091_/Q _20861_/X VGND VGND VPWR VPWR _24091_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14448__A _14448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22632_ _22478_/X _22629_/X _23160_/Q _22626_/X VGND VGND VPWR VPWR _23160_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22665__A _22658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22563_ _22444_/X _22558_/X _13283_/B _22562_/X VGND VGND VPWR VPWR _23206_/D sky130_fd_sc_hd__o22a_4
XFILLER_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16663__A _16646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24302_ _24302_/CLK _24302_/D HRESETn VGND VGND VPWR VPWR _24302_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15185__A1 _13951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21514_ _21304_/X _21513_/X _14684_/B _21510_/X VGND VGND VPWR VPWR _23802_/D sky130_fd_sc_hd__o22a_4
X_22494_ _22508_/A VGND VGND VPWR VPWR _22494_/X sky130_fd_sc_hd__buf_2
XFILLER_21_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21258__B2 _21252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22455__B1 _15454_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24233_ _24127_/CLK _19408_/X HRESETn VGND VGND VPWR VPWR _24233_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15279__A _14897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21445_ _21438_/A VGND VGND VPWR VPWR _21445_/X sky130_fd_sc_hd__buf_2
XFILLER_163_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24359__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24164_ _24184_/CLK _19945_/X HRESETn VGND VGND VPWR VPWR _24164_/Q sky130_fd_sc_hd__dfrtp_4
X_21376_ _21405_/A VGND VGND VPWR VPWR _21391_/A sky130_fd_sc_hd__buf_2
X_23115_ _24074_/CLK _23115_/D VGND VGND VPWR VPWR _12564_/B sky130_fd_sc_hd__dfxtp_4
X_20327_ _20264_/X VGND VGND VPWR VPWR _20761_/A sky130_fd_sc_hd__buf_2
XFILLER_163_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24095_ _23880_/CLK _20802_/X VGND VGND VPWR VPWR _24095_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_116_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_15_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23046_ _23036_/X _17667_/A _23019_/X _23045_/X VGND VGND VPWR VPWR _23047_/A sky130_fd_sc_hd__a211o_4
X_20258_ _20257_/X VGND VGND VPWR VPWR _20259_/A sky130_fd_sc_hd__buf_2
XFILLER_131_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13527__A _12773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21430__B2 _21424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20189_ _24466_/Q IRQ[29] _20188_/X VGND VGND VPWR VPWR _20190_/B sky130_fd_sc_hd__a21boi_4
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14750_ _12190_/A _14834_/B VGND VGND VPWR VPWR _14752_/B sky130_fd_sc_hd__or2_4
X_23948_ _23728_/CLK _23948_/D VGND VGND VPWR VPWR _12357_/B sky130_fd_sc_hd__dfxtp_4
X_11962_ _12103_/A _21937_/A VGND VGND VPWR VPWR _11962_/X sky130_fd_sc_hd__or2_4
XFILLER_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_1_HCLK clkbuf_1_1_0_HCLK/X VGND VGND VPWR VPWR clkbuf_2_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21733__A2 _21727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13701_ _13710_/A VGND VGND VPWR VPWR _14541_/A sky130_fd_sc_hd__buf_2
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14681_ _14660_/A _14676_/X _14681_/C VGND VGND VPWR VPWR _14682_/C sky130_fd_sc_hd__or3_4
X_23879_ _23111_/CLK _23879_/D VGND VGND VPWR VPWR _23879_/Q sky130_fd_sc_hd__dfxtp_4
X_11893_ _16711_/A _11718_/B VGND VGND VPWR VPWR _11893_/X sky130_fd_sc_hd__or2_4
XANTENNA__14358__A _11681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16420_ _16160_/A _16393_/X _16400_/X _16411_/X _16419_/X VGND VGND VPWR VPWR _16420_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13262__A _13261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13632_ _13632_/A _23998_/Q VGND VGND VPWR VPWR _13633_/C sky130_fd_sc_hd__or2_4
XFILLER_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16351_ _16342_/A _16283_/B VGND VGND VPWR VPWR _16351_/X sky130_fd_sc_hd__or2_4
XFILLER_13_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13563_ _13563_/A _13563_/B _13563_/C VGND VGND VPWR VPWR _13564_/C sky130_fd_sc_hd__or3_4
XANTENNA__21497__B2 _21496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15302_ _13593_/A _15300_/X _15302_/C VGND VGND VPWR VPWR _15302_/X sky130_fd_sc_hd__and3_4
X_12514_ _12514_/A _12514_/B VGND VGND VPWR VPWR _12515_/C sky130_fd_sc_hd__or2_4
X_19070_ _24352_/Q _11525_/X _19064_/Y VGND VGND VPWR VPWR _19070_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_157_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16282_ _16282_/A _16282_/B VGND VGND VPWR VPWR _16282_/X sky130_fd_sc_hd__or2_4
XFILLER_125_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13494_ _15903_/A _23365_/Q VGND VGND VPWR VPWR _13497_/B sky130_fd_sc_hd__or2_4
XANTENNA__20095__A _17820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18021_ _17009_/A VGND VGND VPWR VPWR _18148_/A sky130_fd_sc_hd__buf_2
X_15233_ _14663_/A _15233_/B _15232_/X VGND VGND VPWR VPWR _15233_/X sky130_fd_sc_hd__and3_4
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12445_ _12445_/A VGND VGND VPWR VPWR _13011_/A sky130_fd_sc_hd__buf_2
XANTENNA__12606__A _13052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15164_ _15269_/A _15164_/B _15163_/X VGND VGND VPWR VPWR _15168_/B sky130_fd_sc_hd__and3_4
XFILLER_165_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12376_ _15851_/A _12376_/B VGND VGND VPWR VPWR _12377_/C sky130_fd_sc_hd__or2_4
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14115_ _15007_/A VGND VGND VPWR VPWR _14165_/A sky130_fd_sc_hd__buf_2
XFILLER_114_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15917__A _15915_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19972_ _17974_/X _17055_/A _19971_/X _17919_/X _18769_/X VGND VGND VPWR VPWR _19972_/X
+ sky130_fd_sc_hd__a32o_4
X_15095_ _15095_/A _23381_/Q VGND VGND VPWR VPWR _15095_/X sky130_fd_sc_hd__or2_4
XFILLER_153_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14821__A _15112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18923_ _15784_/X _18920_/X _24388_/Q _18921_/X VGND VGND VPWR VPWR _24388_/D sky130_fd_sc_hd__o22a_4
X_14046_ _12581_/A _23552_/Q VGND VGND VPWR VPWR _14047_/C sky130_fd_sc_hd__or2_4
XFILLER_171_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13437__A _13431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18854_ _12419_/X _18849_/X _24428_/Q _18850_/X VGND VGND VPWR VPWR _18854_/X sky130_fd_sc_hd__o22a_4
XFILLER_94_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21972__A2 _21967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17805_ _17109_/X VGND VGND VPWR VPWR _17805_/X sky130_fd_sc_hd__buf_2
XFILLER_95_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15997_ _15993_/A _15995_/X _15997_/C VGND VGND VPWR VPWR _15997_/X sky130_fd_sc_hd__and3_4
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18785_ _18785_/A VGND VGND VPWR VPWR _18786_/A sky130_fd_sc_hd__buf_2
XANTENNA__16748__A _11868_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15652__A _15651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17736_ _17736_/A VGND VGND VPWR VPWR _17737_/A sky130_fd_sc_hd__inv_2
X_14948_ _14769_/A _14944_/X _14947_/X VGND VGND VPWR VPWR _14948_/X sky130_fd_sc_hd__or3_4
XFILLER_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17667_ _17667_/A _17576_/Y VGND VGND VPWR VPWR _17667_/X sky130_fd_sc_hd__or2_4
X_14879_ _14012_/A _14855_/X _14863_/X _14870_/X _14878_/X VGND VGND VPWR VPWR _14879_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14268__A _14278_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13172__A _13304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19406_ _19324_/A VGND VGND VPWR VPWR _19406_/X sky130_fd_sc_hd__buf_2
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16618_ _16656_/A _16615_/X _16617_/X VGND VGND VPWR VPWR _16618_/X sky130_fd_sc_hd__and3_4
XFILLER_78_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17598_ _17459_/Y _17469_/A _17467_/X VGND VGND VPWR VPWR _17598_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__24215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21488__B2 _21482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19337_ _19335_/X _17896_/X _19335_/X _24274_/Q VGND VGND VPWR VPWR _19337_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23807__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16549_ _16556_/A _16549_/B _16549_/C VGND VGND VPWR VPWR _16550_/C sky130_fd_sc_hd__and3_4
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13900__A _14390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19268_ _19252_/A _19252_/B _19267_/Y VGND VGND VPWR VPWR _24303_/D sky130_fd_sc_hd__o21a_4
X_18219_ _18032_/X VGND VGND VPWR VPWR _18219_/X sky130_fd_sc_hd__buf_2
XANTENNA__15099__A _14682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19199_ _19142_/X VGND VGND VPWR VPWR _19199_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12516__A _12516_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21230_ _20980_/X _21226_/X _15156_/B _21195_/A VGND VGND VPWR VPWR _23959_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21161_ _20633_/X _21155_/X _24005_/Q _21159_/X VGND VGND VPWR VPWR _24005_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15827__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20112_ _11585_/D _20119_/A _20111_/X _20124_/B VGND VGND VPWR VPWR _20112_/X sky130_fd_sc_hd__or4_4
X_21092_ _20361_/X _21090_/X _24050_/Q _21087_/X VGND VGND VPWR VPWR _24050_/D sky130_fd_sc_hd__o22a_4
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13347__A _13385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20043_ _18328_/X _20031_/X _20041_/Y _20042_/X VGND VGND VPWR VPWR _20043_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12251__A _12251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21963__A2 _21960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23802_ _24090_/CLK _23802_/D VGND VGND VPWR VPWR _14684_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21994_ _21988_/Y _21993_/X _21811_/X _21993_/X VGND VGND VPWR VPWR _21994_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21715__A2 _21713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23733_ _23904_/CLK _23733_/D VGND VGND VPWR VPWR _23733_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ _20944_/Y _20873_/X _20561_/B _20697_/X VGND VGND VPWR VPWR _20945_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13082__A _13099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ _24080_/CLK _23664_/D VGND VGND VPWR VPWR _16439_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_6_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _24411_/Q _20316_/X VGND VGND VPWR VPWR _20876_/Y sky130_fd_sc_hd__nand2_4
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22615_ _22608_/A VGND VGND VPWR VPWR _22615_/X sky130_fd_sc_hd__buf_2
XANTENNA__21479__B2 _21475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23595_ _24012_/CLK _21907_/X VGND VGND VPWR VPWR _12619_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16393__A _15934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22140__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19541__B1 HRDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13810__A _12477_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22546_ _22416_/X _22544_/X _16621_/B _22541_/X VGND VGND VPWR VPWR _22546_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22477_ _22476_/X _22474_/X _14774_/B _22469_/X VGND VGND VPWR VPWR _23257_/D sky130_fd_sc_hd__o22a_4
X_12230_ _12269_/A VGND VGND VPWR VPWR _12273_/A sky130_fd_sc_hd__buf_2
X_24216_ _24471_/CLK _19431_/X HRESETn VGND VGND VPWR VPWR _24216_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21428_ _21243_/X _21427_/X _23859_/Q _21424_/X VGND VGND VPWR VPWR _23859_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21100__B1 _24044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21651__A1 _21594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24147_ _24127_/CLK _20054_/Y HRESETn VGND VGND VPWR VPWR _24147_/Q sky130_fd_sc_hd__dfrtp_4
X_12161_ _11694_/X _12157_/X _12161_/C VGND VGND VPWR VPWR _12161_/X sky130_fd_sc_hd__or3_4
XANTENNA__21651__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21359_ _21338_/A VGND VGND VPWR VPWR _21359_/X sky130_fd_sc_hd__buf_2
XANTENNA__18113__A _18310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24078_ _24078_/CLK _24078_/D VGND VGND VPWR VPWR _24078_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12092_ _16710_/A _12092_/B _12091_/X VGND VGND VPWR VPWR _12092_/X sky130_fd_sc_hd__or3_4
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13257__A _13235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23029_ _23029_/A VGND VGND VPWR VPWR HADDR[21] sky130_fd_sc_hd__inv_2
X_15920_ _15521_/X _15656_/X VGND VGND VPWR VPWR _15920_/X sky130_fd_sc_hd__or2_4
XFILLER_7_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12161__A _11694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21954__A2 _21953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15851_ _15851_/A _15790_/B VGND VGND VPWR VPWR _15851_/X sky130_fd_sc_hd__or2_4
XANTENNA__21474__A _21489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16568__A _16568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15472__A _12587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14802_ _14674_/A _14720_/B VGND VGND VPWR VPWR _14802_/X sky130_fd_sc_hd__or2_4
X_15782_ _12676_/A _15782_/B _15781_/X VGND VGND VPWR VPWR _15783_/C sky130_fd_sc_hd__or3_4
XANTENNA__24262__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18570_ _17760_/X _17731_/X _17727_/X VGND VGND VPWR VPWR _18570_/X sky130_fd_sc_hd__o21a_4
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12994_ _11872_/A _12990_/X _12994_/C VGND VGND VPWR VPWR _12994_/X sky130_fd_sc_hd__or3_4
XFILLER_57_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17521_ _17518_/Y _17022_/X _17029_/X _17520_/X VGND VGND VPWR VPWR _17522_/B sky130_fd_sc_hd__o22a_4
X_14733_ _11931_/A _14729_/X _14732_/X VGND VGND VPWR VPWR _14733_/X sky130_fd_sc_hd__or3_4
X_11945_ _16744_/A _21080_/A VGND VGND VPWR VPWR _11947_/B sky130_fd_sc_hd__or2_4
XFILLER_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18783__A _12027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ _18418_/A _17437_/Y _17444_/Y _17451_/Y VGND VGND VPWR VPWR _17452_/X sky130_fd_sc_hd__a211o_4
XFILLER_73_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14664_ _14819_/A _14583_/B VGND VGND VPWR VPWR _14667_/B sky130_fd_sc_hd__or2_4
X_11876_ _16145_/A VGND VGND VPWR VPWR _11876_/X sky130_fd_sc_hd__buf_2
XANTENNA__20818__A _20818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16403_ _16402_/X _16403_/B VGND VGND VPWR VPWR _16403_/X sky130_fd_sc_hd__or2_4
X_13615_ _12474_/A VGND VGND VPWR VPWR _13990_/A sky130_fd_sc_hd__buf_2
XANTENNA__22667__B1 _15826_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17383_ _17383_/A VGND VGND VPWR VPWR _18406_/B sky130_fd_sc_hd__inv_2
X_14595_ _15401_/A _14595_/B _14595_/C VGND VGND VPWR VPWR _14596_/C sky130_fd_sc_hd__and3_4
XANTENNA__22131__A2 _22123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16334_ _11727_/A VGND VGND VPWR VPWR _16342_/A sky130_fd_sc_hd__buf_2
XFILLER_125_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13720__A _13720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19122_ _19109_/X _19121_/X _18959_/A _11514_/A VGND VGND VPWR VPWR _24343_/D sky130_fd_sc_hd__a2bb2o_4
X_13546_ _13546_/A _13546_/B VGND VGND VPWR VPWR _13547_/C sky130_fd_sc_hd__or2_4
XFILLER_125_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20256__C _16922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19053_ _19053_/A VGND VGND VPWR VPWR _19053_/Y sky130_fd_sc_hd__inv_2
X_16265_ _15936_/X _16263_/X _16264_/X VGND VGND VPWR VPWR _16265_/X sky130_fd_sc_hd__and3_4
XFILLER_125_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13477_ _12895_/A _13477_/B VGND VGND VPWR VPWR _13477_/X sky130_fd_sc_hd__or2_4
XANTENNA__12336__A _12336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15216_ _14615_/A _15212_/X _15216_/C VGND VGND VPWR VPWR _15216_/X sky130_fd_sc_hd__or3_4
X_18004_ _18099_/A _18097_/A _17586_/X VGND VGND VPWR VPWR _18004_/X sky130_fd_sc_hd__o21a_4
X_12428_ _12428_/A VGND VGND VPWR VPWR _12862_/A sky130_fd_sc_hd__buf_2
X_16196_ _16219_/A _16196_/B VGND VGND VPWR VPWR _16196_/X sky130_fd_sc_hd__or2_4
XANTENNA__20445__A2 _21007_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24342__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15147_ _14170_/A _15147_/B VGND VGND VPWR VPWR _15147_/X sky130_fd_sc_hd__or2_4
XANTENNA__15647__A _14348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12359_ _12339_/X _12357_/X _12358_/X VGND VGND VPWR VPWR _12359_/X sky130_fd_sc_hd__and3_4
XANTENNA__21642__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19955_ _23083_/D VGND VGND VPWR VPWR _19956_/A sky130_fd_sc_hd__buf_2
X_15078_ _15078_/A _15075_/X _15077_/X VGND VGND VPWR VPWR _15082_/B sky130_fd_sc_hd__and3_4
XFILLER_102_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18906_ _18897_/A VGND VGND VPWR VPWR _18906_/X sky130_fd_sc_hd__buf_2
X_14029_ _14075_/A _24032_/Q VGND VGND VPWR VPWR _14032_/B sky130_fd_sc_hd__or2_4
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19886_ _19467_/X _19885_/X _19516_/X _19823_/B VGND VGND VPWR VPWR _19886_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_6_61_0_HCLK clkbuf_6_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21384__A _21391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18271__B1 _18060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18837_ _18837_/A _18837_/B VGND VGND VPWR VPWR _18837_/X sky130_fd_sc_hd__or2_4
XANTENNA__16478__A _16370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15382__A _15382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24467__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18768_ _18768_/A VGND VGND VPWR VPWR _18768_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17719_ _17718_/A _17418_/X VGND VGND VPWR VPWR _17720_/B sky130_fd_sc_hd__nor2_4
XFILLER_82_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18699_ _16970_/A _18698_/X _18630_/X VGND VGND VPWR VPWR _18699_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18693__A _17801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22370__A2 _22369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20730_ _20730_/A _20730_/B VGND VGND VPWR VPWR _20730_/X sky130_fd_sc_hd__or2_4
XFILLER_91_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20661_ _20229_/X VGND VGND VPWR VPWR _20661_/X sky130_fd_sc_hd__buf_2
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14726__A _14331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18326__B2 _18325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22400_ _22163_/X _22397_/X _15264_/B _22394_/X VGND VGND VPWR VPWR _23288_/D sky130_fd_sc_hd__o22a_4
XFILLER_149_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20592_ _24263_/Q _20443_/X _20591_/X VGND VGND VPWR VPWR _20592_/X sky130_fd_sc_hd__o21a_4
X_23380_ _23476_/CLK _23380_/D VGND VGND VPWR VPWR _11745_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_137_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22943__A _22931_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22331_ _23339_/Q VGND VGND VPWR VPWR _23339_/D sky130_fd_sc_hd__buf_2
XANTENNA__12246__A _12298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22262_ _22226_/A VGND VGND VPWR VPWR _22262_/X sky130_fd_sc_hd__buf_2
XANTENNA__20463__A _22113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24135__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24001_ _23908_/CLK _24001_/D VGND VGND VPWR VPWR _24001_/Q sky130_fd_sc_hd__dfxtp_4
X_21213_ _20659_/X _21212_/X _15688_/B _21209_/X VGND VGND VPWR VPWR _23972_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15557__A _14418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21633__B2 _21631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22193_ _22120_/X _22187_/X _12731_/B _22191_/X VGND VGND VPWR VPWR _23434_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14461__A _12428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21144_ _20378_/X _21141_/X _24017_/Q _21138_/X VGND VGND VPWR VPWR _24017_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15312__A1 _14302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22189__A2 _22187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21075_ _20938_/X _21073_/X _24057_/Q _21070_/X VGND VGND VPWR VPWR _24057_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24285__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21936__A2 _21909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20026_ _20026_/A VGND VGND VPWR VPWR _20026_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13805__A _12445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24137__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11637__B1 NMI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21977_ _21867_/X _21974_/X _13819_/B _21971_/X VGND VGND VPWR VPWR _23549_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22837__B _17284_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23716_ _23523_/CLK _23716_/D VGND VGND VPWR VPWR _23716_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11730_ _16080_/A VGND VGND VPWR VPWR _12156_/A sky130_fd_sc_hd__buf_2
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20372__A1 _17957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20928_ _20782_/X _20927_/X _11519_/A _20789_/X VGND VGND VPWR VPWR _20928_/X sky130_fd_sc_hd__o22a_4
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20638__A _20638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23014__A _22949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _15457_/A VGND VGND VPWR VPWR _14369_/A sky130_fd_sc_hd__buf_2
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23647_ _23679_/CLK _21792_/X VGND VGND VPWR VPWR _23647_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20859_ _20859_/A VGND VGND VPWR VPWR _20860_/A sky130_fd_sc_hd__buf_2
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14636__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _13400_/A _13400_/B _13400_/C VGND VGND VPWR VPWR _13416_/B sky130_fd_sc_hd__and3_4
XANTENNA__13540__A _12949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ _14366_/A _14380_/B VGND VGND VPWR VPWR _14383_/B sky130_fd_sc_hd__or2_4
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11592_ _11592_/A VGND VGND VPWR VPWR _11592_/X sky130_fd_sc_hd__buf_2
X_23578_ _24090_/CLK _23578_/D VGND VGND VPWR VPWR _14645_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22853__A _22799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ _13475_/A _13331_/B _13331_/C VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__or3_4
Xclkbuf_2_1_0_HCLK clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22529_ _22489_/A VGND VGND VPWR VPWR _22529_/X sky130_fd_sc_hd__buf_2
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ _16066_/A _16048_/X _16050_/C VGND VGND VPWR VPWR _16050_/X sky130_fd_sc_hd__and3_4
XANTENNA__15551__A1 _14480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13262_ _13261_/X VGND VGND VPWR VPWR _13262_/X sky130_fd_sc_hd__buf_2
XFILLER_157_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15001_ _13957_/A _23989_/Q VGND VGND VPWR VPWR _15002_/C sky130_fd_sc_hd__or2_4
X_12213_ _12213_/A VGND VGND VPWR VPWR _15439_/A sky130_fd_sc_hd__buf_2
XANTENNA__11995__A _11943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15467__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13193_ _11668_/A VGND VGND VPWR VPWR _15517_/A sky130_fd_sc_hd__buf_2
XFILLER_151_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12144_ _12168_/A _12142_/X _12144_/C VGND VGND VPWR VPWR _12144_/X sky130_fd_sc_hd__and3_4
XANTENNA__15186__B _15122_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19740_ _19740_/A _19808_/A VGND VGND VPWR VPWR _19741_/B sky130_fd_sc_hd__and2_4
X_16952_ _17702_/A VGND VGND VPWR VPWR _17675_/A sky130_fd_sc_hd__inv_2
X_12075_ _11984_/X _12074_/X VGND VGND VPWR VPWR _12075_/X sky130_fd_sc_hd__and2_4
XFILLER_110_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15903_ _15903_/A _15833_/B VGND VGND VPWR VPWR _15905_/B sky130_fd_sc_hd__or2_4
X_19671_ HRDATA[25] VGND VGND VPWR VPWR _20422_/B sky130_fd_sc_hd__buf_2
X_16883_ _16831_/A _16882_/X _16831_/A _16882_/X VGND VGND VPWR VPWR _16884_/D sky130_fd_sc_hd__a2bb2o_4
X_18622_ _24475_/Q VGND VGND VPWR VPWR _18622_/Y sky130_fd_sc_hd__inv_2
X_15834_ _12895_/A _15834_/B VGND VGND VPWR VPWR _15834_/X sky130_fd_sc_hd__or2_4
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18553_ _18553_/A _18148_/B VGND VGND VPWR VPWR _18553_/Y sky130_fd_sc_hd__nand2_4
XFILLER_46_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12977_ _12977_/A _12977_/B _12977_/C VGND VGND VPWR VPWR _12978_/C sky130_fd_sc_hd__and3_4
X_15765_ _11689_/X _15761_/X _15764_/X VGND VGND VPWR VPWR _15765_/X sky130_fd_sc_hd__or3_4
XANTENNA__17359__A2 _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17504_ _17504_/A VGND VGND VPWR VPWR _18336_/B sky130_fd_sc_hd__inv_2
XANTENNA__19402__A _19402_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11928_ _11928_/A VGND VGND VPWR VPWR _11929_/A sky130_fd_sc_hd__inv_2
X_14716_ _14325_/A _14716_/B VGND VGND VPWR VPWR _14718_/B sky130_fd_sc_hd__or2_4
X_15696_ _13170_/A _15696_/B _15695_/X VGND VGND VPWR VPWR _15700_/B sky130_fd_sc_hd__and3_4
X_18484_ _18376_/A _17445_/B VGND VGND VPWR VPWR _18484_/Y sky130_fd_sc_hd__nor2_4
XFILLER_61_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17435_ _17635_/B VGND VGND VPWR VPWR _17435_/Y sky130_fd_sc_hd__inv_2
X_14647_ _15595_/A VGND VGND VPWR VPWR _14647_/X sky130_fd_sc_hd__buf_2
X_11859_ _11625_/A VGND VGND VPWR VPWR _14012_/A sky130_fd_sc_hd__buf_2
XANTENNA__14546__A _11813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22104__A2 _22099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13450__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17366_ _18415_/A VGND VGND VPWR VPWR _17396_/A sky130_fd_sc_hd__inv_2
X_14578_ _14296_/A _23450_/Q VGND VGND VPWR VPWR _14578_/X sky130_fd_sc_hd__or2_4
XANTENNA__21312__B1 _15146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19105_ _24378_/Q VGND VGND VPWR VPWR _19105_/Y sky130_fd_sc_hd__inv_2
X_13529_ _13529_/A _13529_/B _13529_/C VGND VGND VPWR VPWR _13530_/C sky130_fd_sc_hd__and3_4
X_16317_ _11727_/A VGND VGND VPWR VPWR _16318_/A sky130_fd_sc_hd__buf_2
XFILLER_174_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17297_ _17297_/A _17297_/B VGND VGND VPWR VPWR _17297_/X sky130_fd_sc_hd__and2_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16248_ _16157_/A _16248_/B VGND VGND VPWR VPWR _16248_/X sky130_fd_sc_hd__or2_4
XFILLER_118_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23065__B1 _22929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19036_ _24390_/Q VGND VGND VPWR VPWR _19036_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15377__A _15377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16179_ _16210_/A _16179_/B _16179_/C VGND VGND VPWR VPWR _16179_/X sky130_fd_sc_hd__and3_4
XANTENNA__23182__CLK _23246_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21615__B2 _21610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21091__A2 _21090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19938_ _19920_/X VGND VGND VPWR VPWR _19938_/X sky130_fd_sc_hd__buf_2
XFILLER_102_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21918__A2 _21916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19869_ _19879_/D _19868_/X _19665_/A VGND VGND VPWR VPWR _19869_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22003__A _22010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18795__A1 _16523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21900_ _21821_/X _21895_/X _16413_/B _21899_/X VGND VGND VPWR VPWR _21900_/X sky130_fd_sc_hd__o22a_4
X_22880_ _22845_/A _22880_/B VGND VGND VPWR VPWR HWDATA[24] sky130_fd_sc_hd__nor2_4
XANTENNA__16001__A _15969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22938__A _18643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24230__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21831_ _20486_/A VGND VGND VPWR VPWR _21831_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15840__A _12878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21762_ _21791_/A VGND VGND VPWR VPWR _21770_/A sky130_fd_sc_hd__buf_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_68_0_HCLK clkbuf_6_34_0_HCLK/X VGND VGND VPWR VPWR _24182_/CLK sky130_fd_sc_hd__clkbuf_1
X_23501_ _23501_/CLK _22055_/X VGND VGND VPWR VPWR _23501_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20713_ _20713_/A VGND VGND VPWR VPWR _20713_/Y sky130_fd_sc_hd__inv_2
X_24481_ _24134_/CLK _18498_/X HRESETn VGND VGND VPWR VPWR _20071_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14456__A _12455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21693_ _21580_/X _21691_/X _13768_/B _21688_/X VGND VGND VPWR VPWR _21693_/X sky130_fd_sc_hd__o22a_4
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23432_ _23496_/CLK _22196_/X VGND VGND VPWR VPWR _13105_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20644_ _20273_/A VGND VGND VPWR VPWR _20644_/X sky130_fd_sc_hd__buf_2
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23363_ _23908_/CLK _23363_/D VGND VGND VPWR VPWR _15853_/B sky130_fd_sc_hd__dfxtp_4
X_20575_ _20575_/A VGND VGND VPWR VPWR _20575_/X sky130_fd_sc_hd__buf_2
XANTENNA__21854__B2 _21846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16671__A _16659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22314_ _22156_/X _22308_/X _14487_/B _22312_/X VGND VGND VPWR VPWR _22314_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23294_ _23294_/CLK _23294_/D VGND VGND VPWR VPWR _13624_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20409__A2 _20847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15287__A _14269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22245_ _22122_/X _22244_/X _23401_/Q _22241_/X VGND VGND VPWR VPWR _22245_/X sky130_fd_sc_hd__o22a_4
XFILLER_3_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12704__A _12704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22176_ _22176_/A VGND VGND VPWR VPWR _22184_/A sky130_fd_sc_hd__buf_2
XANTENNA__23675__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21127_ _20938_/X _21125_/X _14716_/B _21122_/X VGND VGND VPWR VPWR _21127_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23009__A _22949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18235__B1 _18168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21058_ _20633_/X _21052_/X _24069_/Q _21056_/X VGND VGND VPWR VPWR _21058_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15734__B _23940_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12900_ _12873_/A _12900_/B _12900_/C VGND VGND VPWR VPWR _12904_/B sky130_fd_sc_hd__and3_4
XFILLER_98_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20009_ _18105_/X _20007_/X _20008_/Y _19994_/X VGND VGND VPWR VPWR _20009_/X sky130_fd_sc_hd__o22a_4
X_13880_ _14335_/A _13871_/X _13879_/X VGND VGND VPWR VPWR _13894_/B sky130_fd_sc_hd__or3_4
XANTENNA__21790__B1 _23648_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12831_ _13377_/A _12831_/B _12830_/X VGND VGND VPWR VPWR _12831_/X sky130_fd_sc_hd__and3_4
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15750__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15550_ _14450_/A _15549_/X VGND VGND VPWR VPWR _15550_/X sky130_fd_sc_hd__and2_4
X_12762_ _12762_/A VGND VGND VPWR VPWR _12775_/A sky130_fd_sc_hd__buf_2
XFILLER_55_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21471__B _21370_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14540_/A _14499_/X _14500_/X VGND VGND VPWR VPWR _14505_/B sky130_fd_sc_hd__and3_4
X_11713_ _11712_/X VGND VGND VPWR VPWR _11714_/A sky130_fd_sc_hd__buf_2
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _12626_/A _15481_/B VGND VGND VPWR VPWR _15481_/X sky130_fd_sc_hd__or2_4
XANTENNA__24300__CLK _24302_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12693_ _12693_/A _12774_/B VGND VGND VPWR VPWR _12693_/X sky130_fd_sc_hd__or2_4
XFILLER_43_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _12531_/A _24027_/Q VGND VGND VPWR VPWR _14432_/X sky130_fd_sc_hd__or2_4
X_17220_ _12077_/X _17203_/X _17151_/X _17219_/Y VGND VGND VPWR VPWR _17220_/X sky130_fd_sc_hd__o22a_4
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11643_/Y VGND VGND VPWR VPWR _11644_/X sky130_fd_sc_hd__buf_2
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14085__B _14084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17151_ _12028_/X VGND VGND VPWR VPWR _17151_/X sky130_fd_sc_hd__buf_2
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _12583_/A _14363_/B VGND VGND VPWR VPWR _14363_/X sky130_fd_sc_hd__or2_4
XFILLER_7_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11575_ _11575_/A IRQ[24] VGND VGND VPWR VPWR _11575_/X sky130_fd_sc_hd__and2_4
XFILLER_156_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16102_ _16109_/A _16102_/B VGND VGND VPWR VPWR _16103_/C sky130_fd_sc_hd__or2_4
XFILLER_122_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13314_ _13318_/A _13312_/X _13314_/C VGND VGND VPWR VPWR _13314_/X sky130_fd_sc_hd__and3_4
X_17082_ _17075_/X _17082_/B VGND VGND VPWR VPWR _17083_/B sky130_fd_sc_hd__or2_4
X_14294_ _15022_/A VGND VGND VPWR VPWR _14301_/A sky130_fd_sc_hd__buf_2
XFILLER_122_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16033_ _16033_/A VGND VGND VPWR VPWR _16046_/A sky130_fd_sc_hd__buf_2
X_13245_ _13252_/A _23111_/Q VGND VGND VPWR VPWR _13247_/B sky130_fd_sc_hd__or2_4
XFILLER_170_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12614__A _12977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17277__A1 _17273_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13176_ _13332_/A _23495_/Q VGND VGND VPWR VPWR _13176_/X sky130_fd_sc_hd__or2_4
XFILLER_124_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22270__B2 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21927__A _21906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11561__A2 IRQ[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12127_ _12127_/A _24051_/Q VGND VGND VPWR VPWR _12129_/B sky130_fd_sc_hd__or2_4
XFILLER_151_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17984_ _17824_/X _17982_/X _17813_/X _17983_/X VGND VGND VPWR VPWR _17984_/Y sky130_fd_sc_hd__a22oi_4
X_19723_ _19696_/X _19721_/Y _20866_/B _19573_/A VGND VGND VPWR VPWR _19723_/X sky130_fd_sc_hd__a2bb2o_4
X_16935_ _16935_/A VGND VGND VPWR VPWR _16935_/X sky130_fd_sc_hd__buf_2
X_12058_ _12058_/A _23699_/Q VGND VGND VPWR VPWR _12061_/B sky130_fd_sc_hd__or2_4
XANTENNA__22022__B2 _22021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13445__A _13468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19974__B1 _18009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19654_ _19596_/X _19778_/B _19888_/B VGND VGND VPWR VPWR _19655_/D sky130_fd_sc_hd__o21a_4
X_16866_ _15116_/X VGND VGND VPWR VPWR _16866_/X sky130_fd_sc_hd__buf_2
XFILLER_168_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22758__A SYSTICKCLKDIV[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18605_ _17311_/Y _18604_/X VGND VGND VPWR VPWR _18605_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21662__A _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15817_ _11970_/A _15816_/X VGND VGND VPWR VPWR _15817_/X sky130_fd_sc_hd__and2_4
X_19585_ _24171_/Q _19457_/A HRDATA[23] _19454_/A VGND VGND VPWR VPWR _19585_/X sky130_fd_sc_hd__o22a_4
X_16797_ _16635_/A _16797_/B _16797_/C VGND VGND VPWR VPWR _16801_/B sky130_fd_sc_hd__and3_4
X_18536_ _18111_/A _18364_/X _18533_/Y _18026_/X _22961_/B VGND VGND VPWR VPWR _18536_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_80_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15748_ _11739_/A _15746_/X _15747_/X VGND VGND VPWR VPWR _15748_/X sky130_fd_sc_hd__and3_4
XFILLER_34_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18467_ _18198_/A VGND VGND VPWR VPWR _18467_/X sky130_fd_sc_hd__buf_2
X_15679_ _12702_/A _15735_/B VGND VGND VPWR VPWR _15679_/X sky130_fd_sc_hd__or2_4
XANTENNA__14276__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17418_ _17418_/A _17418_/B VGND VGND VPWR VPWR _17418_/X sky130_fd_sc_hd__and2_4
X_18398_ _18356_/X _18395_/X _18396_/X _18397_/X VGND VGND VPWR VPWR _18398_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22493__A _22489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17349_ _15382_/B _17323_/Y _18689_/A _17348_/X VGND VGND VPWR VPWR _17350_/B sky130_fd_sc_hd__o22a_4
XFILLER_119_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16922__C _16922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20360_ _20360_/A VGND VGND VPWR VPWR _21532_/A sky130_fd_sc_hd__buf_2
X_19019_ _19017_/Y _19018_/Y _11535_/X VGND VGND VPWR VPWR _19019_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20291_ _20269_/X _20285_/X _20343_/A _20290_/X VGND VGND VPWR VPWR _20292_/C sky130_fd_sc_hd__a211o_4
XANTENNA__12524__A _12882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21064__A2 _21059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22030_ _21872_/X _22024_/X _14485_/B _22028_/X VGND VGND VPWR VPWR _22030_/X sky130_fd_sc_hd__o22a_4
XFILLER_161_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22261__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24482__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15835__A _12873_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22013__B2 _22007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23981_ _24045_/CLK _21200_/X VGND VGND VPWR VPWR _23981_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13355__A _13399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22564__A2 _22558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_31_0_HCLK clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22932_ _18657_/X _22930_/Y _19319_/X _22931_/X VGND VGND VPWR VPWR _22933_/C sky130_fd_sc_hd__a211o_4
XFILLER_96_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24323__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22863_ _14767_/Y _22848_/X _22815_/X VGND VGND VPWR VPWR _22863_/X sky130_fd_sc_hd__o21a_4
XFILLER_84_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22316__A2 _22315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16666__A _16678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15570__A _14430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21814_ _21808_/A VGND VGND VPWR VPWR _21839_/A sky130_fd_sc_hd__buf_2
XFILLER_71_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22794_ _24125_/Q VGND VGND VPWR VPWR _22794_/Y sky130_fd_sc_hd__inv_2
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21745_ _21724_/A VGND VGND VPWR VPWR _21745_/X sky130_fd_sc_hd__buf_2
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13090__A _13090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18940__A1 _15251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24473__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11603__A _11603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24464_ _23379_/CLK _24464_/D HRESETn VGND VGND VPWR VPWR _24464_/Q sky130_fd_sc_hd__dfrtp_4
X_21676_ _21551_/X _21670_/X _23722_/Q _21674_/X VGND VGND VPWR VPWR _23722_/D sky130_fd_sc_hd__o22a_4
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23415_ _23864_/CLK _22219_/X VGND VGND VPWR VPWR _15166_/B sky130_fd_sc_hd__dfxtp_4
X_20627_ _20626_/X VGND VGND VPWR VPWR _20627_/Y sky130_fd_sc_hd__inv_2
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24395_ _24428_/CLK _24395_/D HRESETn VGND VGND VPWR VPWR _19007_/A sky130_fd_sc_hd__dfstp_4
XFILLER_138_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23346_ _23204_/CLK _23346_/D VGND VGND VPWR VPWR _23346_/Q sky130_fd_sc_hd__dfxtp_4
X_20558_ _20558_/A VGND VGND VPWR VPWR _21268_/A sky130_fd_sc_hd__buf_2
XFILLER_137_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14633__B _14633_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23277_ _23533_/CLK _22429_/X VGND VGND VPWR VPWR _16090_/B sky130_fd_sc_hd__dfxtp_4
X_20489_ _20257_/X VGND VGND VPWR VPWR _20501_/A sky130_fd_sc_hd__buf_2
XFILLER_98_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12434__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13030_ _12570_/A _13028_/X _13029_/X VGND VGND VPWR VPWR _13030_/X sky130_fd_sc_hd__and3_4
XFILLER_156_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21055__A2 _21052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18456__B1 _18027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22228_ _22222_/Y _22227_/X _22095_/X _22227_/X VGND VGND VPWR VPWR _23412_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22252__B2 _22248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15745__A _12778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22159_ _22147_/A VGND VGND VPWR VPWR _22159_/X sky130_fd_sc_hd__buf_2
XFILLER_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22004__B2 _22000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14981_ _11812_/A _14965_/X _14980_/X VGND VGND VPWR VPWR _14981_/X sky130_fd_sc_hd__or3_4
XFILLER_87_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16720_ _16700_/A _23921_/Q VGND VGND VPWR VPWR _16722_/B sky130_fd_sc_hd__or2_4
X_13932_ _13710_/A _23709_/Q VGND VGND VPWR VPWR _13932_/X sky130_fd_sc_hd__or2_4
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21482__A _21482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16651_ _16675_/A _16646_/X _16651_/C VGND VGND VPWR VPWR _16652_/C sky130_fd_sc_hd__or3_4
X_13863_ _11854_/A _11628_/A _13830_/X _11605_/A _13862_/X VGND VGND VPWR VPWR _13863_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13048__A2 _11629_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22307__A2 _22301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12814_ _13343_/A _12812_/X _12814_/C VGND VGND VPWR VPWR _12815_/C sky130_fd_sc_hd__and3_4
X_15602_ _15611_/A _15602_/B VGND VGND VPWR VPWR _15602_/X sky130_fd_sc_hd__or2_4
X_19370_ _19369_/X _18596_/X _19369_/X _24252_/Q VGND VGND VPWR VPWR _19370_/X sky130_fd_sc_hd__a2bb2o_4
X_13794_ _13952_/A VGND VGND VPWR VPWR _14574_/A sky130_fd_sc_hd__buf_2
X_16582_ _16554_/X _16665_/B VGND VGND VPWR VPWR _16583_/C sky130_fd_sc_hd__or2_4
XFILLER_15_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18321_ _18198_/X _18464_/B _18265_/X _18320_/X VGND VGND VPWR VPWR _18321_/X sky130_fd_sc_hd__a211o_4
XFILLER_76_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12745_ _12745_/A _12743_/X _12745_/C VGND VGND VPWR VPWR _12745_/X sky130_fd_sc_hd__and3_4
X_15533_ _12304_/A _15533_/B VGND VGND VPWR VPWR _15533_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_51_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR _23852_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18931__A1 _17153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15464_ _13774_/A _15462_/X _15464_/C VGND VGND VPWR VPWR _15464_/X sky130_fd_sc_hd__and3_4
X_18252_ _17686_/A _18251_/Y VGND VGND VPWR VPWR _18253_/A sky130_fd_sc_hd__or2_4
X_12676_ _12676_/A _12676_/B _12676_/C VGND VGND VPWR VPWR _12677_/C sky130_fd_sc_hd__or3_4
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _15389_/A VGND VGND VPWR VPWR _14415_/Y sky130_fd_sc_hd__inv_2
X_17203_ _17112_/X _17190_/Y _17137_/X _17202_/Y VGND VGND VPWR VPWR _17203_/X sky130_fd_sc_hd__o22a_4
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _11627_/A VGND VGND VPWR VPWR _11628_/A sky130_fd_sc_hd__buf_2
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15395_ _15395_/A _15458_/B VGND VGND VPWR VPWR _15395_/X sky130_fd_sc_hd__or2_4
XANTENNA__21818__B2 _21810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18183_ _17770_/Y _18182_/X _17703_/X VGND VGND VPWR VPWR _18183_/X sky130_fd_sc_hd__o21a_4
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17134_ _15252_/X _17131_/X _17132_/Y _17133_/X VGND VGND VPWR VPWR _17134_/X sky130_fd_sc_hd__o22a_4
X_14346_ _14512_/A _14343_/X _14345_/X VGND VGND VPWR VPWR _14346_/X sky130_fd_sc_hd__and3_4
XANTENNA__21294__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11558_ _11555_/X _11557_/X VGND VGND VPWR VPWR _11558_/X sky130_fd_sc_hd__or2_4
XFILLER_155_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17065_ _17100_/A VGND VGND VPWR VPWR _17188_/A sky130_fd_sc_hd__inv_2
XFILLER_143_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14277_ _14277_/A VGND VGND VPWR VPWR _14310_/A sky130_fd_sc_hd__buf_2
XFILLER_155_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16016_ _16015_/X VGND VGND VPWR VPWR _16016_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21046__A2 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13228_ _12354_/A _13219_/X _13228_/C VGND VGND VPWR VPWR _13229_/C sky130_fd_sc_hd__and3_4
XANTENNA__23990__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18447__B1 _18060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22243__B2 _22241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13159_ _11970_/A _13158_/X VGND VGND VPWR VPWR _13159_/X sky130_fd_sc_hd__and2_4
XFILLER_170_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23220__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17967_ _18150_/A _17641_/A VGND VGND VPWR VPWR _17967_/X sky130_fd_sc_hd__or2_4
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22546__A2 _22544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13175__A _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19706_ _19659_/Y _19665_/B VGND VGND VPWR VPWR _19787_/A sky130_fd_sc_hd__and2_4
XFILLER_78_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16918_ _16918_/A VGND VGND VPWR VPWR _16918_/X sky130_fd_sc_hd__buf_2
X_17898_ _11642_/X _17897_/X _19988_/A _11642_/X VGND VGND VPWR VPWR _24498_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19637_ _19703_/A HRDATA[10] VGND VGND VPWR VPWR _19637_/X sky130_fd_sc_hd__and2_4
X_16849_ _14266_/B _16848_/X _14263_/X VGND VGND VPWR VPWR _16849_/X sky130_fd_sc_hd__o21a_4
XFILLER_92_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13903__A _14348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19568_ _20339_/B _19573_/A _19519_/X HRDATA[13] VGND VGND VPWR VPWR _19568_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_94_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18519_ _17798_/A VGND VGND VPWR VPWR _18519_/X sky130_fd_sc_hd__buf_2
XFILLER_22_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19797__A _19797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19499_ _19499_/A VGND VGND VPWR VPWR _19528_/B sky130_fd_sc_hd__buf_2
XANTENNA__12519__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18922__A1 _13567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21530_ _21542_/A VGND VGND VPWR VPWR _21530_/X sky130_fd_sc_hd__buf_2
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21461_ _21302_/X _21455_/X _14460_/B _21459_/X VGND VGND VPWR VPWR _21461_/X sky130_fd_sc_hd__o22a_4
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23200_ _23203_/CLK _23200_/D VGND VGND VPWR VPWR _23200_/Q sky130_fd_sc_hd__dfxtp_4
X_20412_ _24271_/Q _20305_/X _20411_/X VGND VGND VPWR VPWR _20412_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17110__A _17109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24180_ _24182_/CLK _24180_/D HRESETn VGND VGND VPWR VPWR _20241_/A sky130_fd_sc_hd__dfrtp_4
X_21392_ _21268_/X _21391_/X _23881_/Q _21388_/X VGND VGND VPWR VPWR _23881_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23131_ _24096_/CLK _22678_/X VGND VGND VPWR VPWR _14523_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16161__A1 _11973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20343_ _20343_/A VGND VGND VPWR VPWR _20343_/X sky130_fd_sc_hd__buf_2
X_23062_ _23036_/X _17904_/X _23048_/X _23061_/X VGND VGND VPWR VPWR _23063_/A sky130_fd_sc_hd__a211o_4
X_20274_ _20274_/A VGND VGND VPWR VPWR _20495_/A sky130_fd_sc_hd__inv_2
XANTENNA__20471__A _20282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22013_ _21843_/X _22010_/X _23527_/Q _22007_/X VGND VGND VPWR VPWR _22013_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15565__A _12186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20796__A1 _20662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23964_ _23592_/CLK _23964_/D VGND VGND VPWR VPWR _23964_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22915_ _18717_/X _22930_/A _22914_/X VGND VGND VPWR VPWR _22915_/X sky130_fd_sc_hd__o21a_4
XFILLER_112_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23895_ _23862_/CLK _23895_/D VGND VGND VPWR VPWR _15155_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16396__A _16011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14909__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13813__A _15405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22846_ _18780_/X _22846_/B VGND VGND VPWR VPWR _22846_/X sky130_fd_sc_hd__or2_4
XFILLER_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22777_ _22777_/A _22778_/B _22793_/A VGND VGND VPWR VPWR _24119_/D sky130_fd_sc_hd__and3_4
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22170__B1 _23445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _12530_/A VGND VGND VPWR VPWR _12531_/A sky130_fd_sc_hd__buf_2
Xclkbuf_6_38_0_HCLK clkbuf_6_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_77_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21728_ _21553_/X _21727_/X _23689_/Q _21724_/X VGND VGND VPWR VPWR _21728_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19500__A _19624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20720__A1 _20635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20720__B2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12461_ _12461_/A VGND VGND VPWR VPWR _12881_/A sky130_fd_sc_hd__buf_2
X_24447_ _24445_/CLK _18820_/X HRESETn VGND VGND VPWR VPWR _11567_/A sky130_fd_sc_hd__dfrtp_4
X_21659_ _21674_/A VGND VGND VPWR VPWR _21667_/A sky130_fd_sc_hd__buf_2
XFILLER_71_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24219__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14200_ _14200_/A _23295_/Q VGND VGND VPWR VPWR _14201_/C sky130_fd_sc_hd__or2_4
XFILLER_71_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15180_ _13953_/A _15180_/B VGND VGND VPWR VPWR _15181_/C sky130_fd_sc_hd__or2_4
X_12392_ _12407_/A _12392_/B VGND VGND VPWR VPWR _12394_/B sky130_fd_sc_hd__or2_4
XANTENNA__15459__B _23746_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24378_ _24382_/CLK _18937_/X HRESETn VGND VGND VPWR VPWR _24378_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_166_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14363__B _14363_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14131_ _14131_/A _23455_/Q VGND VGND VPWR VPWR _14132_/C sky130_fd_sc_hd__or2_4
XFILLER_126_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23329_ _23744_/CLK _22341_/X VGND VGND VPWR VPWR _15539_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_137_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24333__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21477__A _21506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14062_ _11660_/A _14062_/B VGND VGND VPWR VPWR _14062_/X sky130_fd_sc_hd__or2_4
XFILLER_4_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13013_ _12540_/A _13013_/B VGND VGND VPWR VPWR _13013_/X sky130_fd_sc_hd__or2_4
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18870_ _18838_/X VGND VGND VPWR VPWR _18870_/X sky130_fd_sc_hd__buf_2
X_17821_ _17816_/X _17121_/X _17817_/X _17138_/X VGND VGND VPWR VPWR _17821_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12611__B _12611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17752_ _17751_/X VGND VGND VPWR VPWR _17752_/X sky130_fd_sc_hd__buf_2
X_14964_ _15369_/A _14960_/X _14963_/X VGND VGND VPWR VPWR _14964_/X sky130_fd_sc_hd__or3_4
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16703_ _16592_/A _16703_/B _16702_/X VGND VGND VPWR VPWR _16703_/X sky130_fd_sc_hd__or3_4
XANTENNA__21200__A2 _21198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13915_ _14375_/A _13913_/X _13915_/C VGND VGND VPWR VPWR _13920_/B sky130_fd_sc_hd__and3_4
XFILLER_130_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17683_ _17683_/A _17683_/B VGND VGND VPWR VPWR _17775_/C sky130_fd_sc_hd__or2_4
XFILLER_47_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14895_ _14131_/A _14895_/B VGND VGND VPWR VPWR _14896_/C sky130_fd_sc_hd__or2_4
XFILLER_63_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22101__A _20360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19422_ _19418_/X _18537_/Y _19421_/X _24223_/Q VGND VGND VPWR VPWR _24223_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16634_ _16656_/A _16632_/X _16633_/X VGND VGND VPWR VPWR _16642_/B sky130_fd_sc_hd__and3_4
X_13846_ _13639_/A _24093_/Q VGND VGND VPWR VPWR _13847_/C sky130_fd_sc_hd__or2_4
XFILLER_62_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19353_ _19350_/X _18327_/X _19350_/X _24263_/Q VGND VGND VPWR VPWR _19353_/X sky130_fd_sc_hd__a2bb2o_4
X_13777_ _12621_/X _13775_/X _13776_/X VGND VGND VPWR VPWR _13777_/X sky130_fd_sc_hd__and3_4
XFILLER_16_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16565_ _16593_/A _16638_/B VGND VGND VPWR VPWR _16567_/B sky130_fd_sc_hd__or2_4
XANTENNA__12339__A _12338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18904__A1 _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22700__A2 _22694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18304_ _17697_/A _18303_/X _17697_/A _18303_/X VGND VGND VPWR VPWR _18304_/X sky130_fd_sc_hd__a2bb2o_4
X_15516_ _12978_/A _15500_/X _15515_/X VGND VGND VPWR VPWR _15516_/X sky130_fd_sc_hd__or3_4
XFILLER_43_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12728_ _13279_/A _12817_/B VGND VGND VPWR VPWR _12729_/C sky130_fd_sc_hd__or2_4
X_19284_ _24295_/Q _19244_/B _19283_/Y VGND VGND VPWR VPWR _19284_/X sky130_fd_sc_hd__o21a_4
X_16496_ _16370_/X _16492_/X _16495_/X VGND VGND VPWR VPWR _16504_/B sky130_fd_sc_hd__or3_4
XANTENNA__20556__A _20535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18235_ _18095_/X _17459_/A _18233_/X _18168_/X _18234_/Y VGND VGND VPWR VPWR _18235_/X
+ sky130_fd_sc_hd__a32o_4
X_12659_ _12659_/A _12653_/X _12659_/C VGND VGND VPWR VPWR _12660_/C sky130_fd_sc_hd__or3_4
X_15447_ _15447_/A _15505_/B VGND VGND VPWR VPWR _15448_/C sky130_fd_sc_hd__or2_4
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14554__A _14270_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18026__A _24212_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21267__A2 _21257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18166_ _17598_/Y _18166_/B VGND VGND VPWR VPWR _18167_/B sky130_fd_sc_hd__and2_4
XFILLER_172_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15378_ _15378_/A _15378_/B _15378_/C VGND VGND VPWR VPWR _15378_/X sky130_fd_sc_hd__or3_4
XFILLER_50_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17117_ _15382_/B _17115_/X _16821_/B _17116_/X VGND VGND VPWR VPWR _17117_/X sky130_fd_sc_hd__o22a_4
X_14329_ _14329_/A _14400_/B VGND VGND VPWR VPWR _14330_/C sky130_fd_sc_hd__or2_4
X_18097_ _18097_/A VGND VGND VPWR VPWR _18097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12074__A _11939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17048_ _17048_/A _17297_/B VGND VGND VPWR VPWR _17049_/A sky130_fd_sc_hd__or2_4
XANTENNA__22216__B2 _22212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12802__A _13562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21975__B1 _23551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12521__B _23467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18999_ _18993_/X _18998_/X _18993_/X _18994_/A VGND VGND VPWR VPWR _18999_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20961_ _20940_/A _19773_/X VGND VGND VPWR VPWR _20961_/X sky130_fd_sc_hd__or2_4
XFILLER_38_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22700_ _21824_/A _22694_/X _16300_/B _22698_/X VGND VGND VPWR VPWR _22700_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23680_ _24096_/CLK _23680_/D VGND VGND VPWR VPWR _23680_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20892_ _20892_/A VGND VGND VPWR VPWR _20892_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22631_ _22476_/X _22629_/X _14798_/B _22626_/X VGND VGND VPWR VPWR _23161_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12249__A _14450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22562_ _22555_/A VGND VGND VPWR VPWR _22562_/X sky130_fd_sc_hd__buf_2
XANTENNA__20466__A _20231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24301_ _24302_/CLK _19272_/X HRESETn VGND VGND VPWR VPWR _19250_/A sky130_fd_sc_hd__dfrtp_4
X_21513_ _21506_/A VGND VGND VPWR VPWR _21513_/X sky130_fd_sc_hd__buf_2
X_22493_ _22489_/A VGND VGND VPWR VPWR _22508_/A sky130_fd_sc_hd__buf_2
X_24232_ _24127_/CLK _19409_/X HRESETn VGND VGND VPWR VPWR _24232_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21258__A2 _21257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21444_ _21273_/X _21441_/X _23847_/Q _21438_/X VGND VGND VPWR VPWR _23847_/D sky130_fd_sc_hd__o22a_4
XFILLER_148_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22455__B2 _22445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23266__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24163_ _24134_/CLK _24163_/D HRESETn VGND VGND VPWR VPWR _24163_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21375_ _21369_/Y _21374_/X _21241_/X _21374_/X VGND VGND VPWR VPWR _23892_/D sky130_fd_sc_hd__a2bb2o_4
X_23114_ _23852_/CLK _23114_/D VGND VGND VPWR VPWR _12824_/B sky130_fd_sc_hd__dfxtp_4
X_20326_ _20315_/X _20324_/X _11544_/D _20325_/X VGND VGND VPWR VPWR _20326_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21297__A _20841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24094_ _23880_/CLK _20820_/X VGND VGND VPWR VPWR _24094_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22207__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23045_ _23051_/A _23043_/Y _23045_/C VGND VGND VPWR VPWR _23045_/X sky130_fd_sc_hd__and3_4
XANTENNA__15295__A _14272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13808__A _12485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20257_ _20257_/A VGND VGND VPWR VPWR _20257_/X sky130_fd_sc_hd__buf_2
XFILLER_66_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21430__A2 _21427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20188_ _20188_/A _20188_/B VGND VGND VPWR VPWR _20188_/X sky130_fd_sc_hd__or2_4
XFILLER_48_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11961_ _12105_/A _11804_/B VGND VGND VPWR VPWR _11961_/X sky130_fd_sc_hd__or2_4
X_23947_ _23467_/CLK _23947_/D VGND VGND VPWR VPWR _12618_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21194__B2 _21188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13543__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13700_ _13700_/A VGND VGND VPWR VPWR _13710_/A sky130_fd_sc_hd__buf_2
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14680_ _14680_/A _14680_/B _14680_/C VGND VGND VPWR VPWR _14681_/C sky130_fd_sc_hd__and3_4
X_23878_ _23397_/CLK _21396_/X VGND VGND VPWR VPWR _13405_/B sky130_fd_sc_hd__dfxtp_4
X_11892_ _11891_/X VGND VGND VPWR VPWR _16711_/A sky130_fd_sc_hd__buf_2
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21760__A _21767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13631_ _14329_/A VGND VGND VPWR VPWR _13632_/A sky130_fd_sc_hd__buf_2
X_22829_ _22819_/X _17319_/Y VGND VGND VPWR VPWR _22829_/X sky130_fd_sc_hd__or2_4
XFILLER_53_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18772__C _18411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13562_ _13562_/A _13562_/B _13562_/C VGND VGND VPWR VPWR _13563_/C sky130_fd_sc_hd__and3_4
XANTENNA__21497__A2 _21492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16350_ _16333_/A _16282_/B VGND VGND VPWR VPWR _16350_/X sky130_fd_sc_hd__or2_4
XFILLER_160_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12513_ _12513_/A VGND VGND VPWR VPWR _12514_/A sky130_fd_sc_hd__buf_2
XFILLER_160_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15301_ _14296_/A _23640_/Q VGND VGND VPWR VPWR _15302_/C sky130_fd_sc_hd__or2_4
X_16281_ _15952_/A _16279_/X _16280_/X VGND VGND VPWR VPWR _16281_/X sky130_fd_sc_hd__and3_4
XANTENNA__11998__A _11963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13493_ _12955_/A VGND VGND VPWR VPWR _15903_/A sky130_fd_sc_hd__buf_2
XANTENNA__14374__A _13229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20095__B _17817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18020_ _18019_/X VGND VGND VPWR VPWR _18020_/X sky130_fd_sc_hd__buf_2
XFILLER_12_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15232_ _14769_/A _15228_/X _15232_/C VGND VGND VPWR VPWR _15232_/X sky130_fd_sc_hd__or3_4
X_12444_ _12444_/A VGND VGND VPWR VPWR _12445_/A sky130_fd_sc_hd__buf_2
XANTENNA__22446__B2 _22445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22591__A _22598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24191__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20457__B1 _20638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15163_ _15294_/A _15227_/B VGND VGND VPWR VPWR _15163_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_3_0_0_HCLK_A clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12375_ _12923_/A VGND VGND VPWR VPWR _15851_/A sky130_fd_sc_hd__buf_2
X_14114_ _14114_/A VGND VGND VPWR VPWR _14149_/A sky130_fd_sc_hd__buf_2
XFILLER_125_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19971_ _17057_/B _19970_/Y VGND VGND VPWR VPWR _19971_/X sky130_fd_sc_hd__or2_4
X_15094_ _15078_/A _15092_/X _15093_/X VGND VGND VPWR VPWR _15094_/X sky130_fd_sc_hd__and3_4
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15917__B _15916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13718__A _15372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18922_ _13567_/X _18920_/X _24389_/Q _18921_/X VGND VGND VPWR VPWR _18922_/X sky130_fd_sc_hd__o22a_4
X_14045_ _11660_/A _22342_/A VGND VGND VPWR VPWR _14045_/X sky130_fd_sc_hd__or2_4
XFILLER_84_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18853_ _16240_/X _18849_/X _20448_/A _18850_/X VGND VGND VPWR VPWR _24429_/D sky130_fd_sc_hd__o22a_4
XFILLER_67_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17804_ _17804_/A VGND VGND VPWR VPWR _17804_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18784_ _18837_/A _18784_/B VGND VGND VPWR VPWR _18785_/A sky130_fd_sc_hd__or2_4
X_15996_ _15969_/A _24110_/Q VGND VGND VPWR VPWR _15997_/C sky130_fd_sc_hd__or2_4
XFILLER_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17735_ _17735_/A _17734_/X VGND VGND VPWR VPWR _17760_/B sky130_fd_sc_hd__or2_4
X_14947_ _14786_/A _14945_/X _14947_/C VGND VGND VPWR VPWR _14947_/X sky130_fd_sc_hd__and3_4
XANTENNA__14549__A _14547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13453__A _13453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17666_ _17669_/A _17567_/X VGND VGND VPWR VPWR _17666_/X sky130_fd_sc_hd__and2_4
X_14878_ _13981_/A _14878_/B VGND VGND VPWR VPWR _14878_/X sky130_fd_sc_hd__and2_4
XFILLER_169_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14268__B _14337_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21670__A _21677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19405_ _19399_/X _19404_/Y _19402_/X _24234_/Q VGND VGND VPWR VPWR _24234_/D sky130_fd_sc_hd__o22a_4
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16617_ _16662_/A _23762_/Q VGND VGND VPWR VPWR _16617_/X sky130_fd_sc_hd__or2_4
XFILLER_23_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24365__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13829_ _15420_/A _13828_/X VGND VGND VPWR VPWR _13829_/X sky130_fd_sc_hd__and2_4
X_17597_ _17572_/X _18113_/B VGND VGND VPWR VPWR _17641_/C sky130_fd_sc_hd__or2_4
XANTENNA__12069__A _16742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19336_ _19325_/X _17785_/X _19335_/X _24275_/Q VGND VGND VPWR VPWR _24275_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21488__A2 _21485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16548_ _16539_/X _16627_/B VGND VGND VPWR VPWR _16549_/C sky130_fd_sc_hd__or2_4
XANTENNA__20286__A _20264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22685__B2 _22648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_21_0_HCLK clkbuf_6_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19267_ _19253_/B VGND VGND VPWR VPWR _19267_/Y sky130_fd_sc_hd__inv_2
X_16479_ _13384_/A VGND VGND VPWR VPWR _16479_/X sky130_fd_sc_hd__buf_2
XFILLER_31_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14284__A _14310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11701__A _11701_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18218_ _18216_/X _18217_/X _18216_/X _18217_/X VGND VGND VPWR VPWR _19404_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19198_ _24322_/Q _19142_/X _19197_/Y VGND VGND VPWR VPWR _24322_/D sky130_fd_sc_hd__o21a_4
XFILLER_129_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18149_ _23038_/B _18148_/X _23038_/B _18148_/X VGND VGND VPWR VPWR _18149_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21160_ _20613_/X _21155_/X _13294_/B _21159_/X VGND VGND VPWR VPWR _24006_/D sky130_fd_sc_hd__o22a_4
XFILLER_85_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14731__B _14731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20111_ _20108_/Y _20109_/Y _20110_/Y _20111_/D VGND VGND VPWR VPWR _20111_/X sky130_fd_sc_hd__and4_4
XFILLER_104_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12532__A _12875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21091_ _20337_/X _21090_/X _24051_/Q _21087_/X VGND VGND VPWR VPWR _21091_/X sky130_fd_sc_hd__o22a_4
XFILLER_113_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20042_ _19950_/X VGND VGND VPWR VPWR _20042_/X sky130_fd_sc_hd__buf_2
XFILLER_113_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15843__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23801_ _23641_/CLK _21515_/X VGND VGND VPWR VPWR _14758_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21993_ _22000_/A VGND VGND VPWR VPWR _21993_/X sky130_fd_sc_hd__buf_2
XFILLER_67_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14459__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23732_ _23764_/CLK _23732_/D VGND VGND VPWR VPWR _21655_/A sky130_fd_sc_hd__dfxtp_4
X_20944_ HRDATA[3] VGND VGND VPWR VPWR _20944_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_103_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR _23587_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21580__A _20819_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _23246_/CLK _21769_/X VGND VGND VPWR VPWR _16297_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20875_ _20943_/A _20870_/X _20874_/X VGND VGND VPWR VPWR _20875_/X sky130_fd_sc_hd__a21o_4
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16674__A _16678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22614_ _22447_/X _22608_/X _13449_/B _22612_/X VGND VGND VPWR VPWR _22614_/X sky130_fd_sc_hd__o22a_4
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20908__B _20908_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21479__A2 _21478_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23594_ _23531_/CLK _21908_/X VGND VGND VPWR VPWR _12790_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22545_ _22412_/X _22544_/X _12124_/B _22541_/X VGND VGND VPWR VPWR _23219_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13810__B _24029_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12707__A _12298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11611__A _17274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22476_ _20937_/A VGND VGND VPWR VPWR _22476_/X sky130_fd_sc_hd__buf_2
XFILLER_108_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24215_ _24248_/CLK _19432_/X HRESETn VGND VGND VPWR VPWR _24215_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21427_ _21441_/A VGND VGND VPWR VPWR _21427_/X sky130_fd_sc_hd__buf_2
XFILLER_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21100__B2 _21094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24146_ _24134_/CLK _24146_/D HRESETn VGND VGND VPWR VPWR _24146_/Q sky130_fd_sc_hd__dfrtp_4
X_12160_ _12122_/A _12158_/X _12159_/X VGND VGND VPWR VPWR _12161_/C sky130_fd_sc_hd__and3_4
XFILLER_136_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21651__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21358_ _21297_/X _21355_/X _13831_/B _21352_/X VGND VGND VPWR VPWR _23901_/D sky130_fd_sc_hd__o22a_4
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13538__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20309_ _20307_/X _20672_/A _20308_/X VGND VGND VPWR VPWR _20309_/X sky130_fd_sc_hd__a21o_4
X_24077_ _24077_/CLK _21047_/X VGND VGND VPWR VPWR _24077_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12091_ _16732_/A _12089_/X _12091_/C VGND VGND VPWR VPWR _12091_/X sky130_fd_sc_hd__and3_4
XANTENNA__12442__A _13955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21289_ _21287_/X _21281_/X _15601_/B _21288_/X VGND VGND VPWR VPWR _23937_/D sky130_fd_sc_hd__o22a_4
XFILLER_150_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13341__A1 _11858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23028_ _23007_/X _16954_/Y _23019_/X _23027_/X VGND VGND VPWR VPWR _23029_/A sky130_fd_sc_hd__a211o_4
XANTENNA__21403__A2 _21398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22600__B2 _22598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15753__A _12762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15850_ _12373_/X _15789_/B VGND VGND VPWR VPWR _15850_/X sky130_fd_sc_hd__or2_4
X_14801_ _14840_/A _14797_/X _14801_/C VGND VGND VPWR VPWR _14810_/B sky130_fd_sc_hd__or3_4
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15781_ _13123_/A _15781_/B _15781_/C VGND VGND VPWR VPWR _15781_/X sky130_fd_sc_hd__and3_4
X_12993_ _12877_/A _12991_/X _12993_/C VGND VGND VPWR VPWR _12994_/C sky130_fd_sc_hd__and3_4
XANTENNA__21167__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13273__A _12559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17520_ _17493_/A _17520_/B VGND VGND VPWR VPWR _17520_/X sky130_fd_sc_hd__or2_4
XFILLER_57_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14732_ _12468_/A _14730_/X _14732_/C VGND VGND VPWR VPWR _14732_/X sky130_fd_sc_hd__and3_4
X_11944_ _11975_/A VGND VGND VPWR VPWR _16744_/A sky130_fd_sc_hd__buf_2
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18783__B _18888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17451_ _17450_/X VGND VGND VPWR VPWR _17451_/Y sky130_fd_sc_hd__inv_2
X_11875_ _16159_/A VGND VGND VPWR VPWR _16145_/A sky130_fd_sc_hd__buf_2
XFILLER_45_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14663_ _14663_/A VGND VGND VPWR VPWR _14682_/A sky130_fd_sc_hd__buf_2
XFILLER_33_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16584__A _16561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16402_ _16401_/X VGND VGND VPWR VPWR _16402_/X sky130_fd_sc_hd__buf_2
X_13614_ _14297_/A VGND VGND VPWR VPWR _15401_/A sky130_fd_sc_hd__buf_2
X_17382_ _15785_/A _17354_/X _17028_/X _17381_/X VGND VGND VPWR VPWR _17383_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22667__B2 _22662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14594_ _15400_/A _23418_/Q VGND VGND VPWR VPWR _14595_/C sky130_fd_sc_hd__or2_4
X_19121_ _18987_/A _19119_/X _19120_/Y _19106_/X VGND VGND VPWR VPWR _19121_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14816__B _24057_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16333_ _16333_/A _16273_/B VGND VGND VPWR VPWR _16333_/X sky130_fd_sc_hd__or2_4
X_13545_ _12971_/A VGND VGND VPWR VPWR _13546_/A sky130_fd_sc_hd__buf_2
XFILLER_158_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19052_ _19024_/A VGND VGND VPWR VPWR _19052_/X sky130_fd_sc_hd__buf_2
X_13476_ _12894_/A _13476_/B VGND VGND VPWR VPWR _13476_/X sky130_fd_sc_hd__or2_4
X_16264_ _11904_/X _16339_/B VGND VGND VPWR VPWR _16264_/X sky130_fd_sc_hd__or2_4
XFILLER_12_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22419__B2 _22409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18003_ _17546_/Y _18138_/A _17585_/Y VGND VGND VPWR VPWR _18097_/A sky130_fd_sc_hd__o21a_4
XFILLER_173_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15215_ _14656_/A _15215_/B _15214_/X VGND VGND VPWR VPWR _15216_/C sky130_fd_sc_hd__and3_4
X_12427_ _12427_/A VGND VGND VPWR VPWR _12428_/A sky130_fd_sc_hd__buf_2
XFILLER_65_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16195_ _16195_/A VGND VGND VPWR VPWR _16219_/A sky130_fd_sc_hd__buf_2
XFILLER_142_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17846__A1 _17811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12358_ _12370_/A _23596_/Q VGND VGND VPWR VPWR _12358_/X sky130_fd_sc_hd__or2_4
XANTENNA__21642__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15146_ _14165_/A _15146_/B VGND VGND VPWR VPWR _15146_/X sky130_fd_sc_hd__or2_4
XFILLER_99_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13448__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19954_ _11638_/A _19953_/X _23086_/B _11639_/A VGND VGND VPWR VPWR _24163_/D sky130_fd_sc_hd__a2bb2o_4
X_15077_ _15096_/A _23989_/Q VGND VGND VPWR VPWR _15077_/X sky130_fd_sc_hd__or2_4
XANTENNA__12352__A _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12289_ _15442_/A VGND VGND VPWR VPWR _12858_/A sky130_fd_sc_hd__buf_2
X_18905_ _16523_/B _18897_/X _24400_/Q _18900_/X VGND VGND VPWR VPWR _18905_/X sky130_fd_sc_hd__o22a_4
X_14028_ _11659_/A VGND VGND VPWR VPWR _14075_/A sky130_fd_sc_hd__buf_2
X_19885_ _19868_/B _19903_/A _19890_/A _19884_/Y VGND VGND VPWR VPWR _19885_/X sky130_fd_sc_hd__o22a_4
XFILLER_84_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15663__A _12571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24087__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18836_ _18835_/X VGND VGND VPWR VPWR _18837_/B sky130_fd_sc_hd__buf_2
XFILLER_68_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15382__B _15382_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18767_ _19962_/B VGND VGND VPWR VPWR _19973_/A sky130_fd_sc_hd__inv_2
X_15979_ _11971_/X _15978_/X VGND VGND VPWR VPWR _15979_/X sky130_fd_sc_hd__and2_4
XANTENNA__14279__A _12454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21158__B2 _21152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13183__A _13183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17718_ _17718_/A _17418_/X VGND VGND VPWR VPWR _17720_/A sky130_fd_sc_hd__and2_4
X_18698_ _16971_/A _18698_/B VGND VGND VPWR VPWR _18698_/X sky130_fd_sc_hd__and2_4
XFILLER_36_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19771__A1 _19576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17649_ _17085_/A _17647_/B _17648_/X VGND VGND VPWR VPWR _17649_/X sky130_fd_sc_hd__o21a_4
XFILLER_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13911__A _13928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20660_ _20635_/X _20659_/X _15702_/B _20614_/X VGND VGND VPWR VPWR _20660_/X sky130_fd_sc_hd__o22a_4
XFILLER_149_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18326__A2 _18309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19319_ _24129_/Q VGND VGND VPWR VPWR _19319_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20591_ _20398_/X _20577_/X _20537_/X _20590_/Y VGND VGND VPWR VPWR _20591_/X sky130_fd_sc_hd__a211o_4
XFILLER_31_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21330__B2 _21324_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22330_ _12374_/B VGND VGND VPWR VPWR _23340_/D sky130_fd_sc_hd__buf_2
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20744__A _20744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22261_ _22151_/X _22258_/X _13841_/B _22255_/X VGND VGND VPWR VPWR _23389_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14742__A _11932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24000_ _23587_/CLK _24000_/D VGND VGND VPWR VPWR _24000_/Q sky130_fd_sc_hd__dfxtp_4
X_21212_ _21198_/A VGND VGND VPWR VPWR _21212_/X sky130_fd_sc_hd__buf_2
XFILLER_133_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22192_ _22117_/X _22187_/X _12657_/B _22191_/X VGND VGND VPWR VPWR _22192_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21633__A2 _21627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22830__A1 _14086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21143_ _20361_/X _21141_/X _24018_/Q _21138_/X VGND VGND VPWR VPWR _24018_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_7_28_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR _24398_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12262__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21074_ _20915_/X _21073_/X _14587_/B _21070_/X VGND VGND VPWR VPWR _21074_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21397__B2 _21395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20025_ _20016_/X _17703_/A _20022_/X _20024_/X VGND VGND VPWR VPWR _20026_/A sky130_fd_sc_hd__o22a_4
XANTENNA__15573__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23454__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21149__B2 _21145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13093__A _12641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11606__A _11606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11637__A1 _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21976_ _21865_/X _21974_/X _23550_/Q _21971_/X VGND VGND VPWR VPWR _21976_/X sky130_fd_sc_hd__o22a_4
XFILLER_73_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23715_ _23656_/CLK _21686_/X VGND VGND VPWR VPWR _15843_/B sky130_fd_sc_hd__dfxtp_4
X_20927_ _20726_/X _20926_/Y _19230_/A _20347_/X VGND VGND VPWR VPWR _20927_/X sky130_fd_sc_hd__o22a_4
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14917__A _14772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _11660_/A VGND VGND VPWR VPWR _15457_/A sky130_fd_sc_hd__buf_2
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22649__B2 _22648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23646_ _23646_/CLK _23646_/D VGND VGND VPWR VPWR _13776_/B sky130_fd_sc_hd__dfxtp_4
X_20858_ _24220_/Q _20773_/X _20857_/Y VGND VGND VPWR VPWR _20859_/A sky130_fd_sc_hd__o21a_4
XFILLER_148_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _17016_/C VGND VGND VPWR VPWR _11592_/A sky130_fd_sc_hd__inv_2
X_23577_ _23391_/CLK _23577_/D VGND VGND VPWR VPWR _14728_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12437__A _12847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20789_ _20267_/X VGND VGND VPWR VPWR _20789_/X sky130_fd_sc_hd__buf_2
XFILLER_70_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _13330_/A _13328_/X _13330_/C VGND VGND VPWR VPWR _13331_/C sky130_fd_sc_hd__and3_4
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22528_ _22471_/X _22522_/X _14469_/B _22526_/X VGND VGND VPWR VPWR _23227_/D sky130_fd_sc_hd__o22a_4
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _15517_/A _13229_/X _13261_/C VGND VGND VPWR VPWR _13261_/X sky130_fd_sc_hd__and3_4
XANTENNA__15748__A _11739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23030__A _23043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22459_ _22459_/A VGND VGND VPWR VPWR _22459_/X sky130_fd_sc_hd__buf_2
XANTENNA__14652__A _15625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12212_ _11880_/A VGND VGND VPWR VPWR _12698_/A sky130_fd_sc_hd__buf_2
X_15000_ _15000_/A _23669_/Q VGND VGND VPWR VPWR _15000_/X sky130_fd_sc_hd__or2_4
X_13192_ _11857_/A _11630_/A _13160_/X _12264_/X _13191_/X VGND VGND VPWR VPWR _13192_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22821__A1 _17397_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12143_ _12167_/A _23571_/Q VGND VGND VPWR VPWR _12144_/C sky130_fd_sc_hd__or2_4
X_24129_ _24134_/CLK _24129_/D HRESETn VGND VGND VPWR VPWR _24129_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17963__A _16941_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21485__A _21492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16951_ _24155_/Q VGND VGND VPWR VPWR _17667_/A sky130_fd_sc_hd__inv_2
X_12074_ _11939_/X _12074_/B _12074_/C VGND VGND VPWR VPWR _12074_/X sky130_fd_sc_hd__or3_4
XFILLER_173_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22585__B1 _15059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15902_ _13528_/A _15898_/X _15902_/C VGND VGND VPWR VPWR _15910_/B sky130_fd_sc_hd__or3_4
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19670_ _19510_/X _19670_/B VGND VGND VPWR VPWR _19670_/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12900__A _12873_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16882_ _16830_/X _16831_/B _13570_/A VGND VGND VPWR VPWR _16882_/X sky130_fd_sc_hd__o21a_4
X_18621_ _18574_/X _18620_/X _24476_/Q _18574_/X VGND VGND VPWR VPWR _18621_/X sky130_fd_sc_hd__a2bb2o_4
X_15833_ _12894_/A _15833_/B VGND VGND VPWR VPWR _15833_/X sky130_fd_sc_hd__or2_4
X_18552_ _18531_/X _18551_/X _24479_/Q _18531_/X VGND VGND VPWR VPWR _18552_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15764_ _12766_/X _15764_/B _15763_/X VGND VGND VPWR VPWR _15764_/X sky130_fd_sc_hd__and3_4
XFILLER_18_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12976_ _12976_/A _12976_/B _12975_/X VGND VGND VPWR VPWR _12977_/C sky130_fd_sc_hd__or3_4
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20829__A _20828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17503_ _17173_/Y _17503_/B VGND VGND VPWR VPWR _17504_/A sky130_fd_sc_hd__or2_4
XFILLER_166_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14715_ _14297_/A _14713_/X _14714_/X VGND VGND VPWR VPWR _14715_/X sky130_fd_sc_hd__and3_4
X_18483_ _18483_/A _18415_/A VGND VGND VPWR VPWR _18483_/X sky130_fd_sc_hd__or2_4
X_11927_ _11876_/X _11908_/X _11926_/X VGND VGND VPWR VPWR _11927_/X sky130_fd_sc_hd__or3_4
X_15695_ _13139_/A _15760_/B VGND VGND VPWR VPWR _15695_/X sky130_fd_sc_hd__or2_4
XFILLER_45_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13731__A _12576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17434_ _17434_/A _17433_/Y VGND VGND VPWR VPWR _17635_/B sky130_fd_sc_hd__or2_4
X_14646_ _14693_/A _14646_/B _14646_/C VGND VGND VPWR VPWR _14646_/X sky130_fd_sc_hd__and3_4
X_11858_ _11858_/A VGND VGND VPWR VPWR _11858_/X sky130_fd_sc_hd__buf_2
XFILLER_61_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17365_ _17365_/A _18466_/A VGND VGND VPWR VPWR _18415_/A sky130_fd_sc_hd__or2_4
XANTENNA__12347__A _12604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14577_ _13596_/A _14649_/B VGND VGND VPWR VPWR _14577_/X sky130_fd_sc_hd__or2_4
X_11789_ _11746_/X _23604_/Q VGND VGND VPWR VPWR _11790_/C sky130_fd_sc_hd__or2_4
XANTENNA__21312__B2 _21239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19104_ _11520_/A _11519_/X _19099_/Y VGND VGND VPWR VPWR _19104_/Y sky130_fd_sc_hd__a21oi_4
X_16316_ _16316_/A _16251_/B VGND VGND VPWR VPWR _16316_/X sky130_fd_sc_hd__or2_4
X_13528_ _13528_/A _13524_/X _13528_/C VGND VGND VPWR VPWR _13529_/C sky130_fd_sc_hd__or3_4
X_17296_ _17296_/A VGND VGND VPWR VPWR _22687_/A sky130_fd_sc_hd__inv_2
XFILLER_146_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19035_ _24358_/Q _11532_/B _19030_/Y VGND VGND VPWR VPWR _19035_/Y sky130_fd_sc_hd__a21oi_4
X_16247_ _16156_/A _16247_/B VGND VGND VPWR VPWR _16247_/X sky130_fd_sc_hd__or2_4
XANTENNA__15658__A _12687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13459_ _13431_/X _24069_/Q VGND VGND VPWR VPWR _13460_/C sky130_fd_sc_hd__or2_4
XANTENNA__14562__A _14280_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21615__A2 _21613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16178_ _16216_/A _16178_/B VGND VGND VPWR VPWR _16179_/C sky130_fd_sc_hd__or2_4
XFILLER_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14281__B _24028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15129_ _12433_/A _15129_/B VGND VGND VPWR VPWR _15129_/X sky130_fd_sc_hd__or2_4
XFILLER_99_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21395__A _21388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19937_ _19931_/X _24170_/Q _19932_/X _20866_/B VGND VGND VPWR VPWR _24170_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16489__A _13383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21379__B2 _21374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15393__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13906__A _14385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19868_ _19894_/C _19868_/B VGND VGND VPWR VPWR _19868_/X sky130_fd_sc_hd__and2_4
XFILLER_96_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18819_ _17161_/X _18817_/X _24448_/Q _18818_/X VGND VGND VPWR VPWR _18819_/X sky130_fd_sc_hd__o22a_4
X_19799_ _19682_/A _19740_/A VGND VGND VPWR VPWR _19809_/A sky130_fd_sc_hd__or2_4
XFILLER_55_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21830_ _21829_/X _21827_/X _23629_/Q _21822_/X VGND VGND VPWR VPWR _21830_/X sky130_fd_sc_hd__o22a_4
XFILLER_23_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22879__A1 _17574_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17717__A2_N _17360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15840__B _15840_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21761_ _21755_/Y _21760_/X _21526_/X _21760_/X VGND VGND VPWR VPWR _21761_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA_clkbuf_4_3_0_HCLK_A clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14737__A _12484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23500_ _23500_/CLK _23500_/D VGND VGND VPWR VPWR _12293_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13641__A _12186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20712_ _18472_/X _20702_/X _20514_/X _20711_/Y VGND VGND VPWR VPWR _20712_/X sky130_fd_sc_hd__a211o_4
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17113__A _12093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24480_ _24137_/CLK _18532_/X HRESETn VGND VGND VPWR VPWR _24480_/Q sky130_fd_sc_hd__dfrtp_4
X_21692_ _21577_/X _21691_/X _23711_/Q _21688_/X VGND VGND VPWR VPWR _21692_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23431_ _23303_/CLK _23431_/D VGND VGND VPWR VPWR _13241_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20643_ _20639_/X _20642_/X VGND VGND VPWR VPWR _20643_/Y sky130_fd_sc_hd__nand2_4
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21303__B2 _21300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23362_ _23908_/CLK _23362_/D VGND VGND VPWR VPWR _15458_/B sky130_fd_sc_hd__dfxtp_4
X_20574_ _22440_/A VGND VGND VPWR VPWR _20575_/A sky130_fd_sc_hd__buf_2
XANTENNA__21854__A2 _21851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22313_ _22153_/X _22308_/X _14343_/B _22312_/X VGND VGND VPWR VPWR _22313_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15568__A _14431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23293_ _23518_/CLK _23293_/D VGND VGND VPWR VPWR _13811_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14472__A _12266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24252__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20193__B _20192_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21067__B1 _24063_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22244_ _22244_/A VGND VGND VPWR VPWR _22244_/X sky130_fd_sc_hd__buf_2
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22175_ _22208_/A VGND VGND VPWR VPWR _22176_/A sky130_fd_sc_hd__inv_2
XFILLER_121_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21126_ _20915_/X _21125_/X _14563_/B _21122_/X VGND VGND VPWR VPWR _24026_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16399__A _15998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22567__B1 _15796_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13816__A _14319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21057_ _20613_/X _21052_/X _24070_/Q _21056_/X VGND VGND VPWR VPWR _24070_/D sky130_fd_sc_hd__o22a_4
XFILLER_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20008_ _20008_/A VGND VGND VPWR VPWR _20008_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21790__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12830_ _13370_/A _12747_/B VGND VGND VPWR VPWR _12830_/X sky130_fd_sc_hd__or2_4
XFILLER_43_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19735__A1 _20512_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23025__A _23043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12761_ _13055_/A VGND VGND VPWR VPWR _12762_/A sky130_fd_sc_hd__buf_2
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21959_ _21836_/X _21953_/X _12804_/B _21957_/X VGND VGND VPWR VPWR _21959_/X sky130_fd_sc_hd__o22a_4
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14647__A _15595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14500_ _14378_/A _14500_/B VGND VGND VPWR VPWR _14500_/X sky130_fd_sc_hd__or2_4
X_11712_ _13248_/A VGND VGND VPWR VPWR _11712_/X sky130_fd_sc_hd__buf_2
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12571_/A _12692_/B _12691_/X VGND VGND VPWR VPWR _12692_/X sky130_fd_sc_hd__or3_4
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _13053_/A _23330_/Q VGND VGND VPWR VPWR _15482_/B sky130_fd_sc_hd__or2_4
XFILLER_43_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14431_/A _14431_/B _14431_/C VGND VGND VPWR VPWR _14431_/X sky130_fd_sc_hd__and3_4
X_11643_ _11643_/A VGND VGND VPWR VPWR _11643_/Y sky130_fd_sc_hd__inv_2
X_23629_ _24077_/CLK _21830_/X VGND VGND VPWR VPWR _23629_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _17112_/X _17123_/X _17136_/X _17137_/X _17149_/X VGND VGND VPWR VPWR _17150_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14362_ _14369_/A _14362_/B VGND VGND VPWR VPWR _14362_/X sky130_fd_sc_hd__or2_4
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11574_ _24456_/Q IRQ[19] _20178_/A VGND VGND VPWR VPWR _11574_/X sky130_fd_sc_hd__a21o_4
XFILLER_126_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20502__C1 _20501_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17677__B _17464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16101_ _16101_/A VGND VGND VPWR VPWR _16109_/A sky130_fd_sc_hd__buf_2
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _13313_/A _24070_/Q VGND VGND VPWR VPWR _13314_/C sky130_fd_sc_hd__or2_4
XFILLER_156_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17081_ _17017_/B _18772_/A _17090_/B VGND VGND VPWR VPWR _17082_/B sky130_fd_sc_hd__or3_4
X_14293_ _11930_/A VGND VGND VPWR VPWR _15022_/A sky130_fd_sc_hd__buf_2
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16032_ _16057_/A _24046_/Q VGND VGND VPWR VPWR _16032_/X sky130_fd_sc_hd__or2_4
X_13244_ _12354_/A _13236_/X _13243_/X VGND VGND VPWR VPWR _13260_/B sky130_fd_sc_hd__and3_4
XFILLER_171_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14_0_HCLK_A clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13175_ _12851_/A VGND VGND VPWR VPWR _13324_/A sky130_fd_sc_hd__buf_2
XFILLER_108_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22270__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12126_ _11762_/X _12124_/X _12126_/C VGND VGND VPWR VPWR _12126_/X sky130_fd_sc_hd__and3_4
XFILLER_112_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17983_ _17819_/X _17827_/X _17230_/X _17835_/X VGND VGND VPWR VPWR _17983_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_11_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR _23475_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_123_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19722_ HRDATA[22] VGND VGND VPWR VPWR _20866_/B sky130_fd_sc_hd__buf_2
Xclkbuf_7_74_0_HCLK clkbuf_7_74_0_HCLK/A VGND VGND VPWR VPWR _23456_/CLK sky130_fd_sc_hd__clkbuf_1
X_16934_ _16933_/Y VGND VGND VPWR VPWR _16935_/A sky130_fd_sc_hd__buf_2
XFILLER_77_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12057_ _16744_/A VGND VGND VPWR VPWR _12058_/A sky130_fd_sc_hd__buf_2
XANTENNA__22022__A2 _22017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20569__C1 _20568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21230__B1 _15156_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21943__A _21950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19653_ _19857_/B VGND VGND VPWR VPWR _19778_/B sky130_fd_sc_hd__inv_2
XFILLER_78_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16865_ _15386_/X _14848_/Y _16864_/Y _14847_/X VGND VGND VPWR VPWR _16865_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18604_ _17980_/X _17621_/B _18599_/X _18602_/X _18603_/X VGND VGND VPWR VPWR _18604_/X
+ sky130_fd_sc_hd__a32o_4
X_15816_ _12858_/A _15812_/X _15816_/C VGND VGND VPWR VPWR _15816_/X sky130_fd_sc_hd__or3_4
XFILLER_168_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19584_ _19705_/A _19557_/Y VGND VGND VPWR VPWR _19601_/B sky130_fd_sc_hd__and2_4
X_16796_ _16757_/X _23857_/Q VGND VGND VPWR VPWR _16797_/C sky130_fd_sc_hd__or2_4
XFILLER_52_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24125__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18535_ _24141_/Q _18534_/Y _16979_/X VGND VGND VPWR VPWR _22961_/B sky130_fd_sc_hd__o21a_4
X_15747_ _15778_/A _15675_/B VGND VGND VPWR VPWR _15747_/X sky130_fd_sc_hd__or2_4
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12959_ _12971_/A _23433_/Q VGND VGND VPWR VPWR _12960_/C sky130_fd_sc_hd__or2_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14557__A _14270_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13461__A _13475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21533__B2 _21525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18466_ _18466_/A _18415_/C VGND VGND VPWR VPWR _18466_/X sky130_fd_sc_hd__or2_4
X_15678_ _12228_/A _23940_/Q VGND VGND VPWR VPWR _15680_/B sky130_fd_sc_hd__or2_4
X_17417_ _11592_/X _17358_/B _17416_/X _17342_/Y VGND VGND VPWR VPWR _17418_/B sky130_fd_sc_hd__a211o_4
XANTENNA__17868__A _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14629_ _14660_/A _14621_/X _14629_/C VGND VGND VPWR VPWR _14629_/X sky130_fd_sc_hd__or3_4
X_18397_ _18180_/X _17773_/X _18180_/X _17773_/X VGND VGND VPWR VPWR _18397_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12077__A _11984_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24275__CLK _24471_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17348_ _15252_/X _17333_/B _18709_/A _17347_/X VGND VGND VPWR VPWR _17348_/X sky130_fd_sc_hd__o22a_4
XFILLER_174_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14292__A _14292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17279_ _17275_/X VGND VGND VPWR VPWR _17280_/B sky130_fd_sc_hd__buf_2
XANTENNA__12805__A _13349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19018_ _19018_/A VGND VGND VPWR VPWR _19018_/Y sky130_fd_sc_hd__inv_2
X_20290_ _18953_/B _20344_/A VGND VGND VPWR VPWR _20290_/X sky130_fd_sc_hd__and2_4
XANTENNA__22261__A2 _22258_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22014__A _22007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22013__A2 _22010_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23980_ _24012_/CLK _21201_/X VGND VGND VPWR VPWR _23980_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16012__A _15934_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22949__A _22949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22931_ _22931_/A _22931_/B VGND VGND VPWR VPWR _22931_/X sky130_fd_sc_hd__and2_4
XFILLER_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21772__B2 _21767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15851__A _15851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22862_ _22861_/X VGND VGND VPWR VPWR HWDATA[19] sky130_fd_sc_hd__inv_2
XANTENNA__15451__A1 _11969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21813_ _21528_/A VGND VGND VPWR VPWR _21813_/X sky130_fd_sc_hd__buf_2
X_22793_ _22793_/A _22791_/X _22792_/Y VGND VGND VPWR VPWR _22793_/X sky130_fd_sc_hd__and3_4
XANTENNA__13371__A _13379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21744_ _21582_/X _21741_/X _23677_/Q _21738_/X VGND VGND VPWR VPWR _23677_/D sky130_fd_sc_hd__o22a_4
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21675_ _21548_/X _21670_/X _12664_/B _21674_/X VGND VGND VPWR VPWR _23723_/D sky130_fd_sc_hd__o22a_4
XFILLER_12_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24463_ _23379_/CLK _24463_/D HRESETn VGND VGND VPWR VPWR _24463_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16682__A _16682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20626_ _18394_/X _20446_/X _20538_/X _20625_/Y VGND VGND VPWR VPWR _20626_/X sky130_fd_sc_hd__a211o_4
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23414_ _23095_/CLK _23414_/D VGND VGND VPWR VPWR _14891_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_137_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24394_ _24422_/CLK _24394_/D HRESETn VGND VGND VPWR VPWR _24394_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14914__B _14850_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23642__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15298__A _12453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23345_ _23409_/CLK _23345_/D VGND VGND VPWR VPWR _16782_/B sky130_fd_sc_hd__dfxtp_4
X_20557_ _24233_/Q _20534_/X _20556_/X VGND VGND VPWR VPWR _20558_/A sky130_fd_sc_hd__o21a_4
XFILLER_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12715__A _12266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23276_ _23500_/CLK _22431_/X VGND VGND VPWR VPWR _12193_/B sky130_fd_sc_hd__dfxtp_4
X_20488_ _20444_/X _20866_/B _20308_/X VGND VGND VPWR VPWR _20488_/X sky130_fd_sc_hd__a21o_4
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18456__A1 _18022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22227_ _22226_/X VGND VGND VPWR VPWR _22227_/X sky130_fd_sc_hd__buf_2
XANTENNA__22252__A2 _22251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22158_ _22158_/A VGND VGND VPWR VPWR _22158_/X sky130_fd_sc_hd__buf_2
XANTENNA__13546__A _13546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21109_ _20613_/X _21104_/X _13286_/B _21108_/X VGND VGND VPWR VPWR _21109_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22004__A2 _22003_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19405__B1 _19402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14980_ _14614_/A _14972_/X _14979_/X VGND VGND VPWR VPWR _14980_/X sky130_fd_sc_hd__and3_4
X_22089_ _21603_/A VGND VGND VPWR VPWR _22090_/A sky130_fd_sc_hd__buf_2
XANTENNA__12450__A _12194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21763__A _21770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24148__CLK _24271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13931_ _14385_/A _13929_/X _13930_/X VGND VGND VPWR VPWR _13931_/X sky130_fd_sc_hd__and3_4
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15761__A _13099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16650_ _16678_/A _16648_/X _16649_/X VGND VGND VPWR VPWR _16651_/C sky130_fd_sc_hd__and3_4
X_13862_ _11969_/A _13837_/X _13844_/X _13851_/X _13861_/X VGND VGND VPWR VPWR _13862_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24121__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15601_ _15610_/A _15601_/B VGND VGND VPWR VPWR _15603_/B sky130_fd_sc_hd__or2_4
X_12813_ _12801_/A _24074_/Q VGND VGND VPWR VPWR _12814_/C sky130_fd_sc_hd__or2_4
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16581_ _16558_/A _16664_/B VGND VGND VPWR VPWR _16581_/X sky130_fd_sc_hd__or2_4
XANTENNA__14377__A _14377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13793_ _15007_/A VGND VGND VPWR VPWR _13952_/A sky130_fd_sc_hd__buf_2
XANTENNA__21515__B2 _21510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23172__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24298__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18320_ _18320_/A _18319_/Y VGND VGND VPWR VPWR _18320_/X sky130_fd_sc_hd__and2_4
X_15532_ _11886_/A _24033_/Q VGND VGND VPWR VPWR _15532_/X sky130_fd_sc_hd__or2_4
X_12744_ _12311_/A _12825_/B VGND VGND VPWR VPWR _12745_/C sky130_fd_sc_hd__or2_4
XANTENNA__22594__A _22608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18251_ _18251_/A VGND VGND VPWR VPWR _18251_/Y sky130_fd_sc_hd__inv_2
X_15463_ _15487_/A _23778_/Q VGND VGND VPWR VPWR _15464_/C sky130_fd_sc_hd__or2_4
X_12675_ _12977_/A _12667_/X _12675_/C VGND VGND VPWR VPWR _12676_/C sky130_fd_sc_hd__and3_4
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16592__A _16592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _17202_/A VGND VGND VPWR VPWR _17202_/Y sky130_fd_sc_hd__inv_2
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _14334_/X _14413_/Y VGND VGND VPWR VPWR _15389_/A sky130_fd_sc_hd__or2_4
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21818__A2 _21815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18182_ _17775_/C _18181_/X _17700_/X VGND VGND VPWR VPWR _18182_/X sky130_fd_sc_hd__o21a_4
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _11625_/X VGND VGND VPWR VPWR _11627_/A sky130_fd_sc_hd__buf_2
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15394_ _15394_/A _15392_/X _15393_/X VGND VGND VPWR VPWR _15398_/B sky130_fd_sc_hd__and3_4
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _17146_/A VGND VGND VPWR VPWR _17133_/X sky130_fd_sc_hd__buf_2
X_14345_ _14367_/A _14345_/B VGND VGND VPWR VPWR _14345_/X sky130_fd_sc_hd__or2_4
XFILLER_129_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19892__B1 _20216_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ _24458_/Q IRQ[21] _20180_/A VGND VGND VPWR VPWR _11557_/X sky130_fd_sc_hd__a21o_4
XFILLER_144_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17064_ _17090_/A _17059_/X _17062_/X _20216_/D _17251_/B VGND VGND VPWR VPWR _17100_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21938__A _21028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14276_ _15398_/A _14271_/X _14276_/C VGND VGND VPWR VPWR _14276_/X sky130_fd_sc_hd__or3_4
XFILLER_170_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16015_ _11858_/X _11631_/X _15980_/X _11608_/A _16014_/X VGND VGND VPWR VPWR _16015_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15936__A _11882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13227_ _13251_/A _13227_/B _13227_/C VGND VGND VPWR VPWR _13228_/C sky130_fd_sc_hd__or3_4
XANTENNA__22243__A2 _22237_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20561__B _20561_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13158_ _12858_/A _13154_/X _13158_/C VGND VGND VPWR VPWR _13158_/X sky130_fd_sc_hd__or3_4
XFILLER_170_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13456__A _13427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12109_ _11868_/X _12109_/B VGND VGND VPWR VPWR _12109_/X sky130_fd_sc_hd__and2_4
X_13089_ _13089_/A _13006_/B VGND VGND VPWR VPWR _13089_/X sky130_fd_sc_hd__or2_4
XANTENNA__12360__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17966_ _17908_/B _17964_/X _17908_/A _17965_/X VGND VGND VPWR VPWR _17966_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21203__B1 _23979_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19705_ _19705_/A _19705_/B VGND VGND VPWR VPWR _19705_/X sky130_fd_sc_hd__or2_4
XANTENNA__24209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16917_ _16918_/A _16921_/A VGND VGND VPWR VPWR _17096_/A sky130_fd_sc_hd__or2_4
X_17897_ _16935_/X _17893_/X _17653_/X _17896_/X VGND VGND VPWR VPWR _17897_/X sky130_fd_sc_hd__o22a_4
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17958__B1 _17014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21754__B2 _21717_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15671__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19636_ HRDATA[26] VGND VGND VPWR VPWR _20776_/A sky130_fd_sc_hd__buf_2
X_16848_ _15921_/Y _16848_/B VGND VGND VPWR VPWR _16848_/X sky130_fd_sc_hd__and2_4
XFILLER_20_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_4_0_HCLK clkbuf_6_2_0_HCLK/X VGND VGND VPWR VPWR _24342_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19567_ _19518_/A VGND VGND VPWR VPWR _19573_/A sky130_fd_sc_hd__buf_2
X_16779_ _16755_/X _23697_/Q VGND VGND VPWR VPWR _16781_/B sky130_fd_sc_hd__or2_4
XANTENNA__20309__A2 _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14287__A _15400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11704__A _16047_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18518_ _18518_/A VGND VGND VPWR VPWR _18518_/X sky130_fd_sc_hd__buf_2
X_19498_ _19445_/A _19497_/X HRDATA[14] _19461_/A VGND VGND VPWR VPWR _19499_/A sky130_fd_sc_hd__o22a_4
XANTENNA__23665__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18449_ _18330_/X _18436_/Y _18373_/X _18448_/X VGND VGND VPWR VPWR _18449_/X sky130_fd_sc_hd__o22a_4
X_21460_ _21299_/X _21455_/X _14388_/B _21459_/X VGND VGND VPWR VPWR _23836_/D sky130_fd_sc_hd__o22a_4
XFILLER_147_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20411_ _20398_/X _20399_/X _20714_/A _20410_/Y VGND VGND VPWR VPWR _20411_/X sky130_fd_sc_hd__a211o_4
X_21391_ _21391_/A VGND VGND VPWR VPWR _21391_/X sky130_fd_sc_hd__buf_2
XANTENNA__12535__A _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16007__A _13441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23130_ _23641_/CLK _22680_/X VGND VGND VPWR VPWR _14590_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21690__B1 _23712_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20342_ _20260_/A VGND VGND VPWR VPWR _20342_/X sky130_fd_sc_hd__buf_2
XFILLER_162_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15846__A _12911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23061_ _23051_/A _23061_/B _23061_/C VGND VGND VPWR VPWR _23061_/X sky130_fd_sc_hd__and3_4
XANTENNA__19635__B1 _17274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20273_ _20273_/A VGND VGND VPWR VPWR _20273_/X sky130_fd_sc_hd__buf_2
XANTENNA__14750__A _12190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22012_ _21841_/X _22010_/X _23528_/Q _22007_/X VGND VGND VPWR VPWR _23528_/D sky130_fd_sc_hd__o22a_4
XFILLER_161_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12270__A _12690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22679__A _22672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23963_ _23592_/CLK _21225_/X VGND VGND VPWR VPWR _23963_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22914_ _19924_/A _16971_/A _23080_/A VGND VGND VPWR VPWR _22914_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18610__A1 _17980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20953__C1 _20952_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23894_ _23862_/CLK _23894_/D VGND VGND VPWR VPWR _14880_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22845_ _22845_/A _22845_/B VGND VGND VPWR VPWR HWDATA[15] sky130_fd_sc_hd__nor2_4
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11614__A _11965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22776_ _22790_/C VGND VGND VPWR VPWR _22793_/A sky130_fd_sc_hd__buf_2
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22170__B2 _22106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21727_ _21727_/A VGND VGND VPWR VPWR _21727_/X sky130_fd_sc_hd__buf_2
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21658_ _21658_/A VGND VGND VPWR VPWR _21674_/A sky130_fd_sc_hd__inv_2
X_12460_ _12288_/A VGND VGND VPWR VPWR _12461_/A sky130_fd_sc_hd__buf_2
XFILLER_32_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24446_ _23476_/CLK _18821_/X HRESETn VGND VGND VPWR VPWR _24446_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12391_ _11701_/A _12389_/X _12391_/C VGND VGND VPWR VPWR _12391_/X sky130_fd_sc_hd__and3_4
X_20609_ _20466_/X _20599_/Y _20607_/X _20608_/Y _20481_/X VGND VGND VPWR VPWR _20610_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18677__A1 _17805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12445__A _12445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24377_ _24382_/CLK _24377_/D HRESETn VGND VGND VPWR VPWR _24377_/Q sky130_fd_sc_hd__dfstp_4
X_21589_ _21304_/A VGND VGND VPWR VPWR _21589_/X sky130_fd_sc_hd__buf_2
XFILLER_137_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14130_ _14108_/A _23167_/Q VGND VGND VPWR VPWR _14130_/X sky130_fd_sc_hd__or2_4
XFILLER_158_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21758__A _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23328_ _23101_/CLK _23328_/D VGND VGND VPWR VPWR _22342_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14061_ _13696_/A _14059_/X _14061_/C VGND VGND VPWR VPWR _14065_/B sky130_fd_sc_hd__and3_4
X_23259_ _24096_/CLK _22472_/X VGND VGND VPWR VPWR _14484_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13012_ _12498_/A _13012_/B VGND VGND VPWR VPWR _13012_/X sky130_fd_sc_hd__or2_4
XFILLER_134_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13276__A _13276_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21984__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17820_ _17819_/X VGND VGND VPWR VPWR _17820_/X sky130_fd_sc_hd__buf_2
XANTENNA__17971__A _17801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23538__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22589__A _22622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19929__B2 _20364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24302__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17751_ _17751_/A _17751_/B VGND VGND VPWR VPWR _17751_/X sky130_fd_sc_hd__or2_4
XFILLER_88_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14963_ _14786_/A _14961_/X _14962_/X VGND VGND VPWR VPWR _14963_/X sky130_fd_sc_hd__and3_4
XFILLER_59_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21736__B2 _21731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16702_ _16702_/A _16702_/B _16701_/X VGND VGND VPWR VPWR _16702_/X sky130_fd_sc_hd__and3_4
X_13914_ _14377_/A _23965_/Q VGND VGND VPWR VPWR _13915_/C sky130_fd_sc_hd__or2_4
X_17682_ _24151_/Q _17455_/X _17681_/X VGND VGND VPWR VPWR _17683_/B sky130_fd_sc_hd__o21ai_4
X_14894_ _14108_/A _23478_/Q VGND VGND VPWR VPWR _14894_/X sky130_fd_sc_hd__or2_4
XFILLER_48_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19421_ _19406_/X VGND VGND VPWR VPWR _19421_/X sky130_fd_sc_hd__buf_2
XANTENNA__14819__B _14743_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16633_ _16662_/A _23602_/Q VGND VGND VPWR VPWR _16633_/X sky130_fd_sc_hd__or2_4
XFILLER_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13845_ _13675_/A _13845_/B VGND VGND VPWR VPWR _13847_/B sky130_fd_sc_hd__or2_4
XFILLER_63_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19352_ _19350_/X _18304_/X _19350_/X _20570_/A VGND VGND VPWR VPWR _19352_/X sky130_fd_sc_hd__a2bb2o_4
X_16564_ _12001_/A _16562_/X _16564_/C VGND VGND VPWR VPWR _16568_/B sky130_fd_sc_hd__and3_4
X_13776_ _12610_/A _13776_/B VGND VGND VPWR VPWR _13776_/X sky130_fd_sc_hd__or2_4
XFILLER_62_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18303_ _17697_/B _18302_/X _17688_/X VGND VGND VPWR VPWR _18303_/X sky130_fd_sc_hd__o21a_4
X_15515_ _11682_/A _15507_/X _15514_/X VGND VGND VPWR VPWR _15515_/X sky130_fd_sc_hd__and3_4
X_12727_ _12727_/A _12816_/B VGND VGND VPWR VPWR _12727_/X sky130_fd_sc_hd__or2_4
X_19283_ _19245_/B VGND VGND VPWR VPWR _19283_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16495_ _16507_/A _16495_/B _16495_/C VGND VGND VPWR VPWR _16495_/X sky130_fd_sc_hd__and3_4
XANTENNA__18307__A _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18234_ _18234_/A VGND VGND VPWR VPWR _18234_/Y sky130_fd_sc_hd__inv_2
X_15446_ _15446_/A _23714_/Q VGND VGND VPWR VPWR _15446_/X sky130_fd_sc_hd__or2_4
X_12658_ _12670_/A _12655_/X _12658_/C VGND VGND VPWR VPWR _12659_/C sky130_fd_sc_hd__and3_4
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18165_ _17461_/X _18165_/B _18164_/X VGND VGND VPWR VPWR _18166_/B sky130_fd_sc_hd__or3_4
X_11609_ _11608_/X VGND VGND VPWR VPWR _11609_/X sky130_fd_sc_hd__buf_2
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19865__B1 _21184_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15377_ _15377_/A _15369_/X _15377_/C VGND VGND VPWR VPWR _15378_/C sky130_fd_sc_hd__and3_4
X_12589_ _12925_/A VGND VGND VPWR VPWR _12970_/A sky130_fd_sc_hd__buf_2
XANTENNA__12355__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17116_ _17198_/A VGND VGND VPWR VPWR _17116_/X sky130_fd_sc_hd__buf_2
XFILLER_117_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14328_ _13666_/A _14399_/B VGND VGND VPWR VPWR _14330_/B sky130_fd_sc_hd__or2_4
X_18096_ _18116_/B _17640_/X VGND VGND VPWR VPWR _18096_/X sky130_fd_sc_hd__or2_4
XANTENNA__20572__A _20438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24313__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15666__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17047_ _17047_/A VGND VGND VPWR VPWR _17047_/X sky130_fd_sc_hd__buf_2
XFILLER_132_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19617__B1 HRDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14259_ _11812_/A _14259_/B _14258_/X VGND VGND VPWR VPWR _14259_/X sky130_fd_sc_hd__or3_4
XANTENNA__22216__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14570__A _15395_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24388__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21975__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13186__A _11887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18998_ _18987_/X _18996_/X _18997_/Y _18990_/X VGND VGND VPWR VPWR _18998_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_6_44_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_89_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17949_ _17877_/X _17948_/X _17880_/X VGND VGND VPWR VPWR _17949_/X sky130_fd_sc_hd__o21a_4
XFILLER_39_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13914__A _14377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20960_ _20894_/X _20959_/X _24088_/Q _20861_/X VGND VGND VPWR VPWR _24088_/D sky130_fd_sc_hd__o22a_4
XFILLER_26_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19619_ _19619_/A VGND VGND VPWR VPWR _19898_/B sky130_fd_sc_hd__inv_2
XFILLER_4_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20891_ _22471_/A VGND VGND VPWR VPWR _20892_/A sky130_fd_sc_hd__buf_2
XPHY_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22630_ _22473_/X _22629_/X _14649_/B _22626_/X VGND VGND VPWR VPWR _23162_/D sky130_fd_sc_hd__o22a_4
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22152__B2 _22142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22561_ _22442_/X _22558_/X _13204_/B _22555_/X VGND VGND VPWR VPWR _23207_/D sky130_fd_sc_hd__o22a_4
XFILLER_16_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14745__A _12469_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18217__A _18148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24300_ _24302_/CLK _24300_/D HRESETn VGND VGND VPWR VPWR _24300_/Q sky130_fd_sc_hd__dfrtp_4
X_21512_ _21302_/X _21506_/X _14474_/B _21510_/X VGND VGND VPWR VPWR _23803_/D sky130_fd_sc_hd__o22a_4
XFILLER_166_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22492_ _22486_/Y _22491_/X _22410_/X _22491_/X VGND VGND VPWR VPWR _22492_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22962__A _18548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21443_ _21271_/X _21441_/X _23848_/Q _21438_/X VGND VGND VPWR VPWR _23848_/D sky130_fd_sc_hd__o22a_4
X_24231_ _24127_/CLK _19410_/X HRESETn VGND VGND VPWR VPWR _24231_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12265__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24162_ _24472_/CLK _19982_/Y HRESETn VGND VGND VPWR VPWR _19328_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21578__A _21523_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21374_ _21381_/A VGND VGND VPWR VPWR _21374_/X sky130_fd_sc_hd__buf_2
XFILLER_162_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23113_ _24073_/CLK _23113_/D VGND VGND VPWR VPWR _12963_/B sky130_fd_sc_hd__dfxtp_4
X_20325_ _20267_/X VGND VGND VPWR VPWR _20325_/X sky130_fd_sc_hd__buf_2
XANTENNA__15576__A _12434_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24093_ _23880_/CLK _20842_/X VGND VGND VPWR VPWR _24093_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19608__B1 _17398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22207__A2 _22201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14480__A _14480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_126_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR _23337_/CLK sky130_fd_sc_hd__clkbuf_1
X_23044_ _18140_/X _23055_/B VGND VGND VPWR VPWR _23045_/C sky130_fd_sc_hd__or2_4
X_20256_ _17091_/A _16918_/X _16922_/C _11598_/X VGND VGND VPWR VPWR _20257_/A sky130_fd_sc_hd__or4_4
XANTENNA__21966__A1 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21966__B2 _21964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17791__A _18150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18831__A1 _15118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11609__A _11608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20187_ _24464_/Q IRQ[27] _20186_/X VGND VGND VPWR VPWR _20188_/B sky130_fd_sc_hd__a21boi_4
XFILLER_118_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21718__B2 _21717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13824__A _15415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23946_ _23531_/CLK _23946_/D VGND VGND VPWR VPWR _12789_/B sky130_fd_sc_hd__dfxtp_4
X_11960_ _11960_/A VGND VGND VPWR VPWR _12105_/A sky130_fd_sc_hd__buf_2
XANTENNA__21194__A2 _21191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22391__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23877_ _23241_/CLK _21397_/X VGND VGND VPWR VPWR _13480_/B sky130_fd_sc_hd__dfxtp_4
X_11891_ _11890_/X VGND VGND VPWR VPWR _11891_/X sky130_fd_sc_hd__buf_2
X_13630_ _13630_/A VGND VGND VPWR VPWR _14329_/A sky130_fd_sc_hd__buf_2
X_22828_ _22814_/X _22827_/X VGND VGND VPWR VPWR HWDATA[10] sky130_fd_sc_hd__nor2_4
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18347__B1 _18168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22143__B2 _22142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13561_ _13554_/A _23653_/Q VGND VGND VPWR VPWR _13562_/C sky130_fd_sc_hd__or2_4
XFILLER_164_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22759_ _22758_/Y _22773_/B _22758_/Y _22773_/B VGND VGND VPWR VPWR _22759_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15300_ _14295_/A _15300_/B VGND VGND VPWR VPWR _15300_/X sky130_fd_sc_hd__or2_4
XFILLER_73_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12512_ _12512_/A VGND VGND VPWR VPWR _12513_/A sky130_fd_sc_hd__buf_2
X_16280_ _16287_/A _16280_/B VGND VGND VPWR VPWR _16280_/X sky130_fd_sc_hd__or2_4
XFILLER_12_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13492_ _12972_/A VGND VGND VPWR VPWR _13547_/A sky130_fd_sc_hd__buf_2
XFILLER_100_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15231_ _14191_/A _15229_/X _15230_/X VGND VGND VPWR VPWR _15232_/C sky130_fd_sc_hd__and3_4
X_12443_ _15018_/A VGND VGND VPWR VPWR _12444_/A sky130_fd_sc_hd__buf_2
X_24429_ _24428_/CLK _24429_/D HRESETn VGND VGND VPWR VPWR _20448_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22446__A2 _22438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19847__B1 _21134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20457__A1 _18140_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15162_ _15267_/A _15162_/B VGND VGND VPWR VPWR _15164_/B sky130_fd_sc_hd__or2_4
XANTENNA__21654__B1 _23733_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12374_ _12373_/X _12374_/B VGND VGND VPWR VPWR _12377_/B sky130_fd_sc_hd__or2_4
XANTENNA__20392__A _20358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17322__A1 _17319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14113_ _11910_/A VGND VGND VPWR VPWR _14114_/A sky130_fd_sc_hd__buf_2
XFILLER_114_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14390__A _14390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19970_ _17645_/X VGND VGND VPWR VPWR _19970_/Y sky130_fd_sc_hd__inv_2
X_15093_ _15086_/A _23829_/Q VGND VGND VPWR VPWR _15093_/X sky130_fd_sc_hd__or2_4
XANTENNA__23360__CLK _23456_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24486__CLK _24271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18921_ _18928_/A VGND VGND VPWR VPWR _18921_/X sky130_fd_sc_hd__buf_2
X_14044_ _13696_/A _14042_/X _14043_/X VGND VGND VPWR VPWR _14044_/X sky130_fd_sc_hd__and3_4
XFILLER_134_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18852_ _17139_/X _18849_/X _24430_/Q _18850_/X VGND VGND VPWR VPWR _24430_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18822__A1 _13945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17803_ _17793_/X _17795_/X _17799_/X _17803_/D VGND VGND VPWR VPWR _17804_/A sky130_fd_sc_hd__or4_4
XFILLER_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18783_ _12027_/X _18888_/B _11633_/X _18834_/C VGND VGND VPWR VPWR _18784_/B sky130_fd_sc_hd__or4_4
X_15995_ _15967_/A _16076_/B VGND VGND VPWR VPWR _15995_/X sky130_fd_sc_hd__or2_4
XFILLER_121_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17734_ _17734_/A _17280_/X VGND VGND VPWR VPWR _17734_/X sky130_fd_sc_hd__or2_4
X_14946_ _14970_/A _14946_/B VGND VGND VPWR VPWR _14947_/C sky130_fd_sc_hd__or2_4
XFILLER_76_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16110__A _16110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22382__B2 _22380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17665_ _17663_/X _17664_/Y VGND VGND VPWR VPWR _17671_/A sky130_fd_sc_hd__or2_4
X_14877_ _11929_/A _14873_/X _14876_/X VGND VGND VPWR VPWR _14878_/B sky130_fd_sc_hd__or3_4
XFILLER_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16616_ _11836_/A VGND VGND VPWR VPWR _16662_/A sky130_fd_sc_hd__buf_2
X_19404_ _19404_/A VGND VGND VPWR VPWR _19404_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19421__A _19406_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13828_ _11932_/A _13824_/X _13827_/X VGND VGND VPWR VPWR _13828_/X sky130_fd_sc_hd__or3_4
X_17596_ _17562_/A _17595_/Y _17554_/B _18039_/B VGND VGND VPWR VPWR _17642_/B sky130_fd_sc_hd__a211o_4
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19335_ _20200_/A VGND VGND VPWR VPWR _19335_/X sky130_fd_sc_hd__buf_2
X_16547_ _16534_/X _24050_/Q VGND VGND VPWR VPWR _16549_/B sky130_fd_sc_hd__or2_4
X_13759_ _14543_/A _13757_/X _13759_/C VGND VGND VPWR VPWR _13759_/X sky130_fd_sc_hd__and3_4
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22685__A2 _22658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14565__A _15394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19266_ _19253_/A _19253_/B _19265_/Y VGND VGND VPWR VPWR _24304_/D sky130_fd_sc_hd__o21a_4
X_16478_ _16370_/X _16474_/X _16478_/C VGND VGND VPWR VPWR _16478_/X sky130_fd_sc_hd__or3_4
XFILLER_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18217_ _18148_/A _18148_/B _18217_/C VGND VGND VPWR VPWR _18217_/X sky130_fd_sc_hd__and3_4
XFILLER_31_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15429_ _15406_/A _15493_/B VGND VGND VPWR VPWR _15431_/B sky130_fd_sc_hd__or2_4
X_19197_ _19143_/X VGND VGND VPWR VPWR _19197_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19838__B1 _16922_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21398__A _21391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18148_ _18148_/A _18148_/B _18148_/C VGND VGND VPWR VPWR _18148_/X sky130_fd_sc_hd__and3_4
XFILLER_160_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15396__A _15400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18079_ _18283_/A _18079_/B _18079_/C _18079_/D VGND VGND VPWR VPWR _18080_/A sky130_fd_sc_hd__or4_4
XANTENNA__13909__A _13720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12813__A _12801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20110_ _11558_/X VGND VGND VPWR VPWR _20110_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21090_ _21104_/A VGND VGND VPWR VPWR _21090_/X sky130_fd_sc_hd__buf_2
XFILLER_160_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21948__B2 _21943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20041_ _24487_/Q VGND VGND VPWR VPWR _20041_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18813__A1 _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23800_ _23098_/CLK _23800_/D VGND VGND VPWR VPWR _15305_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13644__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24209__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16020__A _16056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21992_ _22007_/A VGND VGND VPWR VPWR _22000_/A sky130_fd_sc_hd__buf_2
XFILLER_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14459__B _14523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23731_ _23119_/CLK _21664_/X VGND VGND VPWR VPWR _23731_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20943_ _20943_/A _20942_/X VGND VGND VPWR VPWR _20943_/X sky130_fd_sc_hd__and2_4
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _23662_/CLK _23662_/D VGND VGND VPWR VPWR _23662_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20874_ _19721_/Y _20873_/X _20866_/B _20843_/B VGND VGND VPWR VPWR _20874_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22613_ _22444_/X _22608_/X _23174_/Q _22612_/X VGND VGND VPWR VPWR _23174_/D sky130_fd_sc_hd__o22a_4
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23593_ _24073_/CLK _21910_/X VGND VGND VPWR VPWR _23593_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14475__A _12470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20196__B _20195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22544_ _22558_/A VGND VGND VPWR VPWR _22544_/X sky130_fd_sc_hd__buf_2
XFILLER_10_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11611__B _11611_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19829__B1 _18780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22475_ _22473_/X _22474_/X _14618_/B _22469_/X VGND VGND VPWR VPWR _23258_/D sky130_fd_sc_hd__o22a_4
XFILLER_136_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23383__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24214_ _24248_/CLK _19434_/X HRESETn VGND VGND VPWR VPWR _24214_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21426_ _21455_/A VGND VGND VPWR VPWR _21441_/A sky130_fd_sc_hd__buf_2
XFILLER_108_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21100__A2 _21097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21101__A _21101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13819__A _12198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24145_ _24134_/CLK _20063_/Y HRESETn VGND VGND VPWR VPWR _24145_/Q sky130_fd_sc_hd__dfrtp_4
X_21357_ _21295_/X _21355_/X _13750_/B _21352_/X VGND VGND VPWR VPWR _21357_/X sky130_fd_sc_hd__o22a_4
XFILLER_2_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12723__A _13277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20308_ _20308_/A VGND VGND VPWR VPWR _20308_/X sky130_fd_sc_hd__buf_2
X_12090_ _12059_/X _12159_/B VGND VGND VPWR VPWR _12091_/C sky130_fd_sc_hd__or2_4
X_24076_ _24074_/CLK _21048_/X VGND VGND VPWR VPWR _24076_/Q sky130_fd_sc_hd__dfxtp_4
X_21288_ _21264_/A VGND VGND VPWR VPWR _21288_/X sky130_fd_sc_hd__buf_2
XFILLER_89_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23027_ _23008_/X _23025_/Y _23027_/C VGND VGND VPWR VPWR _23027_/X sky130_fd_sc_hd__and3_4
X_20239_ _19913_/A HRDATA[31] VGND VGND VPWR VPWR _20239_/X sky130_fd_sc_hd__or2_4
XANTENNA__22600__A2 _22594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24371__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14800_ _14647_/X _14800_/B _14800_/C VGND VGND VPWR VPWR _14801_/C sky130_fd_sc_hd__and3_4
XFILLER_76_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15780_ _11755_/X _15776_/X _15779_/X VGND VGND VPWR VPWR _15781_/C sky130_fd_sc_hd__or3_4
X_12992_ _12876_/A _23752_/Q VGND VGND VPWR VPWR _12993_/C sky130_fd_sc_hd__or2_4
XANTENNA__21167__A2 _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18568__B1 _18563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22364__B2 _22359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14731_ _12502_/A _14731_/B VGND VGND VPWR VPWR _14732_/C sky130_fd_sc_hd__or2_4
X_11943_ _16116_/A VGND VGND VPWR VPWR _11943_/X sky130_fd_sc_hd__buf_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23929_ _23391_/CLK _21308_/X VGND VGND VPWR VPWR _14727_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18783__C _11633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17450_ _15786_/Y _18406_/B _17387_/Y _17449_/X VGND VGND VPWR VPWR _17450_/X sky130_fd_sc_hd__o22a_4
X_14662_ _11675_/A _14642_/X _14662_/C VGND VGND VPWR VPWR _14700_/B sky130_fd_sc_hd__or3_4
X_11874_ _13468_/A VGND VGND VPWR VPWR _16159_/A sky130_fd_sc_hd__buf_2
X_16401_ _12559_/A VGND VGND VPWR VPWR _16401_/X sky130_fd_sc_hd__buf_2
XANTENNA__22116__B2 _22106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13613_ _15018_/A VGND VGND VPWR VPWR _14297_/A sky130_fd_sc_hd__buf_2
X_17381_ _17493_/A _17381_/B VGND VGND VPWR VPWR _17381_/X sky130_fd_sc_hd__or2_4
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14593_ _14307_/A _23386_/Q VGND VGND VPWR VPWR _14595_/B sky130_fd_sc_hd__or2_4
XANTENNA__14385__A _14385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19120_ _19120_/A VGND VGND VPWR VPWR _19120_/Y sky130_fd_sc_hd__inv_2
X_16332_ _11714_/A VGND VGND VPWR VPWR _16333_/A sky130_fd_sc_hd__buf_2
XFILLER_111_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13544_ _13543_/X _23397_/Q VGND VGND VPWR VPWR _13544_/X sky130_fd_sc_hd__or2_4
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17543__A1 _17145_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19051_ _19038_/X _19050_/X _19038_/X _11530_/A VGND VGND VPWR VPWR _24356_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16263_ _11890_/X _16338_/B VGND VGND VPWR VPWR _16263_/X sky130_fd_sc_hd__or2_4
X_13475_ _13475_/A _13475_/B _13475_/C VGND VGND VPWR VPWR _13475_/X sky130_fd_sc_hd__or3_4
XFILLER_127_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_8_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22419__A2 _22414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18002_ _18035_/B _18001_/X VGND VGND VPWR VPWR _18002_/X sky130_fd_sc_hd__or2_4
X_15214_ _14669_/A _15143_/B VGND VGND VPWR VPWR _15214_/X sky130_fd_sc_hd__or2_4
XFILLER_51_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12426_ _12426_/A VGND VGND VPWR VPWR _12427_/A sky130_fd_sc_hd__buf_2
X_16194_ _11727_/A VGND VGND VPWR VPWR _16195_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21611__A2_N _21610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15145_ _13589_/A _15141_/X _15145_/C VGND VGND VPWR VPWR _15145_/X sky130_fd_sc_hd__or3_4
XFILLER_142_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12357_ _11712_/X _12357_/B VGND VGND VPWR VPWR _12357_/X sky130_fd_sc_hd__or2_4
XANTENNA__16105__A _15967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21946__A _21960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19953_ _19953_/A _19952_/Y VGND VGND VPWR VPWR _19953_/X sky130_fd_sc_hd__and2_4
X_15076_ _15076_/A VGND VGND VPWR VPWR _15096_/A sky130_fd_sc_hd__buf_2
X_12288_ _12288_/A VGND VGND VPWR VPWR _15442_/A sky130_fd_sc_hd__buf_2
X_18904_ _17266_/X _18897_/X _24401_/Q _18900_/X VGND VGND VPWR VPWR _24401_/D sky130_fd_sc_hd__o22a_4
X_14027_ _13719_/A _14025_/X _14027_/C VGND VGND VPWR VPWR _14027_/X sky130_fd_sc_hd__and3_4
XFILLER_68_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19884_ _19630_/X VGND VGND VPWR VPWR _19884_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18320__A _18320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18835_ _18834_/X VGND VGND VPWR VPWR _18835_/X sky130_fd_sc_hd__buf_2
XANTENNA__13464__A _13474_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15978_ _15978_/A _15978_/B _15978_/C VGND VGND VPWR VPWR _15978_/X sky130_fd_sc_hd__or3_4
X_18766_ _19965_/B _19964_/B VGND VGND VPWR VPWR _19962_/B sky130_fd_sc_hd__or2_4
XANTENNA__21158__A2 _21155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18559__B1 _18467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21681__A _21674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17717_ _16981_/A _17360_/X _16981_/A _17360_/X VGND VGND VPWR VPWR _17717_/X sky130_fd_sc_hd__a2bb2o_4
X_14929_ _14967_/A _14929_/B VGND VGND VPWR VPWR _14929_/X sky130_fd_sc_hd__or2_4
XANTENNA__20366__B1 _24465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18697_ _18696_/X VGND VGND VPWR VPWR _18697_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17648_ _17094_/Y VGND VGND VPWR VPWR _17648_/X sky130_fd_sc_hd__buf_2
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22107__B2 _22106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17579_ _17578_/X VGND VGND VPWR VPWR _18118_/B sky130_fd_sc_hd__inv_2
XANTENNA__12808__A _13530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14295__A _14295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11712__A _13248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19318_ _24278_/Q _19321_/A _19317_/Y VGND VGND VPWR VPWR _19318_/X sky130_fd_sc_hd__o21a_4
XFILLER_32_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20590_ _20589_/X VGND VGND VPWR VPWR _20590_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21330__A2 _21327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19249_ _24300_/Q _19248_/X VGND VGND VPWR VPWR _19250_/B sky130_fd_sc_hd__and2_4
XFILLER_104_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22260_ _22149_/X _22258_/X _13760_/B _22255_/X VGND VGND VPWR VPWR _22260_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22017__A _22010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21211_ _20633_/X _21205_/X _23973_/Q _21209_/X VGND VGND VPWR VPWR _23973_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17298__B1 _11855_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22191_ _22176_/A VGND VGND VPWR VPWR _22191_/X sky130_fd_sc_hd__buf_2
XFILLER_118_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15848__A1 _13307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21142_ _20337_/X _21141_/X _24019_/Q _21138_/X VGND VGND VPWR VPWR _24019_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21073_ _21033_/A VGND VGND VPWR VPWR _21073_/X sky130_fd_sc_hd__buf_2
XANTENNA__21397__A2 _21391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20024_ _18213_/X _20007_/X _20023_/Y _20018_/X VGND VGND VPWR VPWR _20024_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21149__A2 _21148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_14_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24181__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11637__A2 _11587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21975_ _21862_/X _21974_/X _23551_/Q _21971_/X VGND VGND VPWR VPWR _23551_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16685__A _11671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23714_ _23656_/CLK _23714_/D VGND VGND VPWR VPWR _23714_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20926_ _20926_/A VGND VGND VPWR VPWR _20926_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _23646_/CLK _21794_/X VGND VGND VPWR VPWR _23645_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22649__A2 _22644_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ _20857_/A _20856_/X VGND VGND VPWR VPWR _20857_/Y sky130_fd_sc_hd__nand2_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12718__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11622__A _12188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23576_ _23544_/CLK _23576_/D VGND VGND VPWR VPWR _15333_/B sky130_fd_sc_hd__dfxtp_4
X_11590_ _17060_/A _16921_/A VGND VGND VPWR VPWR _11590_/X sky130_fd_sc_hd__or2_4
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20788_ _20726_/X _20787_/Y _24287_/Q _20584_/X VGND VGND VPWR VPWR _20788_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12437__B _12579_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22527_ _22468_/X _22522_/X _14406_/B _22526_/X VGND VGND VPWR VPWR _22527_/X sky130_fd_sc_hd__o22a_4
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13260_ _12978_/A _13260_/B _13260_/C VGND VGND VPWR VPWR _13261_/C sky130_fd_sc_hd__or3_4
XANTENNA__24146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22458_ _22456_/X _22450_/X _15522_/B _22457_/X VGND VGND VPWR VPWR _22458_/X sky130_fd_sc_hd__o22a_4
X_12211_ _12691_/A _12211_/B _12211_/C VGND VGND VPWR VPWR _12225_/B sky130_fd_sc_hd__and3_4
XANTENNA__13549__A _13529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21409_ _21388_/A VGND VGND VPWR VPWR _21409_/X sky130_fd_sc_hd__buf_2
X_13191_ _13307_/A _13167_/X _13174_/X _13182_/X _13190_/X VGND VGND VPWR VPWR _13191_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12453__A _12453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22389_ _22144_/X _22383_/X _23296_/Q _22387_/X VGND VGND VPWR VPWR _23296_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20293__C1 _20292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12142_ _12166_/A _12142_/B VGND VGND VPWR VPWR _12142_/X sky130_fd_sc_hd__or2_4
X_24128_ _24184_/CLK _22739_/X HRESETn VGND VGND VPWR VPWR _24128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15764__A _12766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24059_ _23592_/CLK _24059_/D VGND VGND VPWR VPWR _24059_/Q sky130_fd_sc_hd__dfxtp_4
X_16950_ _17669_/A VGND VGND VPWR VPWR _16950_/Y sky130_fd_sc_hd__inv_2
X_12073_ _11951_/X _12073_/B _12073_/C VGND VGND VPWR VPWR _12074_/C sky130_fd_sc_hd__and3_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22585__B2 _22548_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15901_ _13547_/A _15899_/X _15900_/X VGND VGND VPWR VPWR _15902_/C sky130_fd_sc_hd__and3_4
X_16881_ _16855_/Y _16857_/B VGND VGND VPWR VPWR _16881_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__13284__A _12561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15832_ _12857_/A _15828_/X _15831_/X VGND VGND VPWR VPWR _15832_/X sky130_fd_sc_hd__or3_4
X_18620_ _17652_/X _18596_/X _16935_/A _18619_/X VGND VGND VPWR VPWR _18620_/X sky130_fd_sc_hd__o22a_4
XFILLER_106_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15763_ _15743_/X _15698_/B VGND VGND VPWR VPWR _15763_/X sky130_fd_sc_hd__or2_4
X_18551_ _18499_/X _18549_/X _18527_/X _18550_/X VGND VGND VPWR VPWR _18551_/X sky130_fd_sc_hd__o22a_4
X_12975_ _12975_/A _12975_/B _12974_/X VGND VGND VPWR VPWR _12975_/X sky130_fd_sc_hd__and3_4
XFILLER_79_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16595__A _16595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17502_ _13342_/Y _17020_/X _17028_/X _17501_/X VGND VGND VPWR VPWR _17503_/B sky130_fd_sc_hd__o22a_4
X_14714_ _14296_/A _14788_/B VGND VGND VPWR VPWR _14714_/X sky130_fd_sc_hd__or2_4
XFILLER_73_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18482_ _18481_/X VGND VGND VPWR VPWR _18482_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11926_ _16713_/A _11926_/B _11926_/C VGND VGND VPWR VPWR _11926_/X sky130_fd_sc_hd__and3_4
X_15694_ _13277_/A _15759_/B VGND VGND VPWR VPWR _15696_/B sky130_fd_sc_hd__or2_4
XFILLER_166_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14827__B _14827_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17433_ _17432_/X VGND VGND VPWR VPWR _17433_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14645_ _14684_/A _14645_/B VGND VGND VPWR VPWR _14646_/C sky130_fd_sc_hd__or2_4
X_11857_ _11857_/A VGND VGND VPWR VPWR _11858_/A sky130_fd_sc_hd__buf_2
XFILLER_166_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12628__A _12975_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17364_ _15653_/X _17445_/B VGND VGND VPWR VPWR _18466_/A sky130_fd_sc_hd__and2_4
XPHY_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14576_ _12444_/A _14574_/X _14575_/X VGND VGND VPWR VPWR _14580_/B sky130_fd_sc_hd__and3_4
XFILLER_159_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_34_0_HCLK clkbuf_7_34_0_HCLK/A VGND VGND VPWR VPWR _23983_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_14_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11788_ _12151_/A _23956_/Q VGND VGND VPWR VPWR _11788_/X sky130_fd_sc_hd__or2_4
XANTENNA__21312__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16315_ _11714_/A VGND VGND VPWR VPWR _16316_/A sky130_fd_sc_hd__buf_2
X_19103_ _19096_/X _19102_/X _19096_/X _11521_/A VGND VGND VPWR VPWR _24347_/D sky130_fd_sc_hd__a2bb2o_4
X_13527_ _12773_/X _13525_/X _13526_/X VGND VGND VPWR VPWR _13528_/C sky130_fd_sc_hd__and3_4
Xclkbuf_7_97_0_HCLK clkbuf_6_48_0_HCLK/X VGND VGND VPWR VPWR _23744_/CLK sky130_fd_sc_hd__clkbuf_1
X_17295_ _17294_/X VGND VGND VPWR VPWR _17301_/A sky130_fd_sc_hd__buf_2
XFILLER_159_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14843__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19034_ _19024_/X _19033_/X _19024_/X _24359_/Q VGND VGND VPWR VPWR _19034_/X sky130_fd_sc_hd__a2bb2o_4
X_16246_ _16246_/A _16246_/B VGND VGND VPWR VPWR _16528_/A sky130_fd_sc_hd__or2_4
X_13458_ _13462_/A _23621_/Q VGND VGND VPWR VPWR _13458_/X sky130_fd_sc_hd__or2_4
XFILLER_127_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13459__A _13431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12409_ _12339_/X _12407_/X _12409_/C VGND VGND VPWR VPWR _12409_/X sky130_fd_sc_hd__and3_4
XANTENNA__21076__B2 _21070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16177_ _16215_/A _16177_/B VGND VGND VPWR VPWR _16179_/B sky130_fd_sc_hd__or2_4
X_13389_ _13370_/A VGND VGND VPWR VPWR _13397_/A sky130_fd_sc_hd__buf_2
XANTENNA__12363__A _12923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24054__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15128_ _13788_/A _15128_/B _15127_/X VGND VGND VPWR VPWR _15128_/X sky130_fd_sc_hd__or3_4
Xclkbuf_3_3_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20580__A _11573_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15674__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22025__B1 _23519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19936_ _19931_/X _24171_/Q _19932_/X _20844_/A VGND VGND VPWR VPWR _24171_/D sky130_fd_sc_hd__o22a_4
X_15059_ _12322_/A _15059_/B VGND VGND VPWR VPWR _15059_/X sky130_fd_sc_hd__or2_4
XANTENNA__21379__A2 _21377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15393__B _15455_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19867_ _19562_/X _19857_/X _19859_/A _19898_/B VGND VGND VPWR VPWR _19867_/X sky130_fd_sc_hd__a211o_4
XANTENNA__13194__A _11675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18818_ _18789_/A VGND VGND VPWR VPWR _18818_/X sky130_fd_sc_hd__buf_2
XFILLER_96_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19798_ _19823_/B _19589_/X VGND VGND VPWR VPWR _19798_/X sky130_fd_sc_hd__and2_4
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18749_ _17986_/X _18747_/Y _17988_/X _18748_/Y VGND VGND VPWR VPWR _18749_/X sky130_fd_sc_hd__o22a_4
XFILLER_64_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13922__A _14377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21760_ _21767_/A VGND VGND VPWR VPWR _21760_/X sky130_fd_sc_hd__buf_2
XFILLER_93_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20711_ _20652_/A _20711_/B VGND VGND VPWR VPWR _20711_/Y sky130_fd_sc_hd__nor2_4
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12538__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21691_ _21658_/A VGND VGND VPWR VPWR _21691_/X sky130_fd_sc_hd__buf_2
X_23430_ _24102_/CLK _23430_/D VGND VGND VPWR VPWR _23430_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20642_ _20307_/X HRDATA[15] _20248_/B _20641_/X VGND VGND VPWR VPWR _20642_/X sky130_fd_sc_hd__a211o_4
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21303__A2 _21293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22500__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20573_ _24232_/Q _20534_/X _20572_/Y VGND VGND VPWR VPWR _22440_/A sky130_fd_sc_hd__o21a_4
X_23361_ _23617_/CLK _23361_/D VGND VGND VPWR VPWR _15525_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20511__B1 _12669_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14753__A _15446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18225__A _18283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22312_ _22291_/A VGND VGND VPWR VPWR _22312_/X sky130_fd_sc_hd__buf_2
XFILLER_118_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23292_ _23772_/CLK _22395_/X VGND VGND VPWR VPWR _14355_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22970__A _22969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13369__A _13378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21067__B2 _21063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22243_ _22120_/X _22237_/X _12819_/B _22241_/X VGND VGND VPWR VPWR _23402_/D sky130_fd_sc_hd__o22a_4
XFILLER_117_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22264__B1 _14462_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12273__A _12273_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11555__A1 _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12752__B1 _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22174_ _22173_/X VGND VGND VPWR VPWR _22208_/A sky130_fd_sc_hd__buf_2
XFILLER_133_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15584__A _15620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21125_ _21118_/A VGND VGND VPWR VPWR _21125_/X sky130_fd_sc_hd__buf_2
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22567__B2 _22562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21056_ _21049_/A VGND VGND VPWR VPWR _21056_/X sky130_fd_sc_hd__buf_2
XFILLER_154_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20007_ _19961_/X VGND VGND VPWR VPWR _20007_/X sky130_fd_sc_hd__buf_2
XFILLER_59_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11617__A _12466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17007__C _17906_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22319__A1 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21790__A2 _21784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22319__B2 _22284_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13832__A _15423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12625_/A VGND VGND VPWR VPWR _13055_/A sky130_fd_sc_hd__buf_2
X_21958_ _21833_/X _21953_/X _12514_/B _21957_/X VGND VGND VPWR VPWR _21958_/X sky130_fd_sc_hd__o22a_4
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _12372_/A VGND VGND VPWR VPWR _13248_/A sky130_fd_sc_hd__buf_2
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _18658_/Y _20702_/X _20753_/X _20908_/Y VGND VGND VPWR VPWR _20909_/X sky130_fd_sc_hd__a211o_4
X_12691_ _12691_/A _12691_/B _12690_/X VGND VGND VPWR VPWR _12691_/X sky130_fd_sc_hd__and3_4
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21889_ _21888_/X VGND VGND VPWR VPWR _21923_/A sky130_fd_sc_hd__buf_2
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A _23771_/Q VGND VGND VPWR VPWR _14431_/C sky130_fd_sc_hd__or2_4
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628_ _23500_/CLK _23628_/D VGND VGND VPWR VPWR _23628_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24327__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11642_ _11642_/A VGND VGND VPWR VPWR _11642_/X sky130_fd_sc_hd__buf_2
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20665__A _17077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _14512_/A _14359_/X _14360_/X VGND VGND VPWR VPWR _14361_/X sky130_fd_sc_hd__and3_4
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23559_ _23723_/CLK _23559_/D VGND VGND VPWR VPWR _23559_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20502__B1 _20638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11573_ _11573_/A IRQ[18] VGND VGND VPWR VPWR _20178_/A sky130_fd_sc_hd__and2_4
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14663__A _14663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16100_ _16099_/X VGND VGND VPWR VPWR _16101_/A sky130_fd_sc_hd__buf_2
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _13309_/A _13388_/B VGND VGND VPWR VPWR _13312_/X sky130_fd_sc_hd__or2_4
XFILLER_35_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17080_ _11643_/A _17077_/Y _11645_/X _17079_/Y VGND VGND VPWR VPWR _17090_/B sky130_fd_sc_hd__a211o_4
XFILLER_168_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14292_ _14292_/A _14292_/B _14292_/C VGND VGND VPWR VPWR _14292_/X sky130_fd_sc_hd__or3_4
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16031_ _16031_/A VGND VGND VPWR VPWR _16057_/A sky130_fd_sc_hd__buf_2
XANTENNA__21058__B2 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13279__A _13279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13243_ _13251_/A _13239_/X _13243_/C VGND VGND VPWR VPWR _13243_/X sky130_fd_sc_hd__or3_4
XFILLER_108_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17974__A _18413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21496__A _21489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13174_ _13338_/A _13170_/X _13173_/X VGND VGND VPWR VPWR _13174_/X sky130_fd_sc_hd__or3_4
XANTENNA__17693__B _17501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12125_ _16775_/A _23795_/Q VGND VGND VPWR VPWR _12126_/C sky130_fd_sc_hd__or2_4
XANTENNA__12911__A _12911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17982_ _17819_/X _17821_/X _17945_/X _17826_/X VGND VGND VPWR VPWR _17982_/X sky130_fd_sc_hd__o22a_4
XFILLER_97_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19721_ HRDATA[6] VGND VGND VPWR VPWR _19721_/Y sky130_fd_sc_hd__inv_2
X_16933_ _16932_/X VGND VGND VPWR VPWR _16933_/Y sky130_fd_sc_hd__inv_2
X_12056_ _11943_/X VGND VGND VPWR VPWR _12061_/A sky130_fd_sc_hd__buf_2
XFILLER_77_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20033__A2 _20031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19652_ _19623_/A _19624_/B VGND VGND VPWR VPWR _19857_/B sky130_fd_sc_hd__or2_4
XANTENNA__21230__B2 _21195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16864_ _15386_/X VGND VGND VPWR VPWR _16864_/Y sky130_fd_sc_hd__inv_2
X_18603_ _17594_/X _18603_/B VGND VGND VPWR VPWR _18603_/X sky130_fd_sc_hd__and2_4
XFILLER_65_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15815_ _12862_/A _15815_/B _15814_/X VGND VGND VPWR VPWR _15816_/C sky130_fd_sc_hd__and3_4
X_19583_ _19504_/B VGND VGND VPWR VPWR _19705_/A sky130_fd_sc_hd__buf_2
X_16795_ _16755_/X _16795_/B VGND VGND VPWR VPWR _16797_/B sky130_fd_sc_hd__or2_4
XANTENNA__22120__A _20530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14838__A _14658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15746_ _15770_/A _15746_/B VGND VGND VPWR VPWR _15746_/X sky130_fd_sc_hd__or2_4
X_18534_ _16978_/X VGND VGND VPWR VPWR _18534_/Y sky130_fd_sc_hd__inv_2
X_12958_ _12970_/A _23401_/Q VGND VGND VPWR VPWR _12960_/B sky130_fd_sc_hd__or2_4
XFILLER_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21533__A2 _21530_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22730__B2 _22726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11909_ _12466_/A VGND VGND VPWR VPWR _11910_/A sky130_fd_sc_hd__inv_2
X_15677_ _13338_/A _15677_/B _15676_/X VGND VGND VPWR VPWR _15677_/X sky130_fd_sc_hd__or3_4
X_18465_ _17920_/X _18319_/Y _17944_/X _18464_/X VGND VGND VPWR VPWR _18465_/X sky130_fd_sc_hd__a211o_4
X_12889_ _12889_/A _12889_/B _12889_/C VGND VGND VPWR VPWR _12890_/C sky130_fd_sc_hd__and3_4
XFILLER_34_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17416_ _17415_/Y _16926_/B _11891_/X _17043_/A VGND VGND VPWR VPWR _17416_/X sky130_fd_sc_hd__a2bb2o_4
X_14628_ _14693_/A _14624_/X _14628_/C VGND VGND VPWR VPWR _14629_/C sky130_fd_sc_hd__and3_4
XFILLER_18_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18396_ _18064_/X VGND VGND VPWR VPWR _18396_/X sky130_fd_sc_hd__buf_2
XFILLER_60_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15669__A _12704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17347_ _17339_/A _17340_/B _17341_/X _17346_/Y VGND VGND VPWR VPWR _17347_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14559_ _15398_/A _14555_/X _14559_/C VGND VGND VPWR VPWR _14559_/X sky130_fd_sc_hd__or3_4
XANTENNA__14573__A _14292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17278_ _11611_/B VGND VGND VPWR VPWR _17280_/A sky130_fd_sc_hd__inv_2
XFILLER_88_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23444__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16229_ _16205_/A _16229_/B _16228_/X VGND VGND VPWR VPWR _16237_/B sky130_fd_sc_hd__or3_4
XANTENNA__13189__A _11872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19017_ _11535_/A VGND VGND VPWR VPWR _19017_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12093__A _12001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13917__A _13877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12821__A _13349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22549__B2 _22548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19919_ _22931_/A VGND VGND VPWR VPWR _22738_/A sky130_fd_sc_hd__buf_2
XFILLER_151_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21221__B2 _21216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22930_ _22930_/A VGND VGND VPWR VPWR _22930_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21772__A2 _21770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22861_ _13049_/Y _22847_/X _22853_/X _22860_/X VGND VGND VPWR VPWR _22861_/X sky130_fd_sc_hd__a211o_4
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14748__A _11913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13652__A _13652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21812_ _21805_/Y _21810_/X _21811_/X _21810_/X VGND VGND VPWR VPWR _23636_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22792_ _22763_/Y _22792_/B VGND VGND VPWR VPWR _22792_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22965__A _22964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22721__B2 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21743_ _21580_/X _21741_/X _13741_/B _21738_/X VGND VGND VPWR VPWR _21743_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24491__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24462_ _23347_/CLK _24462_/D HRESETn VGND VGND VPWR VPWR _24462_/Q sky130_fd_sc_hd__dfrtp_4
X_21674_ _21674_/A VGND VGND VPWR VPWR _21674_/X sky130_fd_sc_hd__buf_2
XANTENNA__20485__A _20485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23413_ _23392_/CLK _23413_/D VGND VGND VPWR VPWR _23413_/Q sky130_fd_sc_hd__dfxtp_4
X_20625_ _20501_/A _20624_/X VGND VGND VPWR VPWR _20625_/Y sky130_fd_sc_hd__nor2_4
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22485__B1 _23253_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15579__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24393_ _24422_/CLK _24393_/D HRESETn VGND VGND VPWR VPWR _19020_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__14483__A _14482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23344_ _23533_/CLK _22326_/X VGND VGND VPWR VPWR _22326_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20556_ _20535_/X _20555_/X VGND VGND VPWR VPWR _20556_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_80_0_HCLK clkbuf_6_40_0_HCLK/X VGND VGND VPWR VPWR _23383_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_153_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13099__A _13099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23275_ _23531_/CLK _22434_/X VGND VGND VPWR VPWR _12579_/B sky130_fd_sc_hd__dfxtp_4
X_20487_ _20418_/X _20486_/X _24108_/Q _20396_/X VGND VGND VPWR VPWR _20487_/X sky130_fd_sc_hd__o22a_4
XFILLER_164_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22226_ _22226_/A VGND VGND VPWR VPWR _22226_/X sky130_fd_sc_hd__buf_2
XFILLER_156_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22205__A _22176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13827__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22157_ _22156_/X _22147_/X _14503_/B _22154_/X VGND VGND VPWR VPWR _23451_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21460__B2 _21459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16203__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12731__A _13301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21108_ _21101_/A VGND VGND VPWR VPWR _21108_/X sky130_fd_sc_hd__buf_2
XANTENNA__19405__A1 _19399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22088_ _11795_/B VGND VGND VPWR VPWR _22088_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17416__B1 _11891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13930_ _14507_/A _13930_/B VGND VGND VPWR VPWR _13930_/X sky130_fd_sc_hd__or2_4
X_21039_ _20337_/X _21038_/X _24083_/Q _21035_/X VGND VGND VPWR VPWR _24083_/D sky130_fd_sc_hd__o22a_4
XFILLER_101_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23036__A _22908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13861_ _15450_/A _13860_/X VGND VGND VPWR VPWR _13861_/X sky130_fd_sc_hd__and2_4
XANTENNA__14658__A _14658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15600_ _13894_/A _15591_/X _15600_/C VGND VGND VPWR VPWR _15600_/X sky130_fd_sc_hd__and3_4
XANTENNA__13562__A _13562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12812_ _12800_/A _12723_/B VGND VGND VPWR VPWR _12812_/X sky130_fd_sc_hd__or2_4
XFILLER_16_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17034__A _17481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23317__CLK _23456_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16580_ _16556_/A _16578_/X _16580_/C VGND VGND VPWR VPWR _16580_/X sky130_fd_sc_hd__and3_4
X_13792_ _13792_/A VGND VGND VPWR VPWR _15007_/A sky130_fd_sc_hd__buf_2
XFILLER_28_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21515__A2 _21513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15531_ _12236_/A _15529_/X _15531_/C VGND VGND VPWR VPWR _15535_/B sky130_fd_sc_hd__and3_4
XANTENNA__20098__C _20192_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12743_ _12240_/A _12824_/B VGND VGND VPWR VPWR _12743_/X sky130_fd_sc_hd__or2_4
XANTENNA__12178__A _16684_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18250_ _18250_/A _18249_/X VGND VGND VPWR VPWR _18251_/A sky130_fd_sc_hd__and2_4
X_15462_ _15486_/A _15399_/B VGND VGND VPWR VPWR _15462_/X sky130_fd_sc_hd__or2_4
XANTENNA__24161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12674_ _12976_/A _12674_/B _12673_/X VGND VGND VPWR VPWR _12675_/C sky130_fd_sc_hd__or3_4
XANTENNA__17688__B _17520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17128_/A _17195_/X _12093_/X _17200_/X VGND VGND VPWR VPWR _17202_/A sky130_fd_sc_hd__o22a_4
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14412_/X VGND VGND VPWR VPWR _14413_/Y sky130_fd_sc_hd__inv_2
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21279__B2 _21276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18181_ _18180_/X _17775_/D _17698_/X VGND VGND VPWR VPWR _18181_/X sky130_fd_sc_hd__o21a_4
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _11625_/A _11869_/A _12299_/A _11886_/A VGND VGND VPWR VPWR _11625_/X sky130_fd_sc_hd__or4_4
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _15393_/A _15455_/B VGND VGND VPWR VPWR _15393_/X sky130_fd_sc_hd__or2_4
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12906__A _12906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14393__A _14512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11810__A _11673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17132_ _16685_/X VGND VGND VPWR VPWR _17132_/Y sky130_fd_sc_hd__inv_2
X_14344_ _13937_/A VGND VGND VPWR VPWR _14367_/A sky130_fd_sc_hd__buf_2
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _11556_/A IRQ[20] VGND VGND VPWR VPWR _20180_/A sky130_fd_sc_hd__and2_4
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17063_ _11595_/A VGND VGND VPWR VPWR _20216_/D sky130_fd_sc_hd__buf_2
XANTENNA__15001__B _23989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14275_ _14280_/A _14275_/B _14275_/C VGND VGND VPWR VPWR _14276_/C sky130_fd_sc_hd__and3_4
X_16014_ _16130_/A _15987_/X _15994_/X _16003_/X _16013_/X VGND VGND VPWR VPWR _16014_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_170_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13226_ _12338_/X _13224_/X _13226_/C VGND VGND VPWR VPWR _13227_/C sky130_fd_sc_hd__and3_4
XFILLER_174_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22115__A _20485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13157_ _12301_/A _13157_/B _13157_/C VGND VGND VPWR VPWR _13158_/C sky130_fd_sc_hd__and3_4
XANTENNA__21451__B2 _21445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12641__A _12641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12108_ _12108_/A _12104_/X _12107_/X VGND VGND VPWR VPWR _12109_/B sky130_fd_sc_hd__or3_4
XFILLER_111_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13088_ _13088_/A _23336_/Q VGND VGND VPWR VPWR _13090_/B sky130_fd_sc_hd__or2_4
X_17965_ _17904_/X _16996_/B VGND VGND VPWR VPWR _17965_/X sky130_fd_sc_hd__and2_4
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19704_ _20844_/A _19573_/X _19703_/X _19638_/X VGND VGND VPWR VPWR _19704_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21203__B2 _21202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16916_ _17060_/A VGND VGND VPWR VPWR _16918_/A sky130_fd_sc_hd__inv_2
X_12039_ _16704_/A _12119_/B VGND VGND VPWR VPWR _12039_/X sky130_fd_sc_hd__or2_4
XFILLER_66_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17958__A1 _16943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17896_ _17781_/X _17895_/X _17781_/X _17895_/X VGND VGND VPWR VPWR _17896_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17958__B2 _17957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21754__A2 _21727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19635_ _19571_/X _19611_/X _19634_/X _17274_/A _19607_/X VGND VGND VPWR VPWR _24207_/D
+ sky130_fd_sc_hd__a32o_4
X_16847_ _15391_/A _13950_/X _15391_/D VGND VGND VPWR VPWR _16848_/B sky130_fd_sc_hd__or3_4
XANTENNA__14568__A _13601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13472__A _13441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19566_ HRDATA[29] VGND VGND VPWR VPWR _20339_/B sky130_fd_sc_hd__buf_2
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16778_ _16768_/A _16778_/B _16777_/X VGND VGND VPWR VPWR _16778_/X sky130_fd_sc_hd__or3_4
XFILLER_168_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22703__B2 _22698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18517_ _18517_/A VGND VGND VPWR VPWR _18518_/A sky130_fd_sc_hd__inv_2
X_15729_ _12780_/X _24036_/Q VGND VGND VPWR VPWR _15729_/X sky130_fd_sc_hd__or2_4
X_19497_ _24178_/Q _19457_/A HRDATA[30] _19454_/A VGND VGND VPWR VPWR _19497_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16783__A _16611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19580__B1 HRDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24348__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18448_ _18437_/X _18442_/Y _18444_/X _18446_/X _18447_/Y VGND VGND VPWR VPWR _18448_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15399__A _14307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22467__B1 _13796_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18379_ _18314_/A _18379_/B _18379_/C _18379_/D VGND VGND VPWR VPWR _18379_/X sky130_fd_sc_hd__or4_4
XFILLER_144_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20410_ _20409_/X VGND VGND VPWR VPWR _20410_/Y sky130_fd_sc_hd__inv_2
X_21390_ _21266_/X _21384_/X _12747_/B _21388_/X VGND VGND VPWR VPWR _21390_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12535__B _23979_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20341_ _20261_/X VGND VGND VPWR VPWR _20341_/X sky130_fd_sc_hd__buf_2
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23060_ _18011_/X _23079_/B VGND VGND VPWR VPWR _23061_/C sky130_fd_sc_hd__or2_4
X_20272_ _20490_/A VGND VGND VPWR VPWR _20273_/A sky130_fd_sc_hd__buf_2
XFILLER_161_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22011_ _21838_/X _22010_/X _12916_/B _22007_/X VGND VGND VPWR VPWR _22011_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17646__B1 _17594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13647__A _15444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21442__B2 _21438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12270__B _23980_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19334__A _23083_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23962_ _24057_/CLK _21227_/X VGND VGND VPWR VPWR _14584_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22913_ _22912_/X VGND VGND VPWR VPWR _23080_/A sky130_fd_sc_hd__buf_2
XFILLER_29_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23893_ _23456_/CLK _23893_/D VGND VGND VPWR VPWR _23893_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22844_ _15785_/A _22836_/X _22817_/X _22843_/X VGND VGND VPWR VPWR _22845_/B sky130_fd_sc_hd__o22a_4
XFILLER_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22775_ _24117_/D VGND VGND VPWR VPWR _22790_/C sky130_fd_sc_hd__inv_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22170__A2 _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21726_ _21551_/X _21720_/X _23690_/Q _21724_/X VGND VGND VPWR VPWR _21726_/X sky130_fd_sc_hd__o22a_4
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20181__A1 _24458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21104__A _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24445_ _24445_/CLK _24445_/D HRESETn VGND VGND VPWR VPWR _24445_/Q sky130_fd_sc_hd__dfrtp_4
X_21657_ _21656_/X VGND VGND VPWR VPWR _21658_/A sky130_fd_sc_hd__buf_2
XANTENNA__12726__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20608_ _20608_/A VGND VGND VPWR VPWR _20608_/Y sky130_fd_sc_hd__inv_2
X_12390_ _12829_/A _12390_/B VGND VGND VPWR VPWR _12391_/C sky130_fd_sc_hd__or2_4
X_24376_ _24388_/CLK _18939_/X HRESETn VGND VGND VPWR VPWR _24376_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_149_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21588_ _21587_/X _21578_/X _23771_/Q _21585_/X VGND VGND VPWR VPWR _21588_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21130__B1 _14859_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23327_ _23671_/CLK _22343_/X VGND VGND VPWR VPWR _14117_/B sky130_fd_sc_hd__dfxtp_4
X_20539_ _20287_/A VGND VGND VPWR VPWR _20539_/X sky130_fd_sc_hd__buf_2
XFILLER_119_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18413__A _18413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14060_ _13705_/A _23840_/Q VGND VGND VPWR VPWR _14061_/C sky130_fd_sc_hd__or2_4
X_23258_ _23194_/CLK _23258_/D VGND VGND VPWR VPWR _14618_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_134_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13011_ _13011_/A _13009_/X _13011_/C VGND VGND VPWR VPWR _13015_/B sky130_fd_sc_hd__and3_4
XANTENNA__13557__A _13543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22209_ _22146_/X _22208_/X _23423_/Q _22205_/X VGND VGND VPWR VPWR _22209_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21433__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17029__A _17028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22630__B1 _14649_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12461__A _12461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23189_ _23904_/CLK _22585_/X VGND VGND VPWR VPWR _15059_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21984__A2 _21981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15772__A _11739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17750_ _24131_/Q VGND VGND VPWR VPWR _17751_/A sky130_fd_sc_hd__inv_2
X_14962_ _14970_/A _14891_/B VGND VGND VPWR VPWR _14962_/X sky130_fd_sc_hd__or2_4
XANTENNA__24265__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21736__A2 _21734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16701_ _16724_/A _16766_/B VGND VGND VPWR VPWR _16701_/X sky130_fd_sc_hd__or2_4
XFILLER_101_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13913_ _14386_/A _13831_/B VGND VGND VPWR VPWR _13913_/X sky130_fd_sc_hd__or2_4
X_17681_ _17681_/A _17456_/Y VGND VGND VPWR VPWR _17681_/X sky130_fd_sc_hd__or2_4
X_14893_ _14991_/A _14893_/B _14892_/X VGND VGND VPWR VPWR _14893_/X sky130_fd_sc_hd__or3_4
XFILLER_74_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11805__A _11836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19420_ _19418_/X _18503_/Y _19418_/X _24224_/Q VGND VGND VPWR VPWR _19420_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16632_ _16654_/A _23954_/Q VGND VGND VPWR VPWR _16632_/X sky130_fd_sc_hd__or2_4
X_13844_ _15412_/A _13844_/B _13844_/C VGND VGND VPWR VPWR _13844_/X sky130_fd_sc_hd__or3_4
XFILLER_16_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19351_ _19347_/X _18274_/X _19350_/X _24265_/Q VGND VGND VPWR VPWR _19351_/X sky130_fd_sc_hd__a2bb2o_4
X_13775_ _12623_/A _13775_/B VGND VGND VPWR VPWR _13775_/X sky130_fd_sc_hd__or2_4
X_16563_ _12015_/A _23602_/Q VGND VGND VPWR VPWR _16564_/C sky130_fd_sc_hd__or2_4
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18302_ _17696_/X _18302_/B VGND VGND VPWR VPWR _18302_/X sky130_fd_sc_hd__and2_4
X_12726_ _12726_/A _12722_/X _12726_/C VGND VGND VPWR VPWR _12726_/X sky130_fd_sc_hd__or3_4
X_15514_ _13063_/A _15510_/X _15513_/X VGND VGND VPWR VPWR _15514_/X sky130_fd_sc_hd__or3_4
X_16494_ _16481_/X _16425_/B VGND VGND VPWR VPWR _16495_/C sky130_fd_sc_hd__or2_4
X_19282_ _24296_/Q _19245_/B _19281_/Y VGND VGND VPWR VPWR _19282_/X sky130_fd_sc_hd__o21a_4
XFILLER_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14835__B _14751_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15445_ _11878_/A _15445_/B _15444_/X VGND VGND VPWR VPWR _15445_/X sky130_fd_sc_hd__and3_4
X_18233_ _17460_/X _18164_/X VGND VGND VPWR VPWR _18233_/X sky130_fd_sc_hd__or2_4
X_12657_ _12943_/A _12657_/B VGND VGND VPWR VPWR _12658_/C sky130_fd_sc_hd__or2_4
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ _11608_/A VGND VGND VPWR VPWR _11608_/X sky130_fd_sc_hd__buf_2
XANTENNA__15012__A _12467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15376_ _11752_/A _15376_/B _15375_/X VGND VGND VPWR VPWR _15377_/C sky130_fd_sc_hd__or3_4
X_18164_ _17638_/Y _17605_/X _17603_/X VGND VGND VPWR VPWR _18164_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21121__B1 _24029_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12588_ _15457_/A VGND VGND VPWR VPWR _12925_/A sky130_fd_sc_hd__buf_2
XFILLER_157_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17115_ _17197_/A VGND VGND VPWR VPWR _17115_/X sky130_fd_sc_hd__buf_2
X_14327_ _12469_/A _14327_/B _14326_/X VGND VGND VPWR VPWR _14327_/X sky130_fd_sc_hd__and3_4
XANTENNA__15947__A _15971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11539_ _18994_/A _18995_/A VGND VGND VPWR VPWR _11540_/B sky130_fd_sc_hd__or2_4
X_18095_ _18095_/A VGND VGND VPWR VPWR _18095_/X sky130_fd_sc_hd__buf_2
XFILLER_171_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21672__B2 _21667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14851__A _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17046_ _17046_/A VGND VGND VPWR VPWR _17047_/A sky130_fd_sc_hd__buf_2
XFILLER_116_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14258_ _11680_/A _14250_/X _14258_/C VGND VGND VPWR VPWR _14258_/X sky130_fd_sc_hd__and3_4
XFILLER_125_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13467__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13209_ _13223_/A _13207_/X _13208_/X VGND VGND VPWR VPWR _13210_/C sky130_fd_sc_hd__and3_4
XANTENNA__22621__B1 _23168_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14189_ _14226_/A VGND VGND VPWR VPWR _14200_/A sky130_fd_sc_hd__buf_2
XFILLER_139_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21975__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21684__A _21677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18997_ _24397_/Q VGND VGND VPWR VPWR _18997_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16778__A _16768_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17948_ _17813_/X _17947_/Y _17240_/X VGND VGND VPWR VPWR _17948_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17879_ _17878_/X _17190_/Y _17240_/X VGND VGND VPWR VPWR _17879_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14298__A _13617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19618_ _19446_/A _19617_/X HRDATA[3] _19461_/X VGND VGND VPWR VPWR _19619_/A sky130_fd_sc_hd__o22a_4
X_20890_ _24219_/Q _20773_/X _20889_/X VGND VGND VPWR VPWR _22471_/A sky130_fd_sc_hd__o21a_4
X_19549_ _19545_/A _19848_/A _19883_/A _19548_/X VGND VGND VPWR VPWR _19550_/D sky130_fd_sc_hd__a211o_4
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22152__A2 _22147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13930__A _14507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22560_ _22440_/X _22558_/X _12995_/B _22555_/X VGND VGND VPWR VPWR _23208_/D sky130_fd_sc_hd__o22a_4
XFILLER_62_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18217__B _18148_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21511_ _21299_/X _21506_/X _14397_/B _21510_/X VGND VGND VPWR VPWR _23804_/D sky130_fd_sc_hd__o22a_4
XFILLER_139_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22491_ _22498_/A VGND VGND VPWR VPWR _22491_/X sky130_fd_sc_hd__buf_2
XFILLER_166_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12546__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24230_ _24134_/CLK _19412_/X HRESETn VGND VGND VPWR VPWR _24230_/Q sky130_fd_sc_hd__dfrtp_4
X_21442_ _21268_/X _21441_/X _23849_/Q _21438_/X VGND VGND VPWR VPWR _21442_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19856__A1 _19823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24138__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15857__A _12373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24161_ _24472_/CLK _19987_/Y HRESETn VGND VGND VPWR VPWR _24161_/Q sky130_fd_sc_hd__dfrtp_4
X_21373_ _21388_/A VGND VGND VPWR VPWR _21381_/A sky130_fd_sc_hd__buf_2
X_23112_ _23880_/CLK _23112_/D VGND VGND VPWR VPWR _13109_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20324_ _20273_/A _20322_/Y _24307_/Q _20323_/X VGND VGND VPWR VPWR _20324_/X sky130_fd_sc_hd__o22a_4
X_24092_ _23592_/CLK _20862_/X VGND VGND VPWR VPWR _24092_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13377__A _13377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23043_ _23043_/A _23043_/B VGND VGND VPWR VPWR _23043_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21415__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12281__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20255_ _20255_/A VGND VGND VPWR VPWR _20255_/X sky130_fd_sc_hd__buf_2
XANTENNA__24288__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21966__A2 _21960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20186_ _20186_/A _20185_/Y VGND VGND VPWR VPWR _20186_/X sky130_fd_sc_hd__or2_4
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18831__A2 _18796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21718__A2 _21713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22915__A1 _18717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23945_ _24073_/CLK _21270_/X VGND VGND VPWR VPWR _23945_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22391__A2 _22390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11625__A _11625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11890_ _11889_/X VGND VGND VPWR VPWR _11890_/X sky130_fd_sc_hd__buf_2
X_23876_ _23523_/CLK _21399_/X VGND VGND VPWR VPWR _15712_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14001__A _11623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22827_ _17425_/Y _22816_/X _22818_/X _22826_/X VGND VGND VPWR VPWR _22827_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14936__A _14772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22143__A2 _22135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13560_ _13515_/X _23237_/Q VGND VGND VPWR VPWR _13562_/B sky130_fd_sc_hd__or2_4
X_22758_ SYSTICKCLKDIV[1] VGND VGND VPWR VPWR _22758_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21351__B1 _23906_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12511_ _12511_/A _23339_/Q VGND VGND VPWR VPWR _12515_/B sky130_fd_sc_hd__or2_4
X_21709_ _21724_/A VGND VGND VPWR VPWR _21717_/A sky130_fd_sc_hd__buf_2
X_13491_ _13542_/A _13488_/X _13490_/X VGND VGND VPWR VPWR _13491_/X sky130_fd_sc_hd__and3_4
XANTENNA__12456__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22689_ _22722_/A VGND VGND VPWR VPWR _22705_/A sky130_fd_sc_hd__inv_2
XFILLER_13_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15230_ _14200_/A _15166_/B VGND VGND VPWR VPWR _15230_/X sky130_fd_sc_hd__or2_4
XANTENNA__24394__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12442_ _13955_/A VGND VGND VPWR VPWR _15018_/A sky130_fd_sc_hd__buf_2
X_24428_ _24428_/CLK _18854_/X HRESETn VGND VGND VPWR VPWR _24428_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15581__A1 _11969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15161_ _14277_/A _15157_/X _15160_/X VGND VGND VPWR VPWR _15161_/X sky130_fd_sc_hd__or3_4
XFILLER_60_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12373_ _12948_/A VGND VGND VPWR VPWR _12373_/X sky130_fd_sc_hd__buf_2
XANTENNA__22851__B1 _22884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24359_ _24398_/CLK _19034_/X HRESETn VGND VGND VPWR VPWR _24359_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21654__B2 _21617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23505__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_50_0_HCLK clkbuf_6_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14112_ _12426_/A _14112_/B _14111_/X VGND VGND VPWR VPWR _14112_/X sky130_fd_sc_hd__and3_4
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15486__B _23906_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15092_ _15075_/A _23125_/Q VGND VGND VPWR VPWR _15092_/X sky130_fd_sc_hd__or2_4
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18920_ _18896_/A VGND VGND VPWR VPWR _18920_/X sky130_fd_sc_hd__buf_2
X_14043_ _14056_/A _24000_/Q VGND VGND VPWR VPWR _14043_/X sky130_fd_sc_hd__or2_4
XANTENNA__12191__A _12191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18851_ _16381_/X _18849_/X _24431_/Q _18850_/X VGND VGND VPWR VPWR _24431_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23655__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16598__A _12001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17802_ _17801_/X _17256_/X VGND VGND VPWR VPWR _17803_/D sky130_fd_sc_hd__and2_4
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18782_ _17048_/A _18782_/B _17406_/Y _17398_/Y VGND VGND VPWR VPWR _18834_/C sky130_fd_sc_hd__or4_4
X_15994_ _15971_/A _15994_/B _15994_/C VGND VGND VPWR VPWR _15994_/X sky130_fd_sc_hd__or3_4
X_17733_ _17732_/A _17276_/X VGND VGND VPWR VPWR _17735_/A sky130_fd_sc_hd__and2_4
X_14945_ _14976_/A _14867_/B VGND VGND VPWR VPWR _14945_/X sky130_fd_sc_hd__or2_4
XFILLER_48_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22382__A2 _22376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19702__A HRDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17664_ _16949_/A _17558_/X _17661_/X VGND VGND VPWR VPWR _17664_/Y sky130_fd_sc_hd__o21ai_4
X_14876_ _13591_/A _14874_/X _14875_/X VGND VGND VPWR VPWR _14876_/X sky130_fd_sc_hd__and3_4
XFILLER_21_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19403_ _19399_/X _19400_/Y _19402_/X _24235_/Q VGND VGND VPWR VPWR _24235_/D sky130_fd_sc_hd__o22a_4
X_16615_ _16654_/A _16615_/B VGND VGND VPWR VPWR _16615_/X sky130_fd_sc_hd__or2_4
X_13827_ _13622_/A _13825_/X _13826_/X VGND VGND VPWR VPWR _13827_/X sky130_fd_sc_hd__and3_4
X_17595_ _17569_/X _18118_/B _17571_/A VGND VGND VPWR VPWR _17595_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__14846__A _14766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19334_ _23083_/D VGND VGND VPWR VPWR _20200_/A sky130_fd_sc_hd__buf_2
XFILLER_16_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13758_ _12583_/A _13758_/B VGND VGND VPWR VPWR _13759_/C sky130_fd_sc_hd__or2_4
X_16546_ _11951_/A VGND VGND VPWR VPWR _16556_/A sky130_fd_sc_hd__buf_2
X_12709_ _12228_/A _12789_/B VGND VGND VPWR VPWR _12709_/X sky130_fd_sc_hd__or2_4
X_19265_ _19254_/B VGND VGND VPWR VPWR _19265_/Y sky130_fd_sc_hd__inv_2
X_16477_ _16163_/X _16475_/X _16476_/X VGND VGND VPWR VPWR _16478_/C sky130_fd_sc_hd__and3_4
XANTENNA__12366__A _15887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21893__B2 _21892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13689_ _13689_/A _13688_/X VGND VGND VPWR VPWR _13689_/X sky130_fd_sc_hd__and2_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18216_ _18190_/A _18217_/C _16991_/B VGND VGND VPWR VPWR _18216_/X sky130_fd_sc_hd__o21a_4
X_15428_ _15405_/A _15428_/B _15427_/X VGND VGND VPWR VPWR _15428_/X sky130_fd_sc_hd__or3_4
X_19196_ _19144_/A _19143_/X _19195_/Y VGND VGND VPWR VPWR _19196_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15677__A _13338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18147_ _17702_/A _18148_/C _18107_/A VGND VGND VPWR VPWR _23038_/B sky130_fd_sc_hd__o21a_4
X_15359_ _13704_/A _23416_/Q VGND VGND VPWR VPWR _15359_/X sky130_fd_sc_hd__or2_4
XFILLER_157_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14581__A _14302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23185__CLK _23281_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15396__B _23746_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18078_ _17801_/X _17569_/X VGND VGND VPWR VPWR _18079_/D sky130_fd_sc_hd__and2_4
XFILLER_132_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17029_ _17028_/X VGND VGND VPWR VPWR _17029_/X sky130_fd_sc_hd__buf_2
XFILLER_144_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21948__A2 _21946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20040_ _18670_/A VGND VGND VPWR VPWR _20040_/X sky130_fd_sc_hd__buf_2
XANTENNA__22070__B2 _22064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21991_ _21991_/A VGND VGND VPWR VPWR _22007_/A sky130_fd_sc_hd__inv_2
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23730_ _23728_/CLK _23730_/D VGND VGND VPWR VPWR _23730_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20942_ _20864_/X _20940_/X _20941_/X HRDATA[11] _20869_/X VGND VGND VPWR VPWR _20942_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_82_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _23501_/CLK _21772_/X VGND VGND VPWR VPWR _16150_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _20873_/A VGND VGND VPWR VPWR _20873_/X sky130_fd_sc_hd__buf_2
XFILLER_42_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14756__A _12288_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22612_ _22605_/A VGND VGND VPWR VPWR _22612_/X sky130_fd_sc_hd__buf_2
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23592_ _23592_/CLK _21911_/X VGND VGND VPWR VPWR _23592_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22973__A _18494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22543_ _22539_/A VGND VGND VPWR VPWR _22558_/A sky130_fd_sc_hd__buf_2
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21884__B2 _21809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12276__A _12727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24404__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11611__C _11611_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22474_ _22462_/A VGND VGND VPWR VPWR _22474_/X sky130_fd_sc_hd__buf_2
X_24213_ _24471_/CLK _24213_/D HRESETn VGND VGND VPWR VPWR _24213_/Q sky130_fd_sc_hd__dfrtp_4
X_21425_ _21419_/Y _21424_/X _21241_/X _21424_/X VGND VGND VPWR VPWR _23860_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21636__B2 _21631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14491__A _12372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24144_ _24127_/CLK _20069_/Y HRESETn VGND VGND VPWR VPWR _16962_/A sky130_fd_sc_hd__dfrtp_4
X_21356_ _21292_/X _21355_/X _23903_/Q _21352_/X VGND VGND VPWR VPWR _23903_/D sky130_fd_sc_hd__o22a_4
XFILLER_162_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20307_ _18779_/X VGND VGND VPWR VPWR _20307_/X sky130_fd_sc_hd__buf_2
X_24075_ _24074_/CLK _21050_/X VGND VGND VPWR VPWR _12647_/B sky130_fd_sc_hd__dfxtp_4
X_21287_ _20745_/A VGND VGND VPWR VPWR _21287_/X sky130_fd_sc_hd__buf_2
XANTENNA__20940__B _20561_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22061__A1 _21838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23026_ _18238_/X _23003_/B VGND VGND VPWR VPWR _23027_/C sky130_fd_sc_hd__or2_4
XFILLER_89_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22061__B2 _22057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20238_ _20241_/A _20844_/A VGND VGND VPWR VPWR _20238_/X sky130_fd_sc_hd__or2_4
XFILLER_103_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13835__A _14319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17307__A _17272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20169_ _20169_/A VGND VGND VPWR VPWR _20169_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18017__B1 _17653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12991_ _12875_/A _12991_/B VGND VGND VPWR VPWR _12991_/X sky130_fd_sc_hd__or2_4
XFILLER_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22364__A2 _22362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14730_ _12495_/A _14798_/B VGND VGND VPWR VPWR _14730_/X sky130_fd_sc_hd__or2_4
XFILLER_91_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11942_ _16713_/A _11942_/B _11942_/C VGND VGND VPWR VPWR _11948_/B sky130_fd_sc_hd__and3_4
X_23928_ _23864_/CLK _23928_/D VGND VGND VPWR VPWR _23928_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23044__A _18140_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14661_ _13928_/A _14652_/X _14660_/X VGND VGND VPWR VPWR _14662_/C sky130_fd_sc_hd__and3_4
X_11873_ _12857_/A VGND VGND VPWR VPWR _13468_/A sky130_fd_sc_hd__buf_2
X_23859_ _23119_/CLK _23859_/D VGND VGND VPWR VPWR _23859_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24303__CLK _24306_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18783__D _18834_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22116__A2 _22111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16400_ _15978_/A _16396_/X _16399_/X VGND VGND VPWR VPWR _16400_/X sky130_fd_sc_hd__or3_4
X_13612_ _11932_/A VGND VGND VPWR VPWR _15405_/A sky130_fd_sc_hd__buf_2
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17380_ _16611_/A _17378_/X _17379_/X VGND VGND VPWR VPWR _17381_/B sky130_fd_sc_hd__o21a_4
X_14592_ _15394_/A _14590_/X _14591_/X VGND VGND VPWR VPWR _14592_/X sky130_fd_sc_hd__and3_4
X_13543_ _12970_/A VGND VGND VPWR VPWR _13543_/X sky130_fd_sc_hd__buf_2
X_16331_ _16314_/X _16331_/B _16330_/X VGND VGND VPWR VPWR _16331_/X sky130_fd_sc_hd__and3_4
XANTENNA__12186__A _12186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18740__B2 _22846_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16262_ _16129_/A _16262_/B _16261_/X VGND VGND VPWR VPWR _16262_/X sky130_fd_sc_hd__or3_4
XANTENNA__21499__A _21492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19050_ _19046_/X _19047_/Y _19048_/Y _19049_/X VGND VGND VPWR VPWR _19050_/X sky130_fd_sc_hd__o22a_4
X_13474_ _13474_/A _13472_/X _13474_/C VGND VGND VPWR VPWR _13475_/C sky130_fd_sc_hd__and3_4
XFILLER_40_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15213_ _14677_/A _15213_/B VGND VGND VPWR VPWR _15215_/B sky130_fd_sc_hd__or2_4
X_18001_ _17640_/X _17641_/C _17595_/Y VGND VGND VPWR VPWR _18001_/X sky130_fd_sc_hd__o21a_4
X_12425_ _12425_/A VGND VGND VPWR VPWR _12426_/A sky130_fd_sc_hd__buf_2
X_16193_ _16202_/A _16193_/B VGND VGND VPWR VPWR _16193_/X sky130_fd_sc_hd__or2_4
XFILLER_126_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15144_ _12444_/A _15142_/X _15144_/C VGND VGND VPWR VPWR _15145_/C sky130_fd_sc_hd__and3_4
X_12356_ _13258_/A VGND VGND VPWR VPWR _15887_/A sky130_fd_sc_hd__buf_2
XFILLER_154_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19952_ _19951_/X VGND VGND VPWR VPWR _19952_/Y sky130_fd_sc_hd__inv_2
X_15075_ _15075_/A _23669_/Q VGND VGND VPWR VPWR _15075_/X sky130_fd_sc_hd__or2_4
X_12287_ _12287_/A VGND VGND VPWR VPWR _12288_/A sky130_fd_sc_hd__buf_2
XFILLER_141_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18903_ _17255_/X _18897_/X _24402_/Q _18900_/X VGND VGND VPWR VPWR _18903_/X sky130_fd_sc_hd__o22a_4
X_14026_ _13705_/A _23776_/Q VGND VGND VPWR VPWR _14027_/C sky130_fd_sc_hd__or2_4
XFILLER_136_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22052__B2 _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19883_ _19883_/A _19690_/B VGND VGND VPWR VPWR _19903_/A sky130_fd_sc_hd__or2_4
XANTENNA__22123__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13745__A _12610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18834_ _11609_/X _18888_/B _18834_/C _18834_/D VGND VGND VPWR VPWR _18834_/X sky130_fd_sc_hd__or4_4
XFILLER_1_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_57_0_HCLK clkbuf_7_57_0_HCLK/A VGND VGND VPWR VPWR _23531_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18765_ _12024_/A _19963_/B VGND VGND VPWR VPWR _19964_/B sky130_fd_sc_hd__and2_4
X_15977_ _16006_/A _15977_/B _15977_/C VGND VGND VPWR VPWR _15978_/C sky130_fd_sc_hd__and3_4
XANTENNA__18559__A1 _18413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17716_ _16981_/A VGND VGND VPWR VPWR _18478_/A sky130_fd_sc_hd__buf_2
X_14928_ _12327_/A VGND VGND VPWR VPWR _14967_/A sky130_fd_sc_hd__buf_2
X_18696_ _18506_/X _18688_/X _18689_/Y _18691_/X _18695_/Y VGND VGND VPWR VPWR _18696_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17647_ _17085_/A _17647_/B VGND VGND VPWR VPWR _17647_/Y sky130_fd_sc_hd__nand2_4
X_14859_ _14096_/A _14859_/B VGND VGND VPWR VPWR _14862_/B sky130_fd_sc_hd__or2_4
XANTENNA__22107__A2 _22099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14576__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17578_ _16242_/X _18114_/B VGND VGND VPWR VPWR _17578_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19317_ _19227_/X VGND VGND VPWR VPWR _19317_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21866__A1 _21865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16529_ _16086_/X _16244_/Y _16088_/A VGND VGND VPWR VPWR _16529_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21866__B2 _21858_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12096__A _12093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19248_ _24299_/Q _19248_/B VGND VGND VPWR VPWR _19248_/X sky130_fd_sc_hd__and2_4
XFILLER_91_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21202__A _21202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21618__B2 _21617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19179_ _19153_/B VGND VGND VPWR VPWR _19179_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12824__A _12800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21210_ _20613_/X _21205_/X _23974_/Q _21209_/X VGND VGND VPWR VPWR _23974_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15200__A _14616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22190_ _22115_/X _22187_/X _12393_/B _22184_/X VGND VGND VPWR VPWR _23436_/D sky130_fd_sc_hd__o22a_4
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21141_ _21155_/A VGND VGND VPWR VPWR _21141_/X sky130_fd_sc_hd__buf_2
XANTENNA__24445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21072_ _20892_/X _21066_/X _24059_/Q _21070_/X VGND VGND VPWR VPWR _24059_/D sky130_fd_sc_hd__o22a_4
XFILLER_59_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18798__A1 _16381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20023_ _20023_/A VGND VGND VPWR VPWR _20023_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17127__A _12061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13655__A _13655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21872__A _20892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23200__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24326__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21974_ _21941_/A VGND VGND VPWR VPWR _21974_/X sky130_fd_sc_hd__buf_2
XFILLER_55_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23713_ _23649_/CLK _21689_/X VGND VGND VPWR VPWR _23713_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20925_ _20447_/A _20922_/Y _20924_/X _19111_/Y _20731_/X VGND VGND VPWR VPWR _20926_/A
+ sky130_fd_sc_hd__a32o_4
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14486__A _12410_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17773__A2 _17493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13390__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11903__A _13427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23644_ _23675_/CLK _21796_/X VGND VGND VPWR VPWR _23644_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24476__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20856_ _20695_/X _20846_/Y _20854_/X _20855_/Y _20714_/X VGND VGND VPWR VPWR _20856_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23575_ _23511_/CLK _21934_/X VGND VGND VPWR VPWR _15147_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20787_ _20787_/A VGND VGND VPWR VPWR _20787_/Y sky130_fd_sc_hd__inv_2
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22526_ _22505_/A VGND VGND VPWR VPWR _22526_/X sky130_fd_sc_hd__buf_2
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22208__A _22208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22457_ _22433_/A VGND VGND VPWR VPWR _22457_/X sky130_fd_sc_hd__buf_2
XANTENNA__16206__A _16222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _12687_/A _23788_/Q VGND VGND VPWR VPWR _12211_/C sky130_fd_sc_hd__or2_4
XANTENNA__15110__A _15103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21408_ _21297_/X _21405_/X _13933_/B _21402_/X VGND VGND VPWR VPWR _21408_/X sky130_fd_sc_hd__o22a_4
X_13190_ _11864_/A _13189_/X VGND VGND VPWR VPWR _13190_/X sky130_fd_sc_hd__and2_4
XFILLER_124_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22388_ _22141_/X _22383_/X _15533_/B _22387_/X VGND VGND VPWR VPWR _23297_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22282__B2 _22277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20293__B1 _20262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12141_ _12129_/A _12141_/B _12141_/C VGND VGND VPWR VPWR _12145_/B sky130_fd_sc_hd__and3_4
X_24127_ _24127_/CLK _22747_/X HRESETn VGND VGND VPWR VPWR _11511_/A sky130_fd_sc_hd__dfrtp_4
X_21339_ _21263_/X _21334_/X _12533_/B _21338_/X VGND VGND VPWR VPWR _23915_/D sky130_fd_sc_hd__o22a_4
XFILLER_2_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19517__A HRDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24186__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23039__A _18178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22034__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24058_ _24057_/CLK _21074_/X VGND VGND VPWR VPWR _14587_/B sky130_fd_sc_hd__dfxtp_4
X_12072_ _11990_/A _12136_/B VGND VGND VPWR VPWR _12073_/C sky130_fd_sc_hd__or2_4
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13565__A _13416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15900_ _13546_/A _15844_/B VGND VGND VPWR VPWR _15900_/X sky130_fd_sc_hd__or2_4
X_23009_ _22949_/A _23009_/B VGND VGND VPWR VPWR _23009_/X sky130_fd_sc_hd__or2_4
XFILLER_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22585__A2 _22558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17037__A _17048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16880_ _16860_/X _16862_/X _16878_/X _16880_/D VGND VGND VPWR VPWR _16880_/X sky130_fd_sc_hd__and4_4
XFILLER_103_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15831_ _12536_/A _15829_/X _15830_/X VGND VGND VPWR VPWR _15831_/X sky130_fd_sc_hd__and3_4
XFILLER_77_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15780__A _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18550_ _17762_/X _17724_/X _17762_/X _17724_/X VGND VGND VPWR VPWR _18550_/X sky130_fd_sc_hd__a2bb2o_4
X_12974_ _12974_/A _12902_/B VGND VGND VPWR VPWR _12974_/X sky130_fd_sc_hd__or2_4
X_15762_ _15741_/X _15762_/B VGND VGND VPWR VPWR _15764_/B sky130_fd_sc_hd__or2_4
XANTENNA__20398__A _20234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17501_ _17493_/A _17501_/B VGND VGND VPWR VPWR _17501_/X sky130_fd_sc_hd__or2_4
XFILLER_46_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14713_ _13596_/A _14713_/B VGND VGND VPWR VPWR _14713_/X sky130_fd_sc_hd__or2_4
X_18481_ _18111_/A _18366_/X _18478_/Y _18026_/X _18480_/X VGND VGND VPWR VPWR _18481_/X
+ sky130_fd_sc_hd__a32o_4
X_11925_ _16742_/A _23764_/Q VGND VGND VPWR VPWR _11926_/C sky130_fd_sc_hd__or2_4
X_15693_ _12726_/A _15689_/X _15692_/X VGND VGND VPWR VPWR _15693_/X sky130_fd_sc_hd__or3_4
XFILLER_46_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12909__A _12513_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11813__A _11813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17432_ _14261_/A _17441_/B VGND VGND VPWR VPWR _17432_/X sky130_fd_sc_hd__or2_4
X_11856_ _11856_/A VGND VGND VPWR VPWR _11857_/A sky130_fd_sc_hd__buf_2
XANTENNA__21006__B HRDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14644_ _14653_/A _14644_/B VGND VGND VPWR VPWR _14646_/B sky130_fd_sc_hd__or2_4
XPHY_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17363_ _17362_/X VGND VGND VPWR VPWR _17365_/A sky130_fd_sc_hd__inv_2
X_14575_ _13799_/A _14645_/B VGND VGND VPWR VPWR _14575_/X sky130_fd_sc_hd__or2_4
XANTENNA__15004__B _23541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11787_ _11742_/X VGND VGND VPWR VPWR _12122_/A sky130_fd_sc_hd__buf_2
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19102_ _19074_/X _19100_/X _19101_/Y _19079_/X VGND VGND VPWR VPWR _19102_/X sky130_fd_sc_hd__o22a_4
X_16314_ _13377_/A VGND VGND VPWR VPWR _16314_/X sky130_fd_sc_hd__buf_2
X_13526_ _13554_/A _23557_/Q VGND VGND VPWR VPWR _13526_/X sky130_fd_sc_hd__or2_4
X_17294_ _18651_/B _17294_/B VGND VGND VPWR VPWR _17294_/X sky130_fd_sc_hd__or2_4
XANTENNA__22118__A _22118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19033_ _19016_/X _19031_/X _19032_/Y _19021_/X VGND VGND VPWR VPWR _19033_/X sky130_fd_sc_hd__o22a_4
X_13457_ _13327_/A _13455_/X _13456_/X VGND VGND VPWR VPWR _13457_/X sky130_fd_sc_hd__and3_4
X_16245_ _16162_/X _16242_/X _16244_/Y VGND VGND VPWR VPWR _16246_/B sky130_fd_sc_hd__a21o_4
XANTENNA__16116__A _16116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12408_ _12363_/X _24108_/Q VGND VGND VPWR VPWR _12409_/C sky130_fd_sc_hd__or2_4
XFILLER_161_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21076__A2 _21073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13388_ _13408_/A _13388_/B VGND VGND VPWR VPWR _13391_/B sky130_fd_sc_hd__or2_4
X_16176_ _13398_/A VGND VGND VPWR VPWR _16210_/A sky130_fd_sc_hd__buf_2
XFILLER_154_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20861__A _20510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_20_0_HCLK clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_20_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15955__A _13462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12339_ _12338_/X VGND VGND VPWR VPWR _12339_/X sky130_fd_sc_hd__buf_2
XFILLER_126_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15127_ _14149_/A _15125_/X _15127_/C VGND VGND VPWR VPWR _15127_/X sky130_fd_sc_hd__and3_4
XFILLER_47_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19935_ _19931_/X _24172_/Q _19932_/X _21007_/B VGND VGND VPWR VPWR _24172_/D sky130_fd_sc_hd__o22a_4
X_15058_ _14074_/A _15058_/B _15057_/X VGND VGND VPWR VPWR _15058_/X sky130_fd_sc_hd__or3_4
XANTENNA__23223__CLK _23904_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22025__B2 _22021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19977__B1 _17653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14009_ _12501_/A _23872_/Q VGND VGND VPWR VPWR _14010_/C sky130_fd_sc_hd__or2_4
XANTENNA__13475__A _13475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19866_ _19865_/X VGND VGND VPWR VPWR _19866_/Y sky130_fd_sc_hd__inv_2
X_18817_ _18786_/A VGND VGND VPWR VPWR _18817_/X sky130_fd_sc_hd__buf_2
X_19797_ _19797_/A VGND VGND VPWR VPWR _19823_/B sky130_fd_sc_hd__inv_2
XFILLER_3_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16786__A _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15690__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18748_ _17982_/X VGND VGND VPWR VPWR _18748_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21000__A2 _20231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18679_ _17318_/A _18679_/B VGND VGND VPWR VPWR _18679_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12819__A _12833_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20710_ _20515_/X _20709_/X _24322_/Q _20522_/X VGND VGND VPWR VPWR _20711_/B sky130_fd_sc_hd__o22a_4
XANTENNA__11723__A _14658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21690_ _21575_/X _21684_/X _23712_/Q _21688_/X VGND VGND VPWR VPWR _21690_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20641_ _20778_/A VGND VGND VPWR VPWR _20641_/X sky130_fd_sc_hd__buf_2
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22500__A2 _22494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23360_ _23456_/CLK _23360_/D VGND VGND VPWR VPWR _23360_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20511__A1 _20418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20572_ _20438_/A _20572_/B VGND VGND VPWR VPWR _20572_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__20511__B2 _20510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22028__A _22007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22311_ _22151_/X _22308_/X _13876_/B _22305_/X VGND VGND VPWR VPWR _23357_/D sky130_fd_sc_hd__o22a_4
XFILLER_164_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23291_ _23772_/CLK _22396_/X VGND VGND VPWR VPWR _14495_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12554__A _12874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22242_ _22117_/X _22237_/X _12655_/B _22241_/X VGND VGND VPWR VPWR _22242_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21067__A2 _21066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21867__A _20841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22264__B2 _22262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12273__B _24076_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12752__A1 _11856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11555__A2 IRQ[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22173_ _21806_/A _22173_/B _22637_/C _20220_/A VGND VGND VPWR VPWR _22173_/X sky130_fd_sc_hd__or4_4
XFILLER_105_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22016__A1 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21124_ _20892_/X _21118_/X _24027_/Q _21122_/X VGND VGND VPWR VPWR _24027_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22016__B2 _22014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13385__A _13385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21055_ _20596_/X _21052_/X _24071_/Q _21049_/X VGND VGND VPWR VPWR _24071_/D sky130_fd_sc_hd__o22a_4
XFILLER_8_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21775__B1 _12672_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22698__A _22698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20006_ _20005_/X VGND VGND VPWR VPWR _20006_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17443__A1 _17162_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16696__A _16561_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_40_0_HCLK clkbuf_6_20_0_HCLK/X VGND VGND VPWR VPWR _23918_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22319__A2 _22315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21957_ _21957_/A VGND VGND VPWR VPWR _21957_/X sky130_fd_sc_hd__buf_2
XANTENNA__12729__A _12704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A VGND VGND VPWR VPWR _12372_/A sky130_fd_sc_hd__buf_2
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11633__A _11632_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20908_ _21017_/A _20908_/B VGND VGND VPWR VPWR _20908_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15105__A _15081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12690_ _12690_/A _23754_/Q VGND VGND VPWR VPWR _12690_/X sky130_fd_sc_hd__or2_4
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _21706_/A _21420_/B _21320_/C _20220_/A VGND VGND VPWR VPWR _21888_/X sky130_fd_sc_hd__or4_4
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23627_ _24074_/CLK _23627_/D VGND VGND VPWR VPWR _12646_/B sky130_fd_sc_hd__dfxtp_4
X_11641_ _20196_/A VGND VGND VPWR VPWR _11642_/A sky130_fd_sc_hd__buf_2
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _24221_/Q _20773_/X _20838_/X VGND VGND VPWR VPWR _20840_/A sky130_fd_sc_hd__o21a_4
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17320__A _21028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14367_/A _14360_/B VGND VGND VPWR VPWR _14360_/X sky130_fd_sc_hd__or2_4
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23558_ _23558_/CLK _23558_/D VGND VGND VPWR VPWR _13297_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20502__A1 _18210_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _20157_/A IRQ[17] _11571_/X VGND VGND VPWR VPWR _11572_/X sky130_fd_sc_hd__a21o_4
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13321_/A _13311_/B _13310_/X VGND VGND VPWR VPWR _13311_/X sky130_fd_sc_hd__and3_4
XFILLER_122_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22509_ _22437_/X _22508_/X _23241_/Q _22505_/X VGND VGND VPWR VPWR _22509_/X sky130_fd_sc_hd__o22a_4
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14291_ _11914_/A _14289_/X _14291_/C VGND VGND VPWR VPWR _14292_/C sky130_fd_sc_hd__and3_4
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23489_ _23649_/CLK _22072_/X VGND VGND VPWR VPWR _15566_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21058__A2 _21052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16030_ _16047_/A VGND VGND VPWR VPWR _16035_/A sky130_fd_sc_hd__buf_2
X_13242_ _12338_/X _13240_/X _13242_/C VGND VGND VPWR VPWR _13243_/C sky130_fd_sc_hd__and3_4
XANTENNA__21777__A _21770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23246__CLK _23246_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11546__A2 IRQ[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13173_ _12738_/A _13173_/B _13172_/X VGND VGND VPWR VPWR _13173_/X sky130_fd_sc_hd__and3_4
XFILLER_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12124_ _16608_/A _12124_/B VGND VGND VPWR VPWR _12124_/X sky130_fd_sc_hd__or2_4
X_17981_ _17980_/X VGND VGND VPWR VPWR _18288_/A sky130_fd_sc_hd__buf_2
XFILLER_46_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13295__A _13330_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19720_ _19571_/X _19704_/X _19718_/X _17811_/X _19719_/X VGND VGND VPWR VPWR _19720_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_78_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16932_ _16932_/A VGND VGND VPWR VPWR _16932_/X sky130_fd_sc_hd__buf_2
X_12055_ _11876_/X VGND VGND VPWR VPWR _16710_/A sky130_fd_sc_hd__buf_2
XFILLER_133_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20569__A1 _18299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19651_ _19589_/X _19596_/X VGND VGND VPWR VPWR _19651_/X sky130_fd_sc_hd__and2_4
XANTENNA__21230__A2 _21226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16863_ _15391_/D _13950_/X _15391_/D _13950_/X VGND VGND VPWR VPWR _16878_/A sky130_fd_sc_hd__a2bb2o_4
X_18602_ _17304_/X _18601_/Y VGND VGND VPWR VPWR _18602_/X sky130_fd_sc_hd__or2_4
X_15814_ _12876_/A _15869_/B VGND VGND VPWR VPWR _15814_/X sky130_fd_sc_hd__or2_4
X_19582_ _19578_/Y _19788_/A VGND VGND VPWR VPWR _19582_/X sky130_fd_sc_hd__and2_4
X_16794_ _16768_/A _16794_/B _16793_/X VGND VGND VPWR VPWR _16794_/X sky130_fd_sc_hd__or3_4
XFILLER_92_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18533_ _18533_/A _18533_/B VGND VGND VPWR VPWR _18533_/Y sky130_fd_sc_hd__nand2_4
XFILLER_92_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15745_ _12778_/X _15742_/X _15744_/X VGND VGND VPWR VPWR _15745_/X sky130_fd_sc_hd__and3_4
XFILLER_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12957_ _12957_/A _12957_/B _12957_/C VGND VGND VPWR VPWR _12957_/X sky130_fd_sc_hd__and3_4
XANTENNA__12639__A _12945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22730__A2 _22729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18464_ _18411_/A _18464_/B VGND VGND VPWR VPWR _18464_/X sky130_fd_sc_hd__and2_4
X_11908_ _16595_/A _11893_/X _11908_/C VGND VGND VPWR VPWR _11908_/X sky130_fd_sc_hd__and3_4
X_15676_ _12738_/A _15674_/X _15675_/X VGND VGND VPWR VPWR _15676_/X sky130_fd_sc_hd__and3_4
X_12888_ _12868_/A _24073_/Q VGND VGND VPWR VPWR _12889_/C sky130_fd_sc_hd__or2_4
XFILLER_33_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17415_ _22039_/B VGND VGND VPWR VPWR _17415_/Y sky130_fd_sc_hd__inv_2
X_14627_ _14684_/A _14627_/B VGND VGND VPWR VPWR _14628_/C sky130_fd_sc_hd__or2_4
X_11839_ _11760_/X VGND VGND VPWR VPWR _16768_/A sky130_fd_sc_hd__buf_2
X_18395_ _18330_/X _18372_/X _18373_/X _18394_/X VGND VGND VPWR VPWR _18395_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24021__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17346_ _16866_/X _17346_/B VGND VGND VPWR VPWR _17346_/Y sky130_fd_sc_hd__nor2_4
XFILLER_18_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14558_ _14280_/A _14556_/X _14558_/C VGND VGND VPWR VPWR _14559_/C sky130_fd_sc_hd__and3_4
XFILLER_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13509_ _13520_/A _13502_/X _13509_/C VGND VGND VPWR VPWR _13510_/C sky130_fd_sc_hd__or3_4
XANTENNA__12374__A _12373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17277_ _17273_/Y _17018_/X _17026_/X _17276_/X VGND VGND VPWR VPWR _17306_/A sky130_fd_sc_hd__o22a_4
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14489_ _14540_/A _14487_/X _14489_/C VGND VGND VPWR VPWR _14490_/C sky130_fd_sc_hd__and3_4
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19016_ _19016_/A VGND VGND VPWR VPWR _19016_/X sky130_fd_sc_hd__buf_2
X_16228_ _16220_/A _16226_/X _16227_/X VGND VGND VPWR VPWR _16228_/X sky130_fd_sc_hd__and3_4
XFILLER_146_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22246__B2 _22241_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24171__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15685__A _11970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16159_ _16159_/A _16159_/B _16159_/C VGND VGND VPWR VPWR _16159_/X sky130_fd_sc_hd__or3_4
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23739__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22549__A2 _22544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19918_ _19438_/A VGND VGND VPWR VPWR _22931_/A sky130_fd_sc_hd__buf_2
XFILLER_151_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19849_ _19849_/A _19849_/B _19849_/C VGND VGND VPWR VPWR _19849_/X sky130_fd_sc_hd__and3_4
XFILLER_25_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_27_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_27_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13933__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22860_ _17319_/Y _22848_/X _22849_/X VGND VGND VPWR VPWR _22860_/X sky130_fd_sc_hd__o21a_4
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21811_ _21526_/A VGND VGND VPWR VPWR _21811_/X sky130_fd_sc_hd__buf_2
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22791_ _22763_/Y _22792_/B VGND VGND VPWR VPWR _22791_/X sky130_fd_sc_hd__or2_4
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18925__A1 _17169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22721__A2 _22715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21742_ _21577_/X _21741_/X _23679_/Q _21738_/X VGND VGND VPWR VPWR _21742_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19620__A _19624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24461_ _23379_/CLK _18800_/X HRESETn VGND VGND VPWR VPWR _11575_/A sky130_fd_sc_hd__dfrtp_4
X_21673_ _21546_/X _21670_/X _23724_/Q _21667_/X VGND VGND VPWR VPWR _23724_/D sky130_fd_sc_hd__o22a_4
XFILLER_145_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14764__A _13853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17140__A _17139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23412_ _23476_/CLK _23412_/D VGND VGND VPWR VPWR _11827_/B sky130_fd_sc_hd__dfxtp_4
X_20624_ _20539_/X _20623_/X _24325_/Q _20549_/X VGND VGND VPWR VPWR _20624_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24392_ _24422_/CLK _24392_/D HRESETn VGND VGND VPWR VPWR _24392_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__23269__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22485__B2 _22421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23343_ _23918_/CLK _23343_/D VGND VGND VPWR VPWR _16266_/B sky130_fd_sc_hd__dfxtp_4
X_20555_ _24265_/Q _20443_/X _20554_/X VGND VGND VPWR VPWR _20555_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12284__A _13276_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23274_ _23531_/CLK _23274_/D VGND VGND VPWR VPWR _12759_/B sky130_fd_sc_hd__dfxtp_4
X_20486_ _20486_/A VGND VGND VPWR VPWR _20486_/X sky130_fd_sc_hd__buf_2
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22225_ _22258_/A VGND VGND VPWR VPWR _22226_/A sky130_fd_sc_hd__inv_2
XANTENNA__15595__A _15595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22156_ _22471_/A VGND VGND VPWR VPWR _22156_/X sky130_fd_sc_hd__buf_2
XANTENNA__21460__A2 _21455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_109_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR _23939_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21107_ _20596_/X _21104_/X _24039_/Q _21101_/X VGND VGND VPWR VPWR _21107_/X sky130_fd_sc_hd__o22a_4
XFILLER_160_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22087_ _21885_/X _22060_/A _23477_/Q _22042_/X VGND VGND VPWR VPWR _22087_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14004__A _12287_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21038_ _21045_/A VGND VGND VPWR VPWR _21038_/X sky130_fd_sc_hd__buf_2
XANTENNA__18613__B1 _18009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13860_ _14331_/A _13856_/X _13859_/X VGND VGND VPWR VPWR _13860_/X sky130_fd_sc_hd__or3_4
XFILLER_170_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12811_ _12773_/X _12809_/X _12810_/X VGND VGND VPWR VPWR _12811_/X sky130_fd_sc_hd__and3_4
XANTENNA__12459__A _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22989_ _23048_/A VGND VGND VPWR VPWR _22989_/X sky130_fd_sc_hd__buf_2
X_13791_ _13791_/A VGND VGND VPWR VPWR _15394_/A sky130_fd_sc_hd__buf_2
XANTENNA__18916__A1 _12980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15530_ _12258_/A _23777_/Q VGND VGND VPWR VPWR _15531_/C sky130_fd_sc_hd__or2_4
X_12742_ _13306_/A _12738_/X _12742_/C VGND VGND VPWR VPWR _12742_/X sky130_fd_sc_hd__or3_4
XFILLER_76_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12673_ _12975_/A _12671_/X _12673_/C VGND VGND VPWR VPWR _12673_/X sky130_fd_sc_hd__and3_4
X_15461_ _12578_/A _15456_/X _15460_/X VGND VGND VPWR VPWR _15461_/X sky130_fd_sc_hd__or3_4
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17160_/A _17196_/X _17119_/X _17199_/X VGND VGND VPWR VPWR _17200_/X sky130_fd_sc_hd__o22a_4
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _15517_/A _14412_/B _14412_/C VGND VGND VPWR VPWR _14412_/X sky130_fd_sc_hd__and3_4
X_11624_ _12213_/A VGND VGND VPWR VPWR _11886_/A sky130_fd_sc_hd__buf_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17050__A _17418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21279__A2 _21269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18180_ _17768_/X VGND VGND VPWR VPWR _18180_/X sky130_fd_sc_hd__buf_2
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _12530_/A _15454_/B VGND VGND VPWR VPWR _15392_/X sky130_fd_sc_hd__or2_4
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24194__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20487__B1 _24108_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ _17144_/A VGND VGND VPWR VPWR _17131_/X sky130_fd_sc_hd__buf_2
XFILLER_129_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11555_ _24460_/Q IRQ[23] _20182_/A VGND VGND VPWR VPWR _11555_/X sky130_fd_sc_hd__a21o_4
X_14343_ _14519_/A _14343_/B VGND VGND VPWR VPWR _14343_/X sky130_fd_sc_hd__or2_4
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12194__A _12194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24130__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17062_ _11644_/X _17077_/A _17078_/C _17062_/D VGND VGND VPWR VPWR _17062_/X sky130_fd_sc_hd__or4_4
X_14274_ _12454_/A _14345_/B VGND VGND VPWR VPWR _14275_/C sky130_fd_sc_hd__or2_4
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22228__B2 _22227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16013_ _11865_/X _16013_/B VGND VGND VPWR VPWR _16013_/X sky130_fd_sc_hd__and2_4
X_13225_ _13256_/A _23559_/Q VGND VGND VPWR VPWR _13226_/C sky130_fd_sc_hd__or2_4
XANTENNA__21300__A _21264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12922__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21987__B1 _23541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13156_ _13184_/A _13217_/B VGND VGND VPWR VPWR _13157_/C sky130_fd_sc_hd__or2_4
XANTENNA__21451__A2 _21448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12107_ _12001_/X _12107_/B _12107_/C VGND VGND VPWR VPWR _12107_/X sky130_fd_sc_hd__and3_4
XFILLER_151_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13087_ _13058_/A VGND VGND VPWR VPWR _13090_/A sky130_fd_sc_hd__buf_2
X_17964_ _17904_/X _17964_/B VGND VGND VPWR VPWR _17964_/X sky130_fd_sc_hd__and2_4
XANTENNA__19705__A _19705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19703_ _19703_/A HRDATA[7] VGND VGND VPWR VPWR _19703_/X sky130_fd_sc_hd__and2_4
XANTENNA__21203__A2 _21198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16915_ _16915_/A _17060_/B _16915_/C _16915_/D VGND VGND VPWR VPWR _16915_/X sky130_fd_sc_hd__or4_4
X_12038_ _16711_/A VGND VGND VPWR VPWR _16704_/A sky130_fd_sc_hd__buf_2
XANTENNA__22400__B2 _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17895_ _17783_/X _17894_/Y VGND VGND VPWR VPWR _17895_/X sky130_fd_sc_hd__and2_4
XANTENNA__14849__A _12188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20411__B1 _20714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19634_ _19781_/A _19614_/X _19634_/C _19633_/X VGND VGND VPWR VPWR _19634_/X sky130_fd_sc_hd__or4_4
X_16846_ _15919_/D _16845_/X _15919_/D _16845_/X VGND VGND VPWR VPWR _16846_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19565_ _19848_/A _19565_/B VGND VGND VPWR VPWR _19565_/X sky130_fd_sc_hd__or2_4
X_16777_ _16767_/A _16774_/X _16776_/X VGND VGND VPWR VPWR _16777_/X sky130_fd_sc_hd__and3_4
XFILLER_111_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13989_ _11931_/A _13989_/B _13989_/C VGND VGND VPWR VPWR _13989_/X sky130_fd_sc_hd__or3_4
XANTENNA__22703__A2 _22701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18516_ _17975_/X _18264_/Y _17870_/X _18515_/Y VGND VGND VPWR VPWR _18516_/X sky130_fd_sc_hd__a211o_4
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15728_ _13090_/A _15726_/X _15727_/X VGND VGND VPWR VPWR _15728_/X sky130_fd_sc_hd__and3_4
X_19496_ _19480_/X _19495_/X HRDATA[13] _19484_/X VGND VGND VPWR VPWR _19624_/A sky130_fd_sc_hd__o22a_4
XFILLER_33_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18447_ _17396_/D _18445_/X _18060_/X VGND VGND VPWR VPWR _18447_/Y sky130_fd_sc_hd__a21oi_4
X_15659_ _11881_/A _15659_/B _15658_/X VGND VGND VPWR VPWR _15659_/X sky130_fd_sc_hd__and3_4
XANTENNA__24289__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14584__A _12454_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15399__B _15399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18378_ _18378_/A _17496_/Y VGND VGND VPWR VPWR _18379_/D sky130_fd_sc_hd__and2_4
XANTENNA__22467__B2 _22457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17329_ _11935_/A _17297_/X _19863_/A _17039_/X VGND VGND VPWR VPWR _17329_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17343__B1 _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23561__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20340_ _20251_/X _20339_/X _20235_/X VGND VGND VPWR VPWR _20340_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__22219__A1 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21690__A2 _21684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22219__B2 _22184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13928__A _13928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20271_ _20270_/X VGND VGND VPWR VPWR _20490_/A sky130_fd_sc_hd__inv_2
XANTENNA__12832__A _13556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22010_ _22010_/A VGND VGND VPWR VPWR _22010_/X sky130_fd_sc_hd__buf_2
XANTENNA__21442__A2 _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13647__B _13738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12551__B _12655_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19615__A _19450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15121__A2 _17339_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23961_ _24057_/CLK _23961_/D VGND VGND VPWR VPWR _14737_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22041__A _22041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22912_ _20218_/A VGND VGND VPWR VPWR _22912_/X sky130_fd_sc_hd__buf_2
X_23892_ _23764_/CLK _23892_/D VGND VGND VPWR VPWR _23892_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22976__A _22975_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22843_ _20700_/A _17273_/Y VGND VGND VPWR VPWR _22843_/X sky130_fd_sc_hd__or2_4
XANTENNA__18769__A1_N _17015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12279__A _12279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22155__B1 _14363_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19350__A _19340_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22774_ _22773_/A _22773_/B VGND VGND VPWR VPWR _22778_/B sky130_fd_sc_hd__nand2_4
XFILLER_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21725_ _21548_/X _21720_/X _12500_/B _21724_/X VGND VGND VPWR VPWR _21725_/X sky130_fd_sc_hd__o22a_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20181__A2 IRQ[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21656_ _21806_/A _21656_/B _21706_/C _21236_/D VGND VGND VPWR VPWR _21656_/X sky130_fd_sc_hd__or4_4
X_24444_ _24445_/CLK _24444_/D HRESETn VGND VGND VPWR VPWR _24444_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23904__CLK _23904_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22458__B2 _22457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20607_ _18350_/X _20469_/X _20514_/X _20606_/Y VGND VGND VPWR VPWR _20607_/X sky130_fd_sc_hd__a211o_4
X_24375_ _24388_/CLK _24375_/D HRESETn VGND VGND VPWR VPWR _19120_/A sky130_fd_sc_hd__dfstp_4
X_21587_ _20892_/A VGND VGND VPWR VPWR _21587_/X sky130_fd_sc_hd__buf_2
XANTENNA__21130__B2 _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23326_ _23650_/CLK _22344_/X VGND VGND VPWR VPWR _23326_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_165_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20538_ _20233_/Y VGND VGND VPWR VPWR _20538_/X sky130_fd_sc_hd__buf_2
XFILLER_125_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23257_ _23194_/CLK _23257_/D VGND VGND VPWR VPWR _14774_/B sky130_fd_sc_hd__dfxtp_4
X_20469_ _20260_/A VGND VGND VPWR VPWR _20469_/X sky130_fd_sc_hd__buf_2
XFILLER_152_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13010_ _13010_/A _23592_/Q VGND VGND VPWR VPWR _13011_/C sky130_fd_sc_hd__or2_4
X_22208_ _22208_/A VGND VGND VPWR VPWR _22208_/X sky130_fd_sc_hd__buf_2
XANTENNA__21433__A2 _21427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22630__B2 _22626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23188_ _23475_/CLK _22592_/X VGND VGND VPWR VPWR _11793_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22139_ _20718_/A VGND VGND VPWR VPWR _22139_/X sky130_fd_sc_hd__buf_2
XFILLER_0_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14961_ _14976_/A _14961_/B VGND VGND VPWR VPWR _14961_/X sky130_fd_sc_hd__or2_4
XANTENNA__24354__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21197__B2 _21195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14669__A _14669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16700_ _16700_/A _24049_/Q VGND VGND VPWR VPWR _16702_/B sky130_fd_sc_hd__or2_4
XFILLER_130_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13912_ _11675_/A _13912_/B _13912_/C VGND VGND VPWR VPWR _13945_/B sky130_fd_sc_hd__or3_4
X_17680_ _16989_/A VGND VGND VPWR VPWR _17681_/A sky130_fd_sc_hd__buf_2
X_14892_ _14114_/A _14890_/X _14892_/C VGND VGND VPWR VPWR _14892_/X sky130_fd_sc_hd__and3_4
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16631_ _11786_/X VGND VGND VPWR VPWR _16786_/A sky130_fd_sc_hd__buf_2
Xclkbuf_6_10_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_10_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13843_ _15411_/A _13841_/X _13843_/C VGND VGND VPWR VPWR _13844_/C sky130_fd_sc_hd__and3_4
X_19350_ _19340_/A VGND VGND VPWR VPWR _19350_/X sky130_fd_sc_hd__buf_2
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16562_ _11960_/A _23954_/Q VGND VGND VPWR VPWR _16562_/X sky130_fd_sc_hd__or2_4
X_13774_ _13774_/A _13774_/B _13774_/C VGND VGND VPWR VPWR _13778_/B sky130_fd_sc_hd__and3_4
XANTENNA__22697__B2 _22691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18301_ _18301_/A _17773_/X _18180_/X VGND VGND VPWR VPWR _18302_/B sky130_fd_sc_hd__or3_4
X_15513_ _13051_/A _15511_/X _15512_/X VGND VGND VPWR VPWR _15513_/X sky130_fd_sc_hd__and3_4
XFILLER_43_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12725_ _12704_/A _12725_/B _12725_/C VGND VGND VPWR VPWR _12726_/C sky130_fd_sc_hd__and3_4
X_19281_ _19246_/B VGND VGND VPWR VPWR _19281_/Y sky130_fd_sc_hd__inv_2
X_16493_ _16479_/X _16424_/B VGND VGND VPWR VPWR _16495_/B sky130_fd_sc_hd__or2_4
XFILLER_30_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18232_ _17807_/X _18229_/Y _18089_/X _18231_/X VGND VGND VPWR VPWR _18232_/X sky130_fd_sc_hd__a211o_4
X_15444_ _15444_/A _15502_/B VGND VGND VPWR VPWR _15444_/X sky130_fd_sc_hd__or2_4
XANTENNA__24311__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12656_ _12610_/A VGND VGND VPWR VPWR _12943_/A sky130_fd_sc_hd__buf_2
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ _11607_/A VGND VGND VPWR VPWR _11608_/A sky130_fd_sc_hd__buf_2
X_18163_ _17975_/X _18157_/Y _18089_/X _18162_/Y VGND VGND VPWR VPWR _18163_/X sky130_fd_sc_hd__a211o_4
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12587_ _12587_/A VGND VGND VPWR VPWR _12670_/A sky130_fd_sc_hd__buf_2
X_15375_ _11697_/A _15373_/X _15375_/C VGND VGND VPWR VPWR _15375_/X sky130_fd_sc_hd__and3_4
XANTENNA__21121__B2 _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20853__B _20852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17114_ _12097_/X VGND VGND VPWR VPWR _17114_/X sky130_fd_sc_hd__buf_2
X_14326_ _13655_/A _14397_/B VGND VGND VPWR VPWR _14326_/X sky130_fd_sc_hd__or2_4
XANTENNA__21672__A2 _21670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11538_ _11538_/A _11538_/B VGND VGND VPWR VPWR _18995_/A sky130_fd_sc_hd__or2_4
X_18094_ _18538_/A VGND VGND VPWR VPWR _18095_/A sky130_fd_sc_hd__buf_2
XANTENNA__13748__A _12616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17045_ _17037_/Y _17040_/X _17297_/B VGND VGND VPWR VPWR _17046_/A sky130_fd_sc_hd__o21ai_4
X_14257_ _13882_/A _14253_/X _14256_/X VGND VGND VPWR VPWR _14258_/C sky130_fd_sc_hd__or3_4
XFILLER_48_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13208_ _13200_/X _13208_/B VGND VGND VPWR VPWR _13208_/X sky130_fd_sc_hd__or2_4
XFILLER_171_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14188_ _14199_/A _23359_/Q VGND VGND VPWR VPWR _14188_/X sky130_fd_sc_hd__or2_4
XFILLER_87_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22621__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13139_ _13139_/A _13208_/B VGND VGND VPWR VPWR _13139_/X sky130_fd_sc_hd__or2_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18996_ _18994_/Y _18995_/Y _11540_/B VGND VGND VPWR VPWR _18996_/X sky130_fd_sc_hd__o21a_4
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17947_ _17947_/A VGND VGND VPWR VPWR _17947_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14579__A _13593_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13483__A _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17878_ _17878_/A VGND VGND VPWR VPWR _17878_/X sky130_fd_sc_hd__buf_2
XANTENNA__14298__B _14362_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19617_ _24167_/Q _19457_/X HRDATA[19] _19454_/X VGND VGND VPWR VPWR _19617_/X sky130_fd_sc_hd__o22a_4
X_16829_ _16905_/B _16826_/X _16905_/B _16826_/X VGND VGND VPWR VPWR _16829_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16794__A _16768_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12099__A _12064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19548_ _19687_/C _19548_/B _19548_/C VGND VGND VPWR VPWR _19548_/X sky130_fd_sc_hd__and3_4
XFILLER_59_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21205__A _21198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19479_ _19479_/A VGND VGND VPWR VPWR _19504_/B sky130_fd_sc_hd__buf_2
XANTENNA__21360__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21510_ _21489_/A VGND VGND VPWR VPWR _21510_/X sky130_fd_sc_hd__buf_2
X_22490_ _22505_/A VGND VGND VPWR VPWR _22498_/A sky130_fd_sc_hd__buf_2
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21441_ _21441_/A VGND VGND VPWR VPWR _21441_/X sky130_fd_sc_hd__buf_2
XANTENNA__21112__B2 _21108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24160_ _24471_/CLK _24160_/D HRESETn VGND VGND VPWR VPWR _24160_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22860__A1 _17319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21372_ _21405_/A VGND VGND VPWR VPWR _21388_/A sky130_fd_sc_hd__inv_2
XFILLER_174_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15857__B _15796_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23111_ _23111_/CLK _23111_/D VGND VGND VPWR VPWR _23111_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13658__A _13658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20323_ _20270_/X VGND VGND VPWR VPWR _20323_/X sky130_fd_sc_hd__buf_2
X_24091_ _23592_/CLK _24091_/D VGND VGND VPWR VPWR _24091_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_162_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23042_ _23042_/A VGND VGND VPWR VPWR HADDR[23] sky130_fd_sc_hd__inv_2
X_20254_ _20253_/Y VGND VGND VPWR VPWR _20255_/A sky130_fd_sc_hd__buf_2
XANTENNA__21415__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21875__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20185_ _24462_/Q IRQ[25] _20184_/X VGND VGND VPWR VPWR _20185_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_77_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21179__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13393__A _13384_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22915__A2 _22930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11906__A _11905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23944_ _23592_/CLK _21272_/X VGND VGND VPWR VPWR _23944_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11625__B _11869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23875_ _23656_/CLK _21400_/X VGND VGND VPWR VPWR _15844_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14001__B _23232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22826_ _22819_/X _17327_/Y VGND VGND VPWR VPWR _22826_/X sky130_fd_sc_hd__or2_4
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17715__A2_N _17368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21115__A _21101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22757_ SYSTICKCLKDIV[0] _22749_/Y _22756_/X VGND VGND VPWR VPWR _22757_/X sky130_fd_sc_hd__a21bo_4
XANTENNA__12737__A _13304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21351__B2 _21345_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12510_ _12510_/A VGND VGND VPWR VPWR _12511_/A sky130_fd_sc_hd__buf_2
XFILLER_164_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15113__A _15091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13490_ _13532_/A _13420_/B VGND VGND VPWR VPWR _13490_/X sky130_fd_sc_hd__or2_4
X_21708_ _21741_/A VGND VGND VPWR VPWR _21724_/A sky130_fd_sc_hd__inv_2
X_22688_ _22687_/X VGND VGND VPWR VPWR _22722_/A sky130_fd_sc_hd__buf_2
X_12441_ _11910_/A VGND VGND VPWR VPWR _13955_/A sky130_fd_sc_hd__buf_2
X_21639_ _21572_/X _21634_/X _23745_/Q _21638_/X VGND VGND VPWR VPWR _23745_/D sky130_fd_sc_hd__o22a_4
X_24427_ _24428_/CLK _24427_/D HRESETn VGND VGND VPWR VPWR _24427_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21103__B2 _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19847__A2 _19687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12372_ _12372_/A VGND VGND VPWR VPWR _12948_/A sky130_fd_sc_hd__buf_2
X_15160_ _13791_/A _15158_/X _15159_/X VGND VGND VPWR VPWR _15160_/X sky130_fd_sc_hd__and3_4
XANTENNA__22851__A1 _17491_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24358_ _24398_/CLK _19039_/X HRESETn VGND VGND VPWR VPWR _24358_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21654__A2 _21620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_1_0_HCLK clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_1_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14111_ _15257_/A _23999_/Q VGND VGND VPWR VPWR _14111_/X sky130_fd_sc_hd__or2_4
X_23309_ _24045_/CLK _23309_/D VGND VGND VPWR VPWR _23309_/Q sky130_fd_sc_hd__dfxtp_4
X_15091_ _15091_/A _15087_/X _15090_/X VGND VGND VPWR VPWR _15091_/X sky130_fd_sc_hd__or3_4
XANTENNA__13568__A _13567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24289_ _24287_/CLK _19296_/X HRESETn VGND VGND VPWR VPWR _24289_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24232__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14042_ _14075_/A _23680_/Q VGND VGND VPWR VPWR _14042_/X sky130_fd_sc_hd__or2_4
XANTENNA__21406__A2 _21405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18807__B1 _24456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22603__B2 _22598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15783__A _12979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18850_ _18843_/A VGND VGND VPWR VPWR _18850_/X sky130_fd_sc_hd__buf_2
XFILLER_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20090__A1 _19402_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17801_ _18461_/A VGND VGND VPWR VPWR _17801_/X sky130_fd_sc_hd__buf_2
XFILLER_171_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18781_ _18780_/X _17060_/B _17091_/A _11598_/X VGND VGND VPWR VPWR _18837_/A sky130_fd_sc_hd__or4_4
X_15993_ _15993_/A _15993_/B _15993_/C VGND VGND VPWR VPWR _15994_/C sky130_fd_sc_hd__and3_4
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17732_ _17732_/A _17276_/X VGND VGND VPWR VPWR _17736_/A sky130_fd_sc_hd__or2_4
XANTENNA__11816__A _11815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14944_ _14925_/X _14942_/X _14943_/X VGND VGND VPWR VPWR _14944_/X sky130_fd_sc_hd__and3_4
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17663_ _17663_/A _17659_/X VGND VGND VPWR VPWR _17663_/X sky130_fd_sc_hd__or2_4
XANTENNA__15007__B _23925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22119__B1 _23467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14875_ _11895_/X _14875_/B VGND VGND VPWR VPWR _14875_/X sky130_fd_sc_hd__or2_4
XFILLER_169_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20393__A2 _20304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19402_ _19402_/A VGND VGND VPWR VPWR _19402_/X sky130_fd_sc_hd__buf_2
X_16614_ _11792_/X VGND VGND VPWR VPWR _16654_/A sky130_fd_sc_hd__buf_2
XFILLER_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13826_ _14329_/A _13901_/B VGND VGND VPWR VPWR _13826_/X sky130_fd_sc_hd__or2_4
X_17594_ _17108_/X VGND VGND VPWR VPWR _17594_/X sky130_fd_sc_hd__buf_2
XFILLER_91_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14846__B _14845_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19333_ _19957_/A VGND VGND VPWR VPWR _23083_/D sky130_fd_sc_hd__buf_2
X_16545_ _12001_/X _16543_/X _16545_/C VGND VGND VPWR VPWR _16550_/B sky130_fd_sc_hd__and3_4
X_13757_ _14541_/A _13757_/B VGND VGND VPWR VPWR _13757_/X sky130_fd_sc_hd__or2_4
XFILLER_90_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21342__B2 _21338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15023__A _15000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12708_ _12708_/A _12708_/B _12708_/C VGND VGND VPWR VPWR _12708_/X sky130_fd_sc_hd__or3_4
X_19264_ _24305_/Q _19254_/B _19263_/Y VGND VGND VPWR VPWR _24305_/D sky130_fd_sc_hd__o21a_4
X_16476_ _16166_/X _16476_/B VGND VGND VPWR VPWR _16476_/X sky130_fd_sc_hd__or2_4
X_13688_ _15449_/A _13684_/X _13687_/X VGND VGND VPWR VPWR _13688_/X sky130_fd_sc_hd__or3_4
XFILLER_15_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18215_ _18019_/X VGND VGND VPWR VPWR _18215_/X sky130_fd_sc_hd__buf_2
XANTENNA__15958__A _13431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15427_ _15408_/A _15427_/B _15427_/C VGND VGND VPWR VPWR _15427_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_17_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR _24271_/CLK sky130_fd_sc_hd__clkbuf_1
X_12639_ _12945_/A _12633_/X _12639_/C VGND VGND VPWR VPWR _12640_/C sky130_fd_sc_hd__or3_4
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19195_ _19144_/X VGND VGND VPWR VPWR _19195_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14862__A _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18334__A _18406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18146_ _16992_/B VGND VGND VPWR VPWR _18148_/C sky130_fd_sc_hd__inv_2
X_15358_ _15326_/A _23384_/Q VGND VGND VPWR VPWR _15360_/B sky130_fd_sc_hd__or2_4
XFILLER_145_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13478__A _12869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14309_ _12470_/A _14309_/B _14309_/C VGND VGND VPWR VPWR _14310_/C sky130_fd_sc_hd__and3_4
X_18077_ _18335_/A _17571_/A VGND VGND VPWR VPWR _18079_/C sky130_fd_sc_hd__and2_4
X_15289_ _14277_/A _15289_/B _15288_/X VGND VGND VPWR VPWR _15289_/X sky130_fd_sc_hd__or3_4
XFILLER_144_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21695__A _21674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17028_ _17027_/X VGND VGND VPWR VPWR _17028_/X sky130_fd_sc_hd__buf_2
XANTENNA__15693__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22070__A2 _22067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20104__A _20124_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18979_ _18959_/X _18977_/X _18978_/X _24368_/Q VGND VGND VPWR VPWR _24368_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21990_ _21990_/A VGND VGND VPWR VPWR _21991_/A sky130_fd_sc_hd__buf_2
XFILLER_152_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14102__A _14138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20941_ _21007_/A _20380_/B VGND VGND VPWR VPWR _20941_/X sky130_fd_sc_hd__or2_4
XANTENNA__21581__B2 _21573_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13941__A _13697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23660_ _24012_/CLK _21773_/X VGND VGND VPWR VPWR _23660_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20872_ _20664_/A _20871_/X _20671_/A VGND VGND VPWR VPWR _20873_/A sky130_fd_sc_hd__o21ai_4
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22611_ _22442_/X _22608_/X _13216_/B _22605_/X VGND VGND VPWR VPWR _22611_/X sky130_fd_sc_hd__o22a_4
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23591_ _23723_/CLK _21912_/X VGND VGND VPWR VPWR _23591_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19361__A1_N _19358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12557__A _12515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16029__A _16056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21333__B2 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22530__B1 _14600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22542_ _22536_/Y _22541_/X _22410_/X _22541_/X VGND VGND VPWR VPWR _23220_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21884__A2 _21875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15868__A _13543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22473_ _22158_/A VGND VGND VPWR VPWR _22473_/X sky130_fd_sc_hd__buf_2
XANTENNA__14772__A _14772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18244__A _17900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24255__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21424_ _21431_/A VGND VGND VPWR VPWR _21424_/X sky130_fd_sc_hd__buf_2
X_24212_ _24184_/CLK _24212_/D HRESETn VGND VGND VPWR VPWR _24212_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21636__A2 _21634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22833__A1 _17353_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13388__A _13408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24143_ _24134_/CLK _20074_/Y HRESETn VGND VGND VPWR VPWR _24143_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21355_ _21322_/A VGND VGND VPWR VPWR _21355_/X sky130_fd_sc_hd__buf_2
XANTENNA__12292__A _13183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20306_ _20234_/X VGND VGND VPWR VPWR _20306_/X sky130_fd_sc_hd__buf_2
X_24074_ _24074_/CLK _21051_/X VGND VGND VPWR VPWR _24074_/Q sky130_fd_sc_hd__dfxtp_4
X_21286_ _21285_/X _21281_/X _15470_/B _21276_/X VGND VGND VPWR VPWR _23938_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23025_ _23043_/A _18216_/X VGND VGND VPWR VPWR _23025_/Y sky130_fd_sc_hd__nand2_4
XFILLER_115_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20237_ _20237_/A VGND VGND VPWR VPWR _20864_/A sky130_fd_sc_hd__buf_2
XANTENNA__22061__A2 _22060_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20168_ IRQ[7] VGND VGND VPWR VPWR _20168_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18017__A1 _16935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12990_ _12862_/A _12990_/B _12990_/C VGND VGND VPWR VPWR _12990_/X sky130_fd_sc_hd__and3_4
X_20099_ _20124_/B _20099_/B _20098_/X _20196_/A VGND VGND VPWR VPWR _20099_/X sky130_fd_sc_hd__or4_4
XFILLER_40_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14012__A _14012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23927_ _23192_/CLK _23927_/D VGND VGND VPWR VPWR _15146_/B sky130_fd_sc_hd__dfxtp_4
X_11941_ _11941_/A _23796_/Q VGND VGND VPWR VPWR _11942_/C sky130_fd_sc_hd__or2_4
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17776__B1 _17768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13851__A _11933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14660_ _14660_/A _14660_/B _14660_/C VGND VGND VPWR VPWR _14660_/X sky130_fd_sc_hd__or3_4
X_11872_ _11872_/A VGND VGND VPWR VPWR _12857_/A sky130_fd_sc_hd__buf_2
X_23858_ _23852_/CLK _23858_/D VGND VGND VPWR VPWR _23858_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13611_ _14292_/A _13602_/X _13610_/X VGND VGND VPWR VPWR _13611_/X sky130_fd_sc_hd__or3_4
X_22809_ _14767_/Y _22804_/X VGND VGND VPWR VPWR HWDATA[4] sky130_fd_sc_hd__nor2_4
X_14591_ _15393_/A _14591_/B VGND VGND VPWR VPWR _14591_/X sky130_fd_sc_hd__or2_4
X_23789_ _24045_/CLK _21545_/X VGND VGND VPWR VPWR _16178_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12467__A _12467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22521__B1 _23232_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22883__B _22882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16330_ _16318_/A _16271_/B VGND VGND VPWR VPWR _16330_/X sky130_fd_sc_hd__or2_4
XFILLER_125_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13542_ _13542_/A _13539_/X _13541_/X VGND VGND VPWR VPWR _13542_/X sky130_fd_sc_hd__and3_4
XFILLER_125_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16261_ _15936_/X _16259_/X _16260_/X VGND VGND VPWR VPWR _16261_/X sky130_fd_sc_hd__and3_4
XANTENNA__15778__A _15778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13473_ _13443_/A _23653_/Q VGND VGND VPWR VPWR _13474_/C sky130_fd_sc_hd__or2_4
XFILLER_51_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14682__A _14682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18000_ _17975_/X _17979_/Y _17870_/X _17999_/Y VGND VGND VPWR VPWR _18000_/X sky130_fd_sc_hd__a211o_4
X_15212_ _14616_/A _15210_/X _15212_/C VGND VGND VPWR VPWR _15212_/X sky130_fd_sc_hd__and3_4
X_12424_ _12466_/A VGND VGND VPWR VPWR _12425_/A sky130_fd_sc_hd__buf_2
X_16192_ _16192_/A VGND VGND VPWR VPWR _16202_/A sky130_fd_sc_hd__buf_2
XANTENNA__22824__A1 _13692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15143_ _13799_/A _15143_/B VGND VGND VPWR VPWR _15144_/C sky130_fd_sc_hd__or2_4
X_12355_ _12596_/A VGND VGND VPWR VPWR _13258_/A sky130_fd_sc_hd__buf_2
XFILLER_153_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19951_ _19950_/X VGND VGND VPWR VPWR _19951_/X sky130_fd_sc_hd__buf_2
X_12286_ _11930_/A VGND VGND VPWR VPWR _12287_/A sky130_fd_sc_hd__buf_2
X_15074_ _15091_/A _15069_/X _15073_/X VGND VGND VPWR VPWR _15074_/X sky130_fd_sc_hd__or3_4
XFILLER_141_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18902_ _12180_/X _18897_/X _24403_/Q _18900_/X VGND VGND VPWR VPWR _24403_/D sky130_fd_sc_hd__o22a_4
X_14025_ _13888_/A _23200_/Q VGND VGND VPWR VPWR _14025_/X sky130_fd_sc_hd__or2_4
XANTENNA__22052__A2 _22046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12930__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19882_ _19607_/X _19881_/X _22039_/B _19700_/X VGND VGND VPWR VPWR _19882_/X sky130_fd_sc_hd__o22a_4
XFILLER_136_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18833_ _12061_/A _12097_/X _12028_/X _12078_/X VGND VGND VPWR VPWR _18834_/D sky130_fd_sc_hd__or4_4
XFILLER_171_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18764_ _12024_/A _19963_/B VGND VGND VPWR VPWR _19965_/B sky130_fd_sc_hd__nor2_4
XANTENNA__15018__A _15018_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15976_ _15959_/A _23470_/Q VGND VGND VPWR VPWR _15977_/C sky130_fd_sc_hd__or2_4
XFILLER_49_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20859__A _20859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17715_ _16982_/A _17368_/X _16982_/A _17368_/X VGND VGND VPWR VPWR _17715_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24128__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14927_ _14973_/A _14859_/B VGND VGND VPWR VPWR _14927_/X sky130_fd_sc_hd__or2_4
XFILLER_76_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18695_ _18694_/X VGND VGND VPWR VPWR _18695_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14857__A _12218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13761__A _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17646_ _17250_/X _18768_/A _17594_/X _17645_/X VGND VGND VPWR VPWR _17647_/B sky130_fd_sc_hd__o22a_4
X_14858_ _14094_/A _14856_/X _14858_/C VGND VGND VPWR VPWR _14863_/B sky130_fd_sc_hd__and3_4
X_13809_ _12445_/A _13809_/B _13809_/C VGND VGND VPWR VPWR _13813_/B sky130_fd_sc_hd__and3_4
X_17577_ _17574_/Y _17024_/A _17031_/A _17576_/Y VGND VGND VPWR VPWR _18114_/B sky130_fd_sc_hd__o22a_4
X_14789_ _15081_/A _14787_/X _14789_/C VGND VGND VPWR VPWR _14789_/X sky130_fd_sc_hd__and3_4
XFILLER_90_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19316_ _19228_/A _19227_/X _19315_/Y VGND VGND VPWR VPWR _24279_/D sky130_fd_sc_hd__o21a_4
XANTENNA__24278__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16528_ _16528_/A _16527_/X VGND VGND VPWR VPWR _16528_/X sky130_fd_sc_hd__or2_4
XFILLER_149_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21866__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15688__A _12721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19247_ _19247_/A _19247_/B VGND VGND VPWR VPWR _19248_/B sky130_fd_sc_hd__and2_4
X_16459_ _11727_/A VGND VGND VPWR VPWR _16491_/A sky130_fd_sc_hd__buf_2
XANTENNA__14592__A _15394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21079__B1 _24053_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21618__A2 _21613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19178_ _19153_/A _19153_/B _19177_/Y VGND VGND VPWR VPWR _19178_/X sky130_fd_sc_hd__o21a_4
XFILLER_157_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18129_ _17848_/A _18123_/X _18125_/X _17809_/A _18128_/X VGND VGND VPWR VPWR _18130_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18495__B2 _18494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13308__A1 _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13001__A _12881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21140_ _21136_/A VGND VGND VPWR VPWR _21155_/A sky130_fd_sc_hd__buf_2
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21071_ _20860_/X _21066_/X _24060_/Q _21070_/X VGND VGND VPWR VPWR _21071_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13936__A _14390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20022_ _19956_/A VGND VGND VPWR VPWR _20022_/X sky130_fd_sc_hd__buf_2
XFILLER_154_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24485__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20769__A _22459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20357__A2 _20340_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0_0_HCLK_A clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21973_ _21860_/X _21967_/X _23552_/Q _21971_/X VGND VGND VPWR VPWR _21973_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14767__A _14766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13671__A _12191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23712_ _23649_/CLK _21690_/X VGND VGND VPWR VPWR _23712_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20924_ _20924_/A _20730_/B VGND VGND VPWR VPWR _20924_/X sky130_fd_sc_hd__or2_4
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23643_ _23675_/CLK _21797_/X VGND VGND VPWR VPWR _14470_/B sky130_fd_sc_hd__dfxtp_4
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20855_ _24252_/Q VGND VGND VPWR VPWR _20855_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21306__A1 _21304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12287__A _12287_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21306__B2 _21300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23574_ _23511_/CLK _23574_/D VGND VGND VPWR VPWR _14934_/B sky130_fd_sc_hd__dfxtp_4
X_20786_ _20676_/X _20783_/Y _20785_/X _19078_/Y _20731_/X VGND VGND VPWR VPWR _20787_/A
+ sky130_fd_sc_hd__a32o_4
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22525_ _22466_/X _22522_/X _13848_/B _22519_/X VGND VGND VPWR VPWR _22525_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22456_ _20744_/A VGND VGND VPWR VPWR _22456_/X sky130_fd_sc_hd__buf_2
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_63_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR _23558_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15110__B _15033_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21407_ _21295_/X _21405_/X _13769_/B _21402_/X VGND VGND VPWR VPWR _21407_/X sky130_fd_sc_hd__o22a_4
X_22387_ _22358_/A VGND VGND VPWR VPWR _22387_/X sky130_fd_sc_hd__buf_2
XANTENNA__22282__A2 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14007__A _12467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12140_ _12164_/A _24019_/Q VGND VGND VPWR VPWR _12141_/C sky130_fd_sc_hd__or2_4
XANTENNA__21490__B1 _12565_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21338_ _21338_/A VGND VGND VPWR VPWR _21338_/X sky130_fd_sc_hd__buf_2
X_24126_ _24127_/CLK _24126_/D HRESETn VGND VGND VPWR VPWR _22910_/B sky130_fd_sc_hd__dfstp_4
XFILLER_123_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12071_ _12102_/A _12135_/B VGND VGND VPWR VPWR _12073_/B sky130_fd_sc_hd__or2_4
X_21269_ _21269_/A VGND VGND VPWR VPWR _21269_/X sky130_fd_sc_hd__buf_2
XANTENNA__19435__B1 _19399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22034__A2 _22031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24057_ _24057_/CLK _24057_/D VGND VGND VPWR VPWR _24057_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16222__A _16222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12750__A _11864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23008_ _22912_/X VGND VGND VPWR VPWR _23008_/X sky130_fd_sc_hd__buf_2
XFILLER_103_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21793__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15830_ _12864_/A _15830_/B VGND VGND VPWR VPWR _15830_/X sky130_fd_sc_hd__or2_4
XANTENNA__24155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23055__A _18062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15761_ _13099_/A _15759_/X _15761_/C VGND VGND VPWR VPWR _15761_/X sky130_fd_sc_hd__and3_4
X_12973_ _12973_/A _23241_/Q VGND VGND VPWR VPWR _12975_/B sky130_fd_sc_hd__or2_4
XFILLER_17_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14677__A _14677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21545__B2 _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17500_ _16768_/A _17378_/X _17379_/X VGND VGND VPWR VPWR _17501_/B sky130_fd_sc_hd__o21a_4
XFILLER_166_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14712_ _13589_/A _14708_/X _14711_/X VGND VGND VPWR VPWR _14712_/X sky130_fd_sc_hd__or3_4
X_18480_ _24143_/Q _18479_/Y _16981_/X VGND VGND VPWR VPWR _18480_/X sky130_fd_sc_hd__o21a_4
X_11924_ _11905_/X VGND VGND VPWR VPWR _16742_/A sky130_fd_sc_hd__buf_2
X_15692_ _13170_/A _15690_/X _15692_/C VGND VGND VPWR VPWR _15692_/X sky130_fd_sc_hd__and3_4
XFILLER_46_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17431_ _17429_/B VGND VGND VPWR VPWR _17441_/B sky130_fd_sc_hd__inv_2
XFILLER_79_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14643_ _13882_/A VGND VGND VPWR VPWR _15625_/A sky130_fd_sc_hd__buf_2
X_11855_ _11855_/A VGND VGND VPWR VPWR _11856_/A sky130_fd_sc_hd__buf_2
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12197__A _15444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17362_ _15653_/X _17445_/B VGND VGND VPWR VPWR _17362_/X sky130_fd_sc_hd__or2_4
XPHY_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14574_ _14574_/A _14644_/B VGND VGND VPWR VPWR _14574_/X sky130_fd_sc_hd__or2_4
XFILLER_82_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11786_ _16222_/A VGND VGND VPWR VPWR _11786_/X sky130_fd_sc_hd__buf_2
XANTENNA__18174__B1 _18168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19101_ _19101_/A VGND VGND VPWR VPWR _19101_/Y sky130_fd_sc_hd__inv_2
X_16313_ _16313_/A _16313_/B _16313_/C VGND VGND VPWR VPWR _16320_/B sky130_fd_sc_hd__and3_4
X_13525_ _13515_/X _22337_/A VGND VGND VPWR VPWR _13525_/X sky130_fd_sc_hd__or2_4
X_17293_ _17292_/X VGND VGND VPWR VPWR _17294_/B sky130_fd_sc_hd__inv_2
XANTENNA__12925__A _12925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17921__B1 _17820_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19032_ _19032_/A VGND VGND VPWR VPWR _19032_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15301__A _14296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16244_ _16243_/X VGND VGND VPWR VPWR _16244_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13456_ _13427_/A _23973_/Q VGND VGND VPWR VPWR _13456_/X sky130_fd_sc_hd__or2_4
XANTENNA__12644__B _23979_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12407_ _12407_/A _12293_/B VGND VGND VPWR VPWR _12407_/X sky130_fd_sc_hd__or2_4
XANTENNA__15020__B _24053_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16175_ _16205_/A _16168_/X _16175_/C VGND VGND VPWR VPWR _16187_/B sky130_fd_sc_hd__or3_4
XFILLER_12_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13387_ _13387_/A VGND VGND VPWR VPWR _13408_/A sky130_fd_sc_hd__buf_2
XFILLER_115_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15126_ _14148_/A _23735_/Q VGND VGND VPWR VPWR _15127_/C sky130_fd_sc_hd__or2_4
X_12338_ _12401_/A VGND VGND VPWR VPWR _12338_/X sky130_fd_sc_hd__buf_2
XFILLER_138_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22134__A _20658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19934_ _19931_/X _24173_/Q _19932_/X _20422_/B VGND VGND VPWR VPWR _19934_/X sky130_fd_sc_hd__o22a_4
X_15057_ _14073_/A _15054_/X _15057_/C VGND VGND VPWR VPWR _15057_/X sky130_fd_sc_hd__and3_4
XANTENNA__22025__A2 _22024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12660__A _12962_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12269_ _12269_/A VGND VGND VPWR VPWR _12690_/A sky130_fd_sc_hd__buf_2
XANTENNA__19977__A1 _16935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14008_ _12188_/A _23712_/Q VGND VGND VPWR VPWR _14008_/X sky130_fd_sc_hd__or2_4
XFILLER_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19865_ _19700_/A _19859_/X _19862_/Y _21184_/C _19552_/X VGND VGND VPWR VPWR _19865_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15971__A _15971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18816_ _15651_/X _18810_/X _24449_/Q _18811_/X VGND VGND VPWR VPWR _24449_/D sky130_fd_sc_hd__o22a_4
X_19796_ _19528_/B _19795_/X _19691_/Y VGND VGND VPWR VPWR _19803_/C sky130_fd_sc_hd__o21a_4
XFILLER_62_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15959_ _15959_/A VGND VGND VPWR VPWR _15960_/A sky130_fd_sc_hd__buf_2
X_18747_ _17815_/X _18746_/X _17820_/X _17818_/X VGND VGND VPWR VPWR _18747_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__14587__A _13601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22733__B1 _15176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13491__A _13542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18678_ _18538_/X _17350_/B _17594_/X _17630_/B VGND VGND VPWR VPWR _18679_/B sky130_fd_sc_hd__o22a_4
XFILLER_97_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17629_ _18693_/B _17628_/X _17326_/B VGND VGND VPWR VPWR _17630_/B sky130_fd_sc_hd__o21a_4
XFILLER_145_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20640_ _16899_/A _20244_/B VGND VGND VPWR VPWR _20778_/A sky130_fd_sc_hd__and2_4
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20571_ _20466_/X _20562_/Y _20569_/X _20570_/Y _20481_/X VGND VGND VPWR VPWR _20572_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12835__A _13349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16307__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22310_ _22149_/X _22308_/X _13605_/B _22305_/X VGND VGND VPWR VPWR _22310_/X sky130_fd_sc_hd__o22a_4
X_23290_ _23290_/CLK _22398_/X VGND VGND VPWR VPWR _14564_/B sky130_fd_sc_hd__dfxtp_4
X_22241_ _22226_/A VGND VGND VPWR VPWR _22241_/X sky130_fd_sc_hd__buf_2
XANTENNA__22264__A2 _22258_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22172_ _21133_/A VGND VGND VPWR VPWR _22637_/C sky130_fd_sc_hd__buf_2
XFILLER_172_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21123_ _20860_/X _21118_/X _24028_/Q _21122_/X VGND VGND VPWR VPWR _21123_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22016__A2 _22010_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13666__A _13666_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12570__A _12570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16042__A _16049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21054_ _20575_/X _21052_/X _24072_/Q _21049_/X VGND VGND VPWR VPWR _24072_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21883__A _21313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21775__B2 _21774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20005_ _19992_/X _17660_/A _19998_/X _20004_/X VGND VGND VPWR VPWR _20005_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17443__A2 _17421_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_HCLK clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21527__B2 _21525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22724__B1 _13765_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21956_ _21831_/X _21953_/X _12376_/B _21950_/X VGND VGND VPWR VPWR _21956_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _20754_/X _20906_/X _19135_/A _20761_/X VGND VGND VPWR VPWR _20908_/B sky130_fd_sc_hd__o22a_4
XFILLER_36_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ _23604_/Q VGND VGND VPWR VPWR _21887_/Y sky130_fd_sc_hd__inv_2
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _23467_/CLK _21837_/X VGND VGND VPWR VPWR _12723_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _19957_/A _11640_/B VGND VGND VPWR VPWR _20196_/A sky130_fd_sc_hd__or2_4
XFILLER_70_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _20935_/A _20837_/X VGND VGND VPWR VPWR _20838_/X sky130_fd_sc_hd__or2_4
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23557_ _23557_/CLK _21966_/X VGND VGND VPWR VPWR _23557_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _24453_/Q IRQ[16] VGND VGND VPWR VPWR _11571_/X sky130_fd_sc_hd__and2_4
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16217__A _16163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20769_ _22459_/A VGND VGND VPWR VPWR _20770_/A sky130_fd_sc_hd__buf_2
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _13313_/A _23974_/Q VGND VGND VPWR VPWR _13310_/X sky130_fd_sc_hd__or2_4
XFILLER_161_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22508_ _22508_/A VGND VGND VPWR VPWR _22508_/X sky130_fd_sc_hd__buf_2
XFILLER_167_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14290_ _12504_/A _23548_/Q VGND VGND VPWR VPWR _14291_/C sky130_fd_sc_hd__or2_4
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23488_ _24096_/CLK _22073_/X VGND VGND VPWR VPWR _23488_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12464__B _23787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ _13253_/A _13241_/B VGND VGND VPWR VPWR _13242_/C sky130_fd_sc_hd__or2_4
X_22439_ _22437_/X _22438_/X _12915_/B _22433_/X VGND VGND VPWR VPWR _23273_/D sky130_fd_sc_hd__o22a_4
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14960__A _11697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13172_ _13304_/A _13241_/B VGND VGND VPWR VPWR _13172_/X sky130_fd_sc_hd__or2_4
XANTENNA__15775__B _15702_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24109_ _24077_/CLK _20465_/X VGND VGND VPWR VPWR _24109_/Q sky130_fd_sc_hd__dfxtp_4
X_12123_ _11694_/X _12123_/B _12123_/C VGND VGND VPWR VPWR _12123_/X sky130_fd_sc_hd__or3_4
XANTENNA__17048__A _17048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17682__A2 _17455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17980_ _17249_/X VGND VGND VPWR VPWR _17980_/X sky130_fd_sc_hd__buf_2
XANTENNA__12480__A _12867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24336__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21215__B1 _15487_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16931_ _16931_/A _17297_/A VGND VGND VPWR VPWR _16932_/A sky130_fd_sc_hd__and2_4
X_12054_ _16592_/A _12054_/B _12054_/C VGND VGND VPWR VPWR _12054_/X sky130_fd_sc_hd__or3_4
XFILLER_104_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21766__B2 _21760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15791__A _12741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19650_ _19578_/Y _19643_/A VGND VGND VPWR VPWR _19655_/B sky130_fd_sc_hd__and2_4
X_16862_ _15391_/A _16861_/X _15391_/A _16861_/X VGND VGND VPWR VPWR _16862_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20974__C1 _20973_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15813_ _12875_/A _15868_/B VGND VGND VPWR VPWR _15815_/B sky130_fd_sc_hd__or2_4
XFILLER_120_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18601_ _17301_/A _18600_/X _17289_/X VGND VGND VPWR VPWR _18601_/Y sky130_fd_sc_hd__a21boi_4
X_19581_ _19581_/A VGND VGND VPWR VPWR _19788_/A sky130_fd_sc_hd__buf_2
X_16793_ _16767_/A _16791_/X _16792_/X VGND VGND VPWR VPWR _16793_/X sky130_fd_sc_hd__and3_4
XFILLER_19_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21518__B2 _21482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18532_ _18453_/X _18530_/X _24480_/Q _18531_/X VGND VGND VPWR VPWR _18532_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15744_ _15743_/X _15744_/B VGND VGND VPWR VPWR _15744_/X sky130_fd_sc_hd__or2_4
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12956_ _12949_/A _23849_/Q VGND VGND VPWR VPWR _12957_/C sky130_fd_sc_hd__or2_4
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18463_ _18462_/X VGND VGND VPWR VPWR _18463_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11907_ _11941_/A _23540_/Q VGND VGND VPWR VPWR _11908_/C sky130_fd_sc_hd__or2_4
X_15675_ _13145_/A _15675_/B VGND VGND VPWR VPWR _15675_/X sky130_fd_sc_hd__or2_4
XFILLER_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12887_ _12867_/A _23625_/Q VGND VGND VPWR VPWR _12889_/B sky130_fd_sc_hd__or2_4
XANTENNA__18607__A _18483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17414_ _17414_/A VGND VGND VPWR VPWR _22039_/B sky130_fd_sc_hd__buf_2
XFILLER_21_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14626_ _14669_/A VGND VGND VPWR VPWR _14684_/A sky130_fd_sc_hd__buf_2
X_11838_ _12169_/A _11838_/B _11838_/C VGND VGND VPWR VPWR _11849_/B sky130_fd_sc_hd__or3_4
XFILLER_57_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18394_ _18375_/X _18380_/Y _18390_/X _18392_/Y _18393_/X VGND VGND VPWR VPWR _18394_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22129__A _20612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21033__A _21033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17345_ _15047_/Y _17025_/A _17025_/Y _17751_/B VGND VGND VPWR VPWR _17346_/B sky130_fd_sc_hd__o22a_4
XFILLER_92_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14557_ _14270_/A _14627_/B VGND VGND VPWR VPWR _14558_/C sky130_fd_sc_hd__or2_4
XANTENNA__12655__A _12942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11769_ _11768_/X VGND VGND VPWR VPWR _11832_/A sky130_fd_sc_hd__buf_2
XFILLER_159_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15031__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13508_ _13503_/X _13505_/X _13507_/X VGND VGND VPWR VPWR _13509_/C sky130_fd_sc_hd__and3_4
X_17276_ _17276_/A _17275_/X VGND VGND VPWR VPWR _17276_/X sky130_fd_sc_hd__or2_4
XFILLER_146_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14488_ _14378_/A _14488_/B VGND VGND VPWR VPWR _14489_/C sky130_fd_sc_hd__or2_4
XFILLER_146_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24316__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19015_ _19010_/X _19014_/X _19010_/X _11536_/A VGND VGND VPWR VPWR _24362_/D sky130_fd_sc_hd__a2bb2o_4
X_16227_ _16219_/A _23885_/Q VGND VGND VPWR VPWR _16227_/X sky130_fd_sc_hd__or2_4
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13439_ _12873_/A VGND VGND VPWR VPWR _13467_/A sky130_fd_sc_hd__buf_2
XANTENNA__22246__A2 _22244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19438__A _19438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14870__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16158_ _16123_/A _16158_/B _16158_/C VGND VGND VPWR VPWR _16159_/C sky130_fd_sc_hd__and3_4
XFILLER_114_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13486__A _12659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15109_ _15081_/A _15107_/X _15108_/X VGND VGND VPWR VPWR _15113_/B sky130_fd_sc_hd__and3_4
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16089_ _16086_/X _16089_/B VGND VGND VPWR VPWR _16246_/A sky130_fd_sc_hd__or2_4
XANTENNA__23340__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19917_ _19906_/X _21007_/A _22904_/D VGND VGND VPWR VPWR _24180_/D sky130_fd_sc_hd__o21ai_4
XFILLER_87_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16797__A _16635_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19848_ _19848_/A _19848_/B VGND VGND VPWR VPWR _19849_/C sky130_fd_sc_hd__or2_4
XFILLER_56_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19779_ _19777_/Y _19811_/B _19675_/A VGND VGND VPWR VPWR _19779_/X sky130_fd_sc_hd__o21a_4
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22706__B1 _12564_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21509__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21810_ _21809_/X VGND VGND VPWR VPWR _21810_/X sky130_fd_sc_hd__buf_2
XANTENNA__15206__A _14677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22790_ _22792_/B _22789_/Y _22790_/C VGND VGND VPWR VPWR _24123_/D sky130_fd_sc_hd__and3_4
XFILLER_37_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14110__A _14110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12549__B _12549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22182__B2 _22177_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21741_ _21741_/A VGND VGND VPWR VPWR _21741_/X sky130_fd_sc_hd__buf_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17421__A _14084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24460_ _23379_/CLK _18801_/X HRESETn VGND VGND VPWR VPWR _24460_/Q sky130_fd_sc_hd__dfrtp_4
X_21672_ _21544_/X _21670_/X _16226_/B _21667_/X VGND VGND VPWR VPWR _21672_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_4_13_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_26_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23411_ _23475_/CLK _23411_/D VGND VGND VPWR VPWR _12158_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20623_ _20540_/X _20622_/X _24357_/Q _20547_/X VGND VGND VPWR VPWR _20623_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12565__A _12513_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24391_ _24422_/CLK _24391_/D HRESETn VGND VGND VPWR VPWR _19032_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__22485__A2 _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16037__A _16187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23342_ _24078_/CLK _23342_/D VGND VGND VPWR VPWR _16048_/B sky130_fd_sc_hd__dfxtp_4
X_20554_ _20398_/X _20536_/X _20537_/X _20553_/Y VGND VGND VPWR VPWR _20554_/X sky130_fd_sc_hd__a211o_4
XFILLER_20_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17361__A1 _17353_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17361__B2 _17360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14175__A1 _13951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15876__A _13546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23273_ _23241_/CLK _23273_/D VGND VGND VPWR VPWR _12915_/B sky130_fd_sc_hd__dfxtp_4
X_20485_ _20485_/A VGND VGND VPWR VPWR _20486_/A sky130_fd_sc_hd__buf_2
X_22224_ _22223_/X VGND VGND VPWR VPWR _22258_/A sky130_fd_sc_hd__buf_2
XFILLER_69_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13396__A _13408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11909__A _12466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22155_ _22153_/X _22147_/X _14363_/B _22154_/X VGND VGND VPWR VPWR _22155_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18861__A1 _13262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21106_ _20575_/X _21104_/X _24040_/Q _21101_/X VGND VGND VPWR VPWR _24040_/D sky130_fd_sc_hd__o22a_4
XFILLER_133_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22086_ _21883_/X _22081_/X _23478_/Q _22042_/X VGND VGND VPWR VPWR _23478_/D sky130_fd_sc_hd__o22a_4
X_21037_ _21033_/A VGND VGND VPWR VPWR _21045_/A sky130_fd_sc_hd__buf_2
XANTENNA__18613__A1 _17890_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21118__A _21118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20022__A _19956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12810_ _12775_/A _23978_/Q VGND VGND VPWR VPWR _12810_/X sky130_fd_sc_hd__or2_4
XANTENNA__15116__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19811__A _19811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13790_ _13954_/A VGND VGND VPWR VPWR _13791_/A sky130_fd_sc_hd__buf_2
XANTENNA__14020__A _13696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22988_ _22987_/X VGND VGND VPWR VPWR HADDR[14] sky130_fd_sc_hd__inv_2
XFILLER_55_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12741_ _12741_/A _12739_/X _12741_/C VGND VGND VPWR VPWR _12742_/C sky130_fd_sc_hd__and3_4
XFILLER_15_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_0_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21939_ _21706_/A _22173_/B _21706_/C _20220_/A VGND VGND VPWR VPWR _21939_/X sky130_fd_sc_hd__or4_4
X_15460_ _12587_/A _15458_/X _15460_/C VGND VGND VPWR VPWR _15460_/X sky130_fd_sc_hd__and3_4
X_12672_ _12974_/A _12672_/B VGND VGND VPWR VPWR _12673_/C sky130_fd_sc_hd__or2_4
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14674__B _14590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _11813_/A _14395_/X _14410_/X VGND VGND VPWR VPWR _14412_/C sky130_fd_sc_hd__or3_4
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _23294_/CLK _23609_/D VGND VGND VPWR VPWR _14739_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A VGND VGND VPWR VPWR _12213_/A sky130_fd_sc_hd__buf_2
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15391_ _15391_/A _13950_/X _15391_/C _15391_/D VGND VGND VPWR VPWR _15391_/X sky130_fd_sc_hd__or4_4
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19877__B1 _19811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22891__B _22891_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20487__A1 _20418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _17160_/A VGND VGND VPWR VPWR _17130_/X sky130_fd_sc_hd__buf_2
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20487__B2 _20396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _13916_/A VGND VGND VPWR VPWR _14519_/A sky130_fd_sc_hd__buf_2
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11554_ _11554_/A IRQ[22] VGND VGND VPWR VPWR _20182_/A sky130_fd_sc_hd__and2_4
XFILLER_168_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20692__A _20692_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24377__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17352__A1 _17272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17061_ _17060_/X VGND VGND VPWR VPWR _17077_/A sky130_fd_sc_hd__buf_2
XANTENNA__15786__A _15783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14273_ _14304_/A _14343_/B VGND VGND VPWR VPWR _14275_/B sky130_fd_sc_hd__or2_4
XANTENNA__14690__A _15616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24489__CLK _24294_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16012_ _15934_/X _16012_/B _16012_/C VGND VGND VPWR VPWR _16013_/B sky130_fd_sc_hd__or3_4
XFILLER_7_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13224_ _13248_/A _13148_/B VGND VGND VPWR VPWR _13224_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_33_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_3_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21987__B2 _21950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11819__A _11762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13155_ _13183_/A _13216_/B VGND VGND VPWR VPWR _13157_/B sky130_fd_sc_hd__or2_4
XANTENNA__18852__A1 _17139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12106_ _12106_/A _23891_/Q VGND VGND VPWR VPWR _12107_/C sky130_fd_sc_hd__or2_4
X_13086_ _13103_/A _13086_/B _13086_/C VGND VGND VPWR VPWR _13091_/B sky130_fd_sc_hd__and3_4
X_17963_ _16941_/X VGND VGND VPWR VPWR _17963_/X sky130_fd_sc_hd__buf_2
XANTENNA__19705__B _19705_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22412__A _20336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21739__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19702_ HRDATA[23] VGND VGND VPWR VPWR _20844_/A sky130_fd_sc_hd__buf_2
X_16914_ _16914_/A VGND VGND VPWR VPWR _16915_/D sky130_fd_sc_hd__inv_2
XANTENNA__18604__A1 _17980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17506__A _17172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12037_ _16713_/A VGND VGND VPWR VPWR _16695_/A sky130_fd_sc_hd__buf_2
XANTENNA__22400__A2 _22397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17894_ _17655_/X VGND VGND VPWR VPWR _17894_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19633_ _19510_/X _19632_/X VGND VGND VPWR VPWR _19633_/X sky130_fd_sc_hd__and2_4
XANTENNA__21028__A _21028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16845_ _15920_/X _16842_/X _15925_/Y VGND VGND VPWR VPWR _16845_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19721__A HRDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19564_ _19521_/Y _19899_/B _19563_/X VGND VGND VPWR VPWR _19565_/B sky130_fd_sc_hd__o21a_4
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16776_ _16811_/A _16776_/B VGND VGND VPWR VPWR _16776_/X sky130_fd_sc_hd__or2_4
X_13988_ _12468_/A _13988_/B _13987_/X VGND VGND VPWR VPWR _13989_/C sky130_fd_sc_hd__and3_4
XFILLER_168_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22164__B2 _22154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15727_ _12762_/A _23780_/Q VGND VGND VPWR VPWR _15727_/X sky130_fd_sc_hd__or2_4
X_18515_ _18288_/A _18266_/X VGND VGND VPWR VPWR _18515_/Y sky130_fd_sc_hd__nor2_4
X_12939_ _12951_/A _23689_/Q VGND VGND VPWR VPWR _12939_/X sky130_fd_sc_hd__or2_4
XFILLER_20_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19495_ _24177_/Q _19481_/X HRDATA[29] _19482_/X VGND VGND VPWR VPWR _19495_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21911__A1 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18337__A _18283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21911__B2 _21906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15658_ _12687_/A _15658_/B VGND VGND VPWR VPWR _15658_/X sky130_fd_sc_hd__or2_4
X_18446_ _17396_/D _18445_/X VGND VGND VPWR VPWR _18446_/X sky130_fd_sc_hd__or2_4
X_14609_ _15415_/A _14607_/X _14609_/C VGND VGND VPWR VPWR _14610_/C sky130_fd_sc_hd__and3_4
XFILLER_159_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18377_ _18377_/A _17497_/X VGND VGND VPWR VPWR _18379_/C sky130_fd_sc_hd__nor2_4
XFILLER_105_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15589_ _15611_/A _23745_/Q VGND VGND VPWR VPWR _15590_/C sky130_fd_sc_hd__or2_4
XFILLER_14_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21675__B1 _12664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_115_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR _23646_/CLK sky130_fd_sc_hd__clkbuf_1
X_17328_ _21133_/A VGND VGND VPWR VPWR _19863_/A sky130_fd_sc_hd__inv_2
XANTENNA__23706__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21698__A _21658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22219__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17259_ _17256_/X _17259_/B VGND VGND VPWR VPWR _17260_/A sky130_fd_sc_hd__or2_4
XANTENNA__24258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20270_ _18889_/B _19948_/X VGND VGND VPWR VPWR _20270_/X sky130_fd_sc_hd__or2_4
XFILLER_115_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14105__A _11898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13944__A _11813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23960_ _23290_/CLK _21229_/X VGND VGND VPWR VPWR _23960_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16320__A _13407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22911_ _22910_/X VGND VGND VPWR VPWR _22930_/A sky130_fd_sc_hd__buf_2
XFILLER_99_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23891_ _23764_/CLK _21378_/X VGND VGND VPWR VPWR _23891_/Q sky130_fd_sc_hd__dfxtp_4
X_22842_ _22845_/A _22842_/B VGND VGND VPWR VPWR HWDATA[14] sky130_fd_sc_hd__nor2_4
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22155__B2 _22154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22773_ _22773_/A _22773_/B VGND VGND VPWR VPWR _22777_/A sky130_fd_sc_hd__or2_4
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21724_ _21724_/A VGND VGND VPWR VPWR _21724_/X sky130_fd_sc_hd__buf_2
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24443_ _24445_/CLK _24443_/D HRESETn VGND VGND VPWR VPWR _24443_/Q sky130_fd_sc_hd__dfrtp_4
X_21655_ _21655_/A VGND VGND VPWR VPWR _21655_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20606_ _20652_/A _20605_/X VGND VGND VPWR VPWR _20606_/Y sky130_fd_sc_hd__nor2_4
X_24374_ _24419_/CLK _24374_/D HRESETn VGND VGND VPWR VPWR _20990_/A sky130_fd_sc_hd__dfstp_4
X_21586_ _21584_/X _21578_/X _23772_/Q _21585_/X VGND VGND VPWR VPWR _21586_/X sky130_fd_sc_hd__o22a_4
XFILLER_165_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21130__A2 _21125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23325_ _23679_/CLK _23325_/D VGND VGND VPWR VPWR _13818_/B sky130_fd_sc_hd__dfxtp_4
X_20537_ _20253_/Y VGND VGND VPWR VPWR _20537_/X sky130_fd_sc_hd__buf_2
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13838__B _13838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20468_ _20251_/A _20467_/X _20306_/X VGND VGND VPWR VPWR _20468_/Y sky130_fd_sc_hd__o21ai_4
X_23256_ _23194_/CLK _23256_/D VGND VGND VPWR VPWR _15253_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_152_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21969__B2 _21964_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22207_ _22144_/X _22201_/X _23424_/Q _22205_/X VGND VGND VPWR VPWR _23424_/D sky130_fd_sc_hd__o22a_4
XFILLER_165_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20399_ _20307_/X _20776_/A _20308_/X VGND VGND VPWR VPWR _20399_/X sky130_fd_sc_hd__a21o_4
XANTENNA__22630__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23187_ _23475_/CLK _23187_/D VGND VGND VPWR VPWR _12135_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22138_ _22137_/X _22135_/X _15869_/B _22130_/X VGND VGND VPWR VPWR _22138_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14960_ _11697_/A _14958_/X _14959_/X VGND VGND VPWR VPWR _14960_/X sky130_fd_sc_hd__and3_4
X_22069_ _21853_/X _22067_/X _15833_/B _22064_/X VGND VGND VPWR VPWR _22069_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21197__A2 _21191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13911_ _13928_/A _13903_/X _13911_/C VGND VGND VPWR VPWR _13912_/C sky130_fd_sc_hd__and3_4
X_14891_ _14110_/A _14891_/B VGND VGND VPWR VPWR _14892_/C sky130_fd_sc_hd__or2_4
XFILLER_43_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16630_ _16683_/A _16619_/X _16629_/X VGND VGND VPWR VPWR _16630_/X sky130_fd_sc_hd__and3_4
X_13842_ _12198_/A _13842_/B VGND VGND VPWR VPWR _13843_/C sky130_fd_sc_hd__or2_4
XFILLER_47_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20687__A _20686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16561_ _16561_/A _16561_/B _16561_/C VGND VGND VPWR VPWR _16561_/X sky130_fd_sc_hd__or3_4
X_13773_ _12927_/A _24094_/Q VGND VGND VPWR VPWR _13774_/C sky130_fd_sc_hd__or2_4
XANTENNA__22697__A2 _22694_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15512_ _12626_/A _15512_/B VGND VGND VPWR VPWR _15512_/X sky130_fd_sc_hd__or2_4
X_18300_ _18187_/X _18278_/X _18219_/X _18299_/X VGND VGND VPWR VPWR _18300_/X sky130_fd_sc_hd__o22a_4
X_12724_ _13279_/A _24074_/Q VGND VGND VPWR VPWR _12725_/C sky130_fd_sc_hd__or2_4
X_19280_ _19246_/A _19246_/B _19279_/Y VGND VGND VPWR VPWR _24297_/D sky130_fd_sc_hd__o21a_4
X_16492_ _16474_/A _16490_/X _16492_/C VGND VGND VPWR VPWR _16492_/X sky130_fd_sc_hd__and3_4
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18770__B1 _17100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18231_ _18562_/A _18230_/Y VGND VGND VPWR VPWR _18231_/X sky130_fd_sc_hd__and2_4
X_15443_ _12190_/A _15501_/B VGND VGND VPWR VPWR _15445_/B sky130_fd_sc_hd__or2_4
X_12655_ _12942_/A _12655_/B VGND VGND VPWR VPWR _12655_/X sky130_fd_sc_hd__or2_4
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ _11606_/A VGND VGND VPWR VPWR _11607_/A sky130_fd_sc_hd__buf_2
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18162_ _18288_/A _18161_/X VGND VGND VPWR VPWR _18162_/Y sky130_fd_sc_hd__nor2_4
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _12580_/A _23640_/Q VGND VGND VPWR VPWR _15375_/C sky130_fd_sc_hd__or2_4
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12586_ _12634_/A VGND VGND VPWR VPWR _12587_/A sky130_fd_sc_hd__buf_2
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22407__A _22462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17113_ _12093_/X VGND VGND VPWR VPWR _17113_/X sky130_fd_sc_hd__buf_2
XFILLER_157_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21311__A _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _14325_/A _14396_/B VGND VGND VPWR VPWR _14327_/B sky130_fd_sc_hd__or2_4
XFILLER_102_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11537_ _19004_/A _11537_/B VGND VGND VPWR VPWR _11538_/B sky130_fd_sc_hd__or2_4
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18093_ _17807_/X _18637_/B _18089_/X _18092_/X VGND VGND VPWR VPWR _18093_/X sky130_fd_sc_hd__a211o_4
XFILLER_157_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17044_ _17357_/B _17044_/B VGND VGND VPWR VPWR _17297_/B sky130_fd_sc_hd__or2_4
X_14256_ _15595_/A _14254_/X _14256_/C VGND VGND VPWR VPWR _14256_/X sky130_fd_sc_hd__and3_4
XANTENNA__12652__B _12549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13207_ _13220_/A _24039_/Q VGND VGND VPWR VPWR _13207_/X sky130_fd_sc_hd__or2_4
X_14187_ _14229_/A VGND VGND VPWR VPWR _14199_/A sky130_fd_sc_hd__buf_2
XFILLER_135_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13138_ _13300_/A _24039_/Q VGND VGND VPWR VPWR _13140_/B sky130_fd_sc_hd__or2_4
XFILLER_140_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18995_ _18995_/A VGND VGND VPWR VPWR _18995_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22142__A _22118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13764__A _12616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13069_ _13055_/A VGND VGND VPWR VPWR _13085_/A sky130_fd_sc_hd__buf_2
X_17946_ _17922_/X _17852_/X _17945_/X _17234_/X VGND VGND VPWR VPWR _17947_/A sky130_fd_sc_hd__o22a_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22385__B2 _22380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21981__A _21941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17877_ _17876_/X VGND VGND VPWR VPWR _17877_/X sky130_fd_sc_hd__buf_2
X_19616_ _19615_/X VGND VGND VPWR VPWR _19690_/B sky130_fd_sc_hd__buf_2
X_16828_ _16905_/A _16827_/X _16905_/A _16827_/X VGND VGND VPWR VPWR _16828_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19547_ _19816_/B _19546_/X VGND VGND VPWR VPWR _19548_/C sky130_fd_sc_hd__or2_4
X_16759_ _16759_/A _16756_/X _16759_/C VGND VGND VPWR VPWR _16759_/X sky130_fd_sc_hd__and3_4
XANTENNA__14595__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19478_ _19446_/A _19477_/X HRDATA[15] _19461_/X VGND VGND VPWR VPWR _19479_/A sky130_fd_sc_hd__o22a_4
XFILLER_22_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21360__A2 _21355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18429_ _17767_/A _18428_/X _17767_/A _18428_/X VGND VGND VPWR VPWR _18429_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15203__B _15146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13004__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21440_ _21266_/X _21434_/X _12817_/B _21438_/X VGND VGND VPWR VPWR _23850_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21112__A2 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21371_ _21370_/X VGND VGND VPWR VPWR _21405_/A sky130_fd_sc_hd__buf_2
XFILLER_163_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16315__A _11714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12843__A _12753_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24360__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23110_ _24102_/CLK _23110_/D VGND VGND VPWR VPWR _23110_/Q sky130_fd_sc_hd__dfxtp_4
X_20322_ _20321_/X VGND VGND VPWR VPWR _20322_/Y sky130_fd_sc_hd__inv_2
X_24090_ _24090_/CLK _20916_/X VGND VGND VPWR VPWR _14598_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_163_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19608__A3 _19606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20253_ _20229_/X VGND VGND VPWR VPWR _20253_/Y sky130_fd_sc_hd__inv_2
X_23041_ _23036_/X _17675_/A _23019_/X _23040_/X VGND VGND VPWR VPWR _23042_/A sky130_fd_sc_hd__a211o_4
XANTENNA__18816__A1 _15651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20184_ _11575_/X _20183_/Y VGND VGND VPWR VPWR _20184_/X sky130_fd_sc_hd__or2_4
XFILLER_135_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21179__A2 _21176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21891__A _21906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23943_ _23111_/CLK _23943_/D VGND VGND VPWR VPWR _23943_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24184__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23874_ _23650_/CLK _23874_/D VGND VGND VPWR VPWR _15505_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_57_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11625__C _12299_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22128__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22825_ _22814_/X _22825_/B VGND VGND VPWR VPWR HWDATA[9] sky130_fd_sc_hd__nor2_4
XFILLER_53_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22756_ _22755_/Y _24121_/Q SYSTICKCLKDIV[2] _22753_/Y VGND VGND VPWR VPWR _22756_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_71_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21351__A2 _21348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21707_ _21706_/X VGND VGND VPWR VPWR _21741_/A sky130_fd_sc_hd__buf_2
XFILLER_73_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22687_ _22687_/A _22687_/B _22637_/C _22637_/D VGND VGND VPWR VPWR _22687_/X sky130_fd_sc_hd__or4_4
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12440_ _12440_/A _12437_/X _12439_/X VGND VGND VPWR VPWR _12440_/X sky130_fd_sc_hd__and3_4
XFILLER_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24426_ _24422_/CLK _24426_/D HRESETn VGND VGND VPWR VPWR _24426_/Q sky130_fd_sc_hd__dfrtp_4
X_21638_ _21624_/A VGND VGND VPWR VPWR _21638_/X sky130_fd_sc_hd__buf_2
XANTENNA__21103__A2 _21097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14952__B _23958_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22227__A _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22300__B2 _22298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13849__A _13676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12371_ _12387_/A _12369_/X _12370_/X VGND VGND VPWR VPWR _12371_/X sky130_fd_sc_hd__and3_4
X_24357_ _24357_/CLK _19045_/X HRESETn VGND VGND VPWR VPWR _24357_/Q sky130_fd_sc_hd__dfstp_4
X_21569_ _21568_/X _21566_/X _15797_/B _21561_/X VGND VGND VPWR VPWR _21569_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12753__A _12752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14110_ _14110_/A VGND VGND VPWR VPWR _15257_/A sky130_fd_sc_hd__buf_2
XFILLER_154_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23308_ _23852_/CLK _22372_/X VGND VGND VPWR VPWR _12223_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20862__B2 _20861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15090_ _15112_/A _15090_/B _15090_/C VGND VGND VPWR VPWR _15090_/X sky130_fd_sc_hd__and3_4
X_24288_ _24292_/CLK _24288_/D HRESETn VGND VGND VPWR VPWR _19237_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_109_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14041_ _11753_/A _14037_/X _14041_/C VGND VGND VPWR VPWR _14041_/X sky130_fd_sc_hd__or3_4
X_23239_ _24039_/CLK _22511_/X VGND VGND VPWR VPWR _13179_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18807__A1 _13266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22603__A2 _22601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23401__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17800_ _18440_/A VGND VGND VPWR VPWR _18461_/A sky130_fd_sc_hd__buf_2
XANTENNA__17056__A _17015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15992_ _15960_/A _23438_/Q VGND VGND VPWR VPWR _15993_/C sky130_fd_sc_hd__or2_4
X_18780_ _18779_/X VGND VGND VPWR VPWR _18780_/X sky130_fd_sc_hd__buf_2
XANTENNA__22367__B2 _22366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17731_ _17727_/A _17399_/X _17727_/X VGND VGND VPWR VPWR _17731_/X sky130_fd_sc_hd__a21bo_4
X_14943_ _14967_/A _23990_/Q VGND VGND VPWR VPWR _14943_/X sky130_fd_sc_hd__or2_4
XFILLER_85_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17662_ _17659_/X _17661_/X VGND VGND VPWR VPWR _17779_/B sky130_fd_sc_hd__nor2_4
X_14874_ _14905_/A _23158_/Q VGND VGND VPWR VPWR _14874_/X sky130_fd_sc_hd__or2_4
XANTENNA__22119__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19401_ _11511_/A VGND VGND VPWR VPWR _19402_/A sky130_fd_sc_hd__buf_2
XFILLER_63_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16613_ _11762_/X VGND VGND VPWR VPWR _16656_/A sky130_fd_sc_hd__buf_2
X_13825_ _13666_/A _13900_/B VGND VGND VPWR VPWR _13825_/X sky130_fd_sc_hd__or2_4
XFILLER_165_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17593_ _17132_/Y _17256_/B _17260_/Y _17592_/X VGND VGND VPWR VPWR _18768_/A sky130_fd_sc_hd__o22a_4
XFILLER_63_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16544_ _12106_/A _23794_/Q VGND VGND VPWR VPWR _16545_/C sky130_fd_sc_hd__or2_4
X_19332_ _19325_/X _19331_/X _24276_/Q _19325_/X VGND VGND VPWR VPWR _24276_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15304__A _14169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13756_ _13756_/A _13756_/B _13756_/C VGND VGND VPWR VPWR _13764_/B sky130_fd_sc_hd__or3_4
XFILLER_91_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21342__A2 _21341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12647__B _12647_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12707_ _12298_/A _12707_/B _12707_/C VGND VGND VPWR VPWR _12708_/C sky130_fd_sc_hd__and3_4
XANTENNA__11551__B IRQ[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16475_ _16164_/X _16415_/B VGND VGND VPWR VPWR _16475_/X sky130_fd_sc_hd__or2_4
X_19263_ _19255_/B VGND VGND VPWR VPWR _19263_/Y sky130_fd_sc_hd__inv_2
X_13687_ _13687_/A _13687_/B _13686_/X VGND VGND VPWR VPWR _13687_/X sky130_fd_sc_hd__and3_4
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15426_ _14319_/A _15490_/B VGND VGND VPWR VPWR _15427_/C sky130_fd_sc_hd__or2_4
XFILLER_19_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18214_ _18145_/X _18213_/X _20023_/A _18145_/X VGND VGND VPWR VPWR _24491_/D sky130_fd_sc_hd__a2bb2o_4
X_12638_ _12944_/A _12638_/B _12637_/X VGND VGND VPWR VPWR _12639_/C sky130_fd_sc_hd__and3_4
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19194_ _24324_/Q _19144_/X _19193_/Y VGND VGND VPWR VPWR _19194_/X sky130_fd_sc_hd__o21a_4
XFILLER_19_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22137__A _20692_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18145_ _17900_/A VGND VGND VPWR VPWR _18145_/X sky130_fd_sc_hd__buf_2
X_15357_ _11654_/A _15357_/B _15357_/C VGND VGND VPWR VPWR _15361_/B sky130_fd_sc_hd__and3_4
XFILLER_102_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ _12569_/A _12665_/B VGND VGND VPWR VPWR _12569_/X sky130_fd_sc_hd__or2_4
XFILLER_145_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14308_ _12485_/A _24060_/Q VGND VGND VPWR VPWR _14309_/C sky130_fd_sc_hd__or2_4
XFILLER_102_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18076_ _18222_/A _18076_/B VGND VGND VPWR VPWR _18079_/B sky130_fd_sc_hd__and2_4
X_15288_ _15269_/A _15286_/X _15288_/C VGND VGND VPWR VPWR _15288_/X sky130_fd_sc_hd__and3_4
XFILLER_172_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17027_ _17026_/X VGND VGND VPWR VPWR _17027_/X sky130_fd_sc_hd__buf_2
XANTENNA__15974__A _16011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14239_ _14623_/A _23391_/Q VGND VGND VPWR VPWR _14239_/X sky130_fd_sc_hd__or2_4
XFILLER_131_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20081__A2 _20079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18978_ _18959_/A VGND VGND VPWR VPWR _18978_/X sky130_fd_sc_hd__buf_2
XFILLER_26_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20104__B _20093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17929_ _18126_/A _17927_/X _17850_/X _17928_/X VGND VGND VPWR VPWR _17930_/A sky130_fd_sc_hd__o22a_4
XFILLER_61_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14102__B _23775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20940_ _20940_/A _20561_/B VGND VGND VPWR VPWR _20940_/X sky130_fd_sc_hd__or2_4
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21581__A2 _21578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21216__A _21202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20871_ _20871_/A _20867_/A VGND VGND VPWR VPWR _20871_/X sky130_fd_sc_hd__and2_4
XANTENNA__12838__A _13367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22610_ _22440_/X _22608_/X _13012_/B _22605_/X VGND VGND VPWR VPWR _23176_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11742__A _16056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15214__A _14669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23590_ _23723_/CLK _23590_/D VGND VGND VPWR VPWR _13365_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__A1 _13192_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6_0_HCLK_A clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21333__A2 _21327_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22530__B2 _22526_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22541_ _22548_/A VGND VGND VPWR VPWR _22541_/X sky130_fd_sc_hd__buf_2
XANTENNA__24273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15868__B _15868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22472_ _22471_/X _22462_/X _14484_/B _22469_/X VGND VGND VPWR VPWR _22472_/X sky130_fd_sc_hd__o22a_4
X_24211_ _23383_/CLK _19514_/Y HRESETn VGND VGND VPWR VPWR _17357_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_72_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21423_ _21438_/A VGND VGND VPWR VPWR _21431_/A sky130_fd_sc_hd__buf_2
XFILLER_120_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24142_ _24137_/CLK _24142_/D HRESETn VGND VGND VPWR VPWR _17718_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_120_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21354_ _21290_/X _21348_/X _14052_/B _21352_/X VGND VGND VPWR VPWR _23904_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20305_ _20229_/X VGND VGND VPWR VPWR _20305_/X sky130_fd_sc_hd__buf_2
X_24073_ _24073_/CLK _21053_/X VGND VGND VPWR VPWR _24073_/Q sky130_fd_sc_hd__dfxtp_4
X_21285_ _21570_/A VGND VGND VPWR VPWR _21285_/X sky130_fd_sc_hd__buf_2
XFILLER_162_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23024_ _23024_/A VGND VGND VPWR VPWR HADDR[20] sky130_fd_sc_hd__inv_2
XANTENNA__22597__B2 _22591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20236_ _11590_/X VGND VGND VPWR VPWR _20863_/A sky130_fd_sc_hd__inv_2
XFILLER_104_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11917__A _12515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20167_ _24444_/Q VGND VGND VPWR VPWR _20167_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20098_ _11636_/Y _20146_/A _20192_/A VGND VGND VPWR VPWR _20098_/X sky130_fd_sc_hd__or3_4
XFILLER_57_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15108__B _24085_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23926_ _23192_/CLK _23926_/D VGND VGND VPWR VPWR _14871_/B sky130_fd_sc_hd__dfxtp_4
X_11940_ _16741_/A _11763_/B VGND VGND VPWR VPWR _11942_/B sky130_fd_sc_hd__or2_4
Xclkbuf_7_23_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR _24472_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_86_0_HCLK clkbuf_7_86_0_HCLK/A VGND VGND VPWR VPWR _23098_/CLK sky130_fd_sc_hd__clkbuf_1
X_11871_ _12186_/A VGND VGND VPWR VPWR _11872_/A sky130_fd_sc_hd__buf_2
X_23857_ _23761_/CLK _23857_/D VGND VGND VPWR VPWR _23857_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13610_ _13657_/A _13610_/B _13609_/X VGND VGND VPWR VPWR _13610_/X sky130_fd_sc_hd__and3_4
XFILLER_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11652__A _13865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22808_ _17319_/Y _22804_/X VGND VGND VPWR VPWR HWDATA[3] sky130_fd_sc_hd__nor2_4
X_14590_ _12530_/A _14590_/B VGND VGND VPWR VPWR _14590_/X sky130_fd_sc_hd__or2_4
X_23788_ _24045_/CLK _21547_/X VGND VGND VPWR VPWR _23788_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20965__A HRDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22521__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13541_ _13540_/X _23845_/Q VGND VGND VPWR VPWR _13541_/X sky130_fd_sc_hd__or2_4
XFILLER_38_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22739_ _19696_/X _22736_/X _22736_/X _23086_/C VGND VGND VPWR VPWR _22739_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16260_ _16287_/A _16260_/B VGND VGND VPWR VPWR _16260_/X sky130_fd_sc_hd__or2_4
X_13472_ _13441_/A _23237_/Q VGND VGND VPWR VPWR _13472_/X sky130_fd_sc_hd__or2_4
XANTENNA__23060__B _23079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15211_ _15198_/X _15211_/B VGND VGND VPWR VPWR _15212_/C sky130_fd_sc_hd__or2_4
X_12423_ _12423_/A _12423_/B VGND VGND VPWR VPWR _12423_/X sky130_fd_sc_hd__or2_4
X_24409_ _24445_/CLK _18881_/X HRESETn VGND VGND VPWR VPWR _24409_/Q sky130_fd_sc_hd__dfrtp_4
X_16191_ _11714_/A VGND VGND VPWR VPWR _16192_/A sky130_fd_sc_hd__buf_2
XFILLER_139_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21088__B2 _21087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11576__A1 _24462_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15142_ _14574_/A _15213_/B VGND VGND VPWR VPWR _15142_/X sky130_fd_sc_hd__or2_4
XFILLER_166_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12354_ _12354_/A VGND VGND VPWR VPWR _13529_/A sky130_fd_sc_hd__buf_2
XFILLER_153_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22037__B1 _23509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19950_ _19949_/X VGND VGND VPWR VPWR _19950_/X sky130_fd_sc_hd__buf_2
X_15073_ _15112_/A _15073_/B _15073_/C VGND VGND VPWR VPWR _15073_/X sky130_fd_sc_hd__and3_4
X_12285_ _12708_/A _12278_/X _12284_/X VGND VGND VPWR VPWR _12285_/X sky130_fd_sc_hd__or3_4
XFILLER_107_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18901_ _11851_/X _18897_/X _24404_/Q _18900_/X VGND VGND VPWR VPWR _24404_/D sky130_fd_sc_hd__o22a_4
X_14024_ _14074_/A _14020_/X _14024_/C VGND VGND VPWR VPWR _14024_/X sky130_fd_sc_hd__or3_4
X_19881_ _19556_/X _19811_/A _19876_/X _19880_/X VGND VGND VPWR VPWR _19881_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20599__B1 _20306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17464__B1 _17418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21260__B2 _21252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18832_ _16866_/X _18796_/A _24437_/Q _18790_/A VGND VGND VPWR VPWR _24437_/D sky130_fd_sc_hd__o22a_4
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18763_ _12021_/Y _17024_/X _17037_/Y _17031_/X VGND VGND VPWR VPWR _19963_/B sky130_fd_sc_hd__o22a_4
XFILLER_96_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15975_ _15956_/A _16041_/B VGND VGND VPWR VPWR _15977_/B sky130_fd_sc_hd__or2_4
XANTENNA__22420__A _22420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21012__A1 _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17714_ _18368_/A _17389_/X _17710_/B VGND VGND VPWR VPWR _17714_/X sky130_fd_sc_hd__a21bo_4
XANTENNA__21012__B2 _20282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14926_ _14772_/A VGND VGND VPWR VPWR _14973_/A sky130_fd_sc_hd__buf_2
X_18694_ _17326_/B _18692_/X _17793_/X _18693_/X VGND VGND VPWR VPWR _18694_/X sky130_fd_sc_hd__a211o_4
XFILLER_63_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13761__B _13761_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17645_ _17256_/X _17644_/X _17258_/A VGND VGND VPWR VPWR _17645_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20771__B1 _24096_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14857_ _12218_/A _23766_/Q VGND VGND VPWR VPWR _14858_/C sky130_fd_sc_hd__or2_4
XFILLER_95_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13808_ _12485_/A _23773_/Q VGND VGND VPWR VPWR _13809_/C sky130_fd_sc_hd__or2_4
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17576_ _17047_/X _17575_/X _17051_/X VGND VGND VPWR VPWR _17576_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__17519__A1 _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14788_ _14820_/A _14788_/B VGND VGND VPWR VPWR _14789_/C sky130_fd_sc_hd__or2_4
XFILLER_51_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19315_ _19228_/X VGND VGND VPWR VPWR _19315_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15969__A _15969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13739_ _12621_/X _13736_/X _13739_/C VGND VGND VPWR VPWR _13739_/X sky130_fd_sc_hd__and3_4
XFILLER_108_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16527_ _16527_/A _16527_/B VGND VGND VPWR VPWR _16527_/X sky130_fd_sc_hd__or2_4
XFILLER_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19246_ _19246_/A _19246_/B VGND VGND VPWR VPWR _19247_/B sky130_fd_sc_hd__and2_4
X_16458_ _16490_/A _16390_/B VGND VGND VPWR VPWR _16458_/X sky130_fd_sc_hd__or2_4
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13489__A _12923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15409_ _12191_/A _23330_/Q VGND VGND VPWR VPWR _15411_/B sky130_fd_sc_hd__or2_4
XANTENNA__21079__B2 _21042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16389_ _16006_/A _16389_/B _16389_/C VGND VGND VPWR VPWR _16389_/X sky130_fd_sc_hd__and3_4
X_19177_ _19154_/B VGND VGND VPWR VPWR _19177_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18128_ _17810_/X _17240_/X _18126_/X _17849_/X _18127_/X VGND VGND VPWR VPWR _18128_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_117_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18059_ _17583_/B _18059_/B VGND VGND VPWR VPWR _18059_/X sky130_fd_sc_hd__or2_4
XFILLER_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21070_ _21049_/A VGND VGND VPWR VPWR _21070_/X sky130_fd_sc_hd__buf_2
XFILLER_28_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20021_ _20020_/X VGND VGND VPWR VPWR _24154_/D sky130_fd_sc_hd__inv_2
XANTENNA__11737__A _12634_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17455__B1 _17418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19995__A2 _19983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17207__B1 _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13952__A _13952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21972_ _21857_/X _21967_/X _15540_/B _21971_/X VGND VGND VPWR VPWR _23553_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23711_ _23646_/CLK _21692_/X VGND VGND VPWR VPWR _23711_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13671__B _13760_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20923_ _20923_/A VGND VGND VPWR VPWR _20924_/A sky130_fd_sc_hd__inv_2
XFILLER_148_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12568__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24454__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24222__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23642_ _23101_/CLK _23642_/D VGND VGND VPWR VPWR _14601_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20854_ _18614_/Y _20702_/X _20753_/X _20853_/Y VGND VGND VPWR VPWR _20854_/X sky130_fd_sc_hd__a211o_4
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21306__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22503__B2 _22498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15879__A _13529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23573_ _23203_/CLK _23573_/D VGND VGND VPWR VPWR _23573_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_167_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20785_ _20785_/A _20730_/B VGND VGND VPWR VPWR _20785_/X sky130_fd_sc_hd__or2_4
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18255__A _18310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22524_ _22464_/X _22522_/X _13775_/B _22519_/X VGND VGND VPWR VPWR _22524_/X sky130_fd_sc_hd__o22a_4
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13399__A _13399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22267__B1 _23385_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22455_ _22454_/X _22450_/X _15454_/B _22445_/X VGND VGND VPWR VPWR _23266_/D sky130_fd_sc_hd__o22a_4
X_21406_ _21292_/X _21405_/X _23871_/Q _21402_/X VGND VGND VPWR VPWR _23871_/D sky130_fd_sc_hd__o22a_4
X_22386_ _22139_/X _22383_/X _15466_/B _22380_/X VGND VGND VPWR VPWR _23298_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22505__A _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24125_ _23416_/CLK _24125_/D HRESETn VGND VGND VPWR VPWR _24125_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21490__B2 _21489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21337_ _21261_/X _21334_/X _12268_/B _21331_/X VGND VGND VPWR VPWR _23916_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16503__A _16362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24056_ _23290_/CLK _21076_/X VGND VGND VPWR VPWR _24056_/Q sky130_fd_sc_hd__dfxtp_4
X_12070_ _11963_/A _12070_/B _12070_/C VGND VGND VPWR VPWR _12074_/B sky130_fd_sc_hd__and3_4
X_21268_ _21268_/A VGND VGND VPWR VPWR _21268_/X sky130_fd_sc_hd__buf_2
XANTENNA__13846__B _24093_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23007_ _22908_/A VGND VGND VPWR VPWR _23007_/X sky130_fd_sc_hd__buf_2
XANTENNA__21242__B2 _21240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20219_ _22039_/A _17415_/Y _21234_/B VGND VGND VPWR VPWR _20220_/A sky130_fd_sc_hd__or3_4
X_21199_ _20441_/X _21198_/X _23982_/Q _21195_/X VGND VGND VPWR VPWR _21199_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14023__A _11736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21793__A2 _21791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15760_ _12783_/X _15760_/B VGND VGND VPWR VPWR _15761_/C sky130_fd_sc_hd__or2_4
XFILLER_58_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12972_ _12972_/A _12972_/B _12971_/X VGND VGND VPWR VPWR _12976_/B sky130_fd_sc_hd__and3_4
XANTENNA__21545__A2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14711_ _14297_/A _14709_/X _14710_/X VGND VGND VPWR VPWR _14711_/X sky130_fd_sc_hd__and3_4
X_11923_ _16741_/A _11745_/B VGND VGND VPWR VPWR _11926_/B sky130_fd_sc_hd__or2_4
X_23909_ _23557_/CLK _23909_/D VGND VGND VPWR VPWR _23909_/Q sky130_fd_sc_hd__dfxtp_4
X_15691_ _13139_/A _15756_/B VGND VGND VPWR VPWR _15692_/C sky130_fd_sc_hd__or2_4
XANTENNA__12478__A _12537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22894__B _22894_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17430_ _17429_/X VGND VGND VPWR VPWR _17434_/A sky130_fd_sc_hd__inv_2
X_14642_ _14841_/A _14629_/X _14642_/C VGND VGND VPWR VPWR _14642_/X sky130_fd_sc_hd__and3_4
X_11854_ _11854_/A VGND VGND VPWR VPWR _11855_/A sky130_fd_sc_hd__buf_2
XANTENNA__24124__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20695__A _20231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17361_ _17353_/Y _17354_/X _17027_/X _17360_/X VGND VGND VPWR VPWR _17445_/B sky130_fd_sc_hd__o22a_4
X_14573_ _14292_/A _14573_/B _14573_/C VGND VGND VPWR VPWR _14573_/X sky130_fd_sc_hd__or3_4
XPHY_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ _11784_/X VGND VGND VPWR VPWR _16222_/A sky130_fd_sc_hd__buf_2
XPHY_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19100_ _19098_/Y _19099_/Y _11521_/X VGND VGND VPWR VPWR _19100_/X sky130_fd_sc_hd__o21a_4
XPHY_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13524_ _13521_/X _13524_/B _13524_/C VGND VGND VPWR VPWR _13524_/X sky130_fd_sc_hd__and3_4
X_16312_ _16195_/A _16248_/B VGND VGND VPWR VPWR _16313_/C sky130_fd_sc_hd__or2_4
XFILLER_41_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17292_ _17290_/X _17292_/B VGND VGND VPWR VPWR _17292_/X sky130_fd_sc_hd__or2_4
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19031_ _19029_/Y _19030_/Y _11533_/X VGND VGND VPWR VPWR _19031_/X sky130_fd_sc_hd__o21a_4
X_16243_ _16162_/X _16243_/B VGND VGND VPWR VPWR _16243_/X sky130_fd_sc_hd__or2_4
X_13455_ _13455_/A _23909_/Q VGND VGND VPWR VPWR _13455_/X sky130_fd_sc_hd__or2_4
XANTENNA__14735__A1 _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12406_ _15894_/A _12400_/X _12406_/C VGND VGND VPWR VPWR _12416_/B sky130_fd_sc_hd__or3_4
XFILLER_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16174_ _16220_/A _16171_/X _16173_/X VGND VGND VPWR VPWR _16175_/C sky130_fd_sc_hd__and3_4
X_13386_ _13410_/A _13384_/X _13386_/C VGND VGND VPWR VPWR _13392_/B sky130_fd_sc_hd__and3_4
XANTENNA__19674__A1 _19469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15125_ _12433_/A _15125_/B VGND VGND VPWR VPWR _15125_/X sky130_fd_sc_hd__or2_4
XFILLER_115_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12337_ _12337_/A VGND VGND VPWR VPWR _12401_/A sky130_fd_sc_hd__buf_2
XANTENNA__21481__B2 _21475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12941__A _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19933_ _19931_/X _24174_/Q _19932_/X _20776_/A VGND VGND VPWR VPWR _19933_/X sky130_fd_sc_hd__o22a_4
XFILLER_5_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15056_ _15086_/A _23733_/Q VGND VGND VPWR VPWR _15057_/C sky130_fd_sc_hd__or2_4
X_12268_ _12689_/A _12268_/B VGND VGND VPWR VPWR _12268_/X sky130_fd_sc_hd__or2_4
XANTENNA__19360__A1_N _19358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14007_ _12467_/A _14007_/B _14007_/C VGND VGND VPWR VPWR _14007_/X sky130_fd_sc_hd__and3_4
XANTENNA__15029__A _15029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19724__A _19724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19864_ _21319_/A VGND VGND VPWR VPWR _21184_/C sky130_fd_sc_hd__buf_2
X_12199_ _12512_/A VGND VGND VPWR VPWR _12569_/A sky130_fd_sc_hd__buf_2
XFILLER_122_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18815_ _17169_/X _18810_/X _20161_/A _18811_/X VGND VGND VPWR VPWR _24450_/D sky130_fd_sc_hd__o22a_4
X_19795_ _19744_/A _19765_/B _19613_/X VGND VGND VPWR VPWR _19795_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14868__A _14110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13772__A _12925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17244__A _12027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24245__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18746_ _17817_/X _18744_/X _18745_/X _17816_/X _17126_/X VGND VGND VPWR VPWR _18746_/X
+ sky130_fd_sc_hd__a32o_4
X_15958_ _13431_/X VGND VGND VPWR VPWR _15959_/A sky130_fd_sc_hd__buf_2
XFILLER_36_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22733__A1 _21311_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22733__B2 _22698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14909_ _11625_/A _14908_/X VGND VGND VPWR VPWR _14909_/X sky130_fd_sc_hd__and2_4
X_18677_ _17805_/X _17979_/Y _17869_/A _18676_/Y VGND VGND VPWR VPWR _18677_/X sky130_fd_sc_hd__a211o_4
X_15889_ _13532_/A _15827_/B VGND VGND VPWR VPWR _15889_/X sky130_fd_sc_hd__or2_4
XANTENNA__12388__A _15887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17628_ _18714_/B _17627_/X _17333_/X VGND VGND VPWR VPWR _17628_/X sky130_fd_sc_hd__o21a_4
XFILLER_23_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15699__A _12298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17559_ _17558_/X VGND VGND VPWR VPWR _17660_/B sky130_fd_sc_hd__inv_2
XFILLER_149_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18075__A _17792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20570_ _20570_/A VGND VGND VPWR VPWR _20570_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19229_ _24280_/Q _19228_/X VGND VGND VPWR VPWR _19313_/A sky130_fd_sc_hd__and2_4
XFILLER_20_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18803__A _18796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22240_ _22115_/X _22237_/X _12392_/B _22234_/X VGND VGND VPWR VPWR _23404_/D sky130_fd_sc_hd__o22a_4
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22171_ _11828_/B VGND VGND VPWR VPWR _22171_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12851__A _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21122_ _21101_/A VGND VGND VPWR VPWR _21122_/X sky130_fd_sc_hd__buf_2
XANTENNA__19417__B2 _24226_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17428__B1 _17028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21053_ _20559_/X _21052_/X _24073_/Q _21049_/X VGND VGND VPWR VPWR _21053_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21224__B2 _21223_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21775__A2 _21770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20004_ _18067_/X _19983_/X _20003_/Y _19994_/X VGND VGND VPWR VPWR _20004_/X sky130_fd_sc_hd__o22a_4
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22060__A _22060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14778__A _15112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13682__A _12190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22724__A1 _20819_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22724__B2 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21955_ _21829_/X _21953_/X _16203_/B _21950_/X VGND VGND VPWR VPWR _21955_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23612__CLK _23675_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12298__A _12298_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16993__A _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _20755_/X _20905_/X _11520_/A _20708_/X VGND VGND VPWR VPWR _20906_/X sky130_fd_sc_hd__o22a_4
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21886_ _21885_/X _21839_/A _23605_/Q _21809_/X VGND VGND VPWR VPWR _21886_/X sky130_fd_sc_hd__o22a_4
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23625_ _24073_/CLK _21840_/X VGND VGND VPWR VPWR _23625_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _24253_/Q _20661_/X _20836_/X VGND VGND VPWR VPWR _20837_/X sky130_fd_sc_hd__o21a_4
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11930__A _11930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23556_ _23588_/CLK _23556_/D VGND VGND VPWR VPWR _15675_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _11564_/X _11570_/B VGND VGND VPWR VPWR _20111_/D sky130_fd_sc_hd__or2_4
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20768_ _24224_/Q _20636_/X _20767_/Y VGND VGND VPWR VPWR _22459_/A sky130_fd_sc_hd__o21a_4
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22507_ _22435_/X _22501_/X _12836_/B _22505_/X VGND VGND VPWR VPWR _23242_/D sky130_fd_sc_hd__o22a_4
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23487_ _23518_/CLK _22075_/X VGND VGND VPWR VPWR _23487_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_161_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20699_ _20339_/B _20844_/B VGND VGND VPWR VPWR _20699_/X sky130_fd_sc_hd__or2_4
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14018__A _13888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20962__B _20776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13240_ _13252_/A _13240_/B VGND VGND VPWR VPWR _13240_/X sky130_fd_sc_hd__or2_4
XFILLER_109_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22438_ _22438_/A VGND VGND VPWR VPWR _22438_/X sky130_fd_sc_hd__buf_2
XANTENNA__24118__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21463__A1 _21304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13171_ _13303_/A _13240_/B VGND VGND VPWR VPWR _13173_/B sky130_fd_sc_hd__or2_4
XANTENNA__21463__B2 _21459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13857__A _15446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12761__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22369_ _22376_/A VGND VGND VPWR VPWR _22369_/X sky130_fd_sc_hd__buf_2
XFILLER_163_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24108_ _24074_/CLK _20487_/X VGND VGND VPWR VPWR _24108_/Q sky130_fd_sc_hd__dfxtp_4
X_12122_ _12122_/A _12119_/X _12121_/X VGND VGND VPWR VPWR _12123_/C sky130_fd_sc_hd__and3_4
XANTENNA__12480__B _12608_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17419__B1 _17020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24039_ _24039_/CLK _21107_/X VGND VGND VPWR VPWR _24039_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21215__B2 _21209_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19544__A _19888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16930_ _11596_/A _16936_/A _11592_/A _16929_/X VGND VGND VPWR VPWR _17297_/A sky130_fd_sc_hd__or4_4
X_12053_ _16725_/A _12053_/B _12052_/X VGND VGND VPWR VPWR _12054_/C sky130_fd_sc_hd__and3_4
XANTENNA__24268__CLK _24495_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21766__A2 _21763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22692__A2_N _22691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16861_ _15391_/D _13950_/X _13949_/A VGND VGND VPWR VPWR _16861_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20974__B1 _20662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14688__A _15620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18600_ _18600_/A _17300_/X VGND VGND VPWR VPWR _18600_/X sky130_fd_sc_hd__or2_4
XANTENNA__13592__A _13965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15812_ _12851_/A _15810_/X _15811_/X VGND VGND VPWR VPWR _15812_/X sky130_fd_sc_hd__and3_4
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19580_ _19445_/A _19579_/X HRDATA[9] _19461_/A VGND VGND VPWR VPWR _19581_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24305__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16792_ _16811_/A _24081_/Q VGND VGND VPWR VPWR _16792_/X sky130_fd_sc_hd__or2_4
XANTENNA__21518__A2 _21513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18531_ _18399_/X VGND VGND VPWR VPWR _18531_/X sky130_fd_sc_hd__buf_2
X_12955_ _12955_/A _23145_/Q VGND VGND VPWR VPWR _12957_/B sky130_fd_sc_hd__or2_4
X_15743_ _13205_/A VGND VGND VPWR VPWR _15743_/X sky130_fd_sc_hd__buf_2
XFILLER_46_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18395__B2 _18394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11906_ _11905_/X VGND VGND VPWR VPWR _11941_/A sky130_fd_sc_hd__buf_2
XFILLER_18_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18462_ _18409_/A _18459_/X _18460_/X _18462_/D VGND VGND VPWR VPWR _18462_/X sky130_fd_sc_hd__or4_4
X_12886_ _12886_/A _12884_/X _12886_/C VGND VGND VPWR VPWR _12886_/X sky130_fd_sc_hd__and3_4
X_15674_ _12735_/A _15746_/B VGND VGND VPWR VPWR _15674_/X sky130_fd_sc_hd__or2_4
XANTENNA__12001__A _12001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_56_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17413_ _17412_/X VGND VGND VPWR VPWR _17436_/B sky130_fd_sc_hd__buf_2
X_11837_ _16647_/A _11837_/B _11837_/C VGND VGND VPWR VPWR _11838_/C sky130_fd_sc_hd__and3_4
X_14625_ _13868_/A VGND VGND VPWR VPWR _14669_/A sky130_fd_sc_hd__buf_2
XANTENNA__22479__B1 _15253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18393_ _17499_/Y _18391_/X _17648_/X VGND VGND VPWR VPWR _18393_/X sky130_fd_sc_hd__o21a_4
XFILLER_159_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12936__A _12943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__A _11768_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _17343_/X VGND VGND VPWR VPWR _17751_/B sky130_fd_sc_hd__inv_2
X_14556_ _14278_/A _23354_/Q VGND VGND VPWR VPWR _14556_/X sky130_fd_sc_hd__or2_4
XANTENNA__21151__B1 _24012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11768_ _16048_/A VGND VGND VPWR VPWR _11768_/X sky130_fd_sc_hd__buf_2
XFILLER_144_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12655__B _12655_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13507_ _13535_/A _23301_/Q VGND VGND VPWR VPWR _13507_/X sky130_fd_sc_hd__or2_4
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15031__B _24085_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14487_ _14506_/A _14487_/B VGND VGND VPWR VPWR _14487_/X sky130_fd_sc_hd__or2_4
X_17275_ _16936_/A _17044_/B VGND VGND VPWR VPWR _17275_/X sky130_fd_sc_hd__and2_4
X_11699_ _12604_/A VGND VGND VPWR VPWR _13223_/A sky130_fd_sc_hd__buf_2
X_19014_ _18987_/X _19012_/Y _19013_/Y _18990_/X VGND VGND VPWR VPWR _19014_/X sky130_fd_sc_hd__o22a_4
X_13438_ _13474_/A _13438_/B _13438_/C VGND VGND VPWR VPWR _13445_/B sky130_fd_sc_hd__and3_4
X_16226_ _16202_/A _16226_/B VGND VGND VPWR VPWR _16226_/X sky130_fd_sc_hd__or2_4
XFILLER_173_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16157_ _16157_/A _23885_/Q VGND VGND VPWR VPWR _16158_/C sky130_fd_sc_hd__or2_4
X_13369_ _13378_/A _23174_/Q VGND VGND VPWR VPWR _13372_/B sky130_fd_sc_hd__or2_4
XANTENNA__21454__B2 _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15108_ _15096_/A _24085_/Q VGND VGND VPWR VPWR _15108_/X sky130_fd_sc_hd__or2_4
X_16088_ _16088_/A VGND VGND VPWR VPWR _16089_/B sky130_fd_sc_hd__inv_2
XANTENNA__21206__B2 _21202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19916_ _23083_/D _19915_/X VGND VGND VPWR VPWR _22904_/D sky130_fd_sc_hd__or2_4
X_15039_ _12467_/A _15039_/B _15039_/C VGND VGND VPWR VPWR _15043_/B sky130_fd_sc_hd__and3_4
XANTENNA__22403__B1 _23285_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19847_ _19471_/X _19687_/C _19844_/Y _21134_/A _19512_/X VGND VGND VPWR VPWR _19847_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_69_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14598__A _13656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19778_ _19683_/A _19778_/B _19711_/A VGND VGND VPWR VPWR _19811_/B sky130_fd_sc_hd__or3_4
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21509__A2 _21506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22706__B2 _22705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18729_ _17341_/X _17346_/Y _17341_/X _17346_/Y VGND VGND VPWR VPWR _18729_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17189__A2 _17187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22182__A2 _22180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13007__A _12570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23785__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21740_ _21575_/X _21734_/X _23680_/Q _21738_/X VGND VGND VPWR VPWR _23680_/D sky130_fd_sc_hd__o22a_4
XFILLER_92_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21671_ _21541_/X _21670_/X _23726_/Q _21667_/X VGND VGND VPWR VPWR _21671_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17421__B _17421_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22039__B _22039_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23410_ _23204_/CLK _22232_/X VGND VGND VPWR VPWR _16664_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20622_ _20490_/X _20621_/Y _19242_/A _20584_/X VGND VGND VPWR VPWR _20622_/X sky130_fd_sc_hd__o22a_4
X_24390_ _24422_/CLK _24390_/D HRESETn VGND VGND VPWR VPWR _24390_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__12565__B _12565_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19886__B2 _19823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23341_ _24077_/CLK _23341_/D VGND VGND VPWR VPWR _23341_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17897__B1 _17653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20553_ _20552_/X VGND VGND VPWR VPWR _20553_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23272_ _23656_/CLK _23272_/D VGND VGND VPWR VPWR _12988_/B sky130_fd_sc_hd__dfxtp_4
X_20484_ _24236_/Q _20420_/X _20483_/Y VGND VGND VPWR VPWR _20485_/A sky130_fd_sc_hd__o21a_4
XANTENNA__17649__B1 _17648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22223_ _21134_/B _21134_/C _21236_/D VGND VGND VPWR VPWR _22223_/X sky130_fd_sc_hd__or3_4
XFILLER_118_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12581__A _12581_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16053__A _16053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20653__C1 _20652_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22154_ _22118_/A VGND VGND VPWR VPWR _22154_/X sky130_fd_sc_hd__buf_2
XANTENNA__21894__A _21923_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21105_ _20559_/X _21104_/X _24041_/Q _21101_/X VGND VGND VPWR VPWR _24041_/D sky130_fd_sc_hd__o22a_4
X_22085_ _21881_/X _22081_/X _15169_/B _22042_/X VGND VGND VPWR VPWR _22085_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21036_ _21026_/Y _21035_/X _20299_/X _21035_/X VGND VGND VPWR VPWR _24084_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19810__A1 _19888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20303__A _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17821__B1 _17817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11925__A _16742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14301__A _14301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22987_ _22977_/X _18368_/A _22959_/X _22986_/X VGND VGND VPWR VPWR _22987_/X sky130_fd_sc_hd__a211o_4
XANTENNA__12110__A1 _12077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12740_ _13333_/A _23658_/Q VGND VGND VPWR VPWR _12741_/C sky130_fd_sc_hd__or2_4
XFILLER_83_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21938_ _21028_/A VGND VGND VPWR VPWR _22173_/B sky130_fd_sc_hd__buf_2
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14955__B _14884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21134__A _21134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12671_ _12973_/A _12671_/B VGND VGND VPWR VPWR _12671_/X sky130_fd_sc_hd__or2_4
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ _20860_/A VGND VGND VPWR VPWR _21869_/X sky130_fd_sc_hd__buf_2
XANTENNA__12756__A _13052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _12576_/A _14402_/X _14410_/C VGND VGND VPWR VPWR _14410_/X sky130_fd_sc_hd__and3_4
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23608_ _23416_/CLK _21880_/X VGND VGND VPWR VPWR _15351_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15132__A _14897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11622_ _12188_/A VGND VGND VPWR VPWR _11623_/A sky130_fd_sc_hd__buf_2
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _14417_/X _14552_/Y _15388_/X _14417_/B _15389_/X VGND VGND VPWR VPWR _15391_/D
+ sky130_fd_sc_hd__o32a_4
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _13720_/A VGND VGND VPWR VPWR _14512_/A sky130_fd_sc_hd__buf_2
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23539_ _23889_/CLK _21997_/X VGND VGND VPWR VPWR _23539_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _24440_/Q IRQ[3] _11552_/Y VGND VGND VPWR VPWR _11553_/X sky130_fd_sc_hd__a21bo_4
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19539__A _19539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22881__B1 _13692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17060_ _17060_/A _17060_/B VGND VGND VPWR VPWR _17060_/X sky130_fd_sc_hd__or2_4
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _14272_/A VGND VGND VPWR VPWR _14280_/A sky130_fd_sc_hd__buf_2
X_16011_ _16011_/A _16011_/B _16011_/C VGND VGND VPWR VPWR _16012_/C sky130_fd_sc_hd__and3_4
X_13223_ _13223_/A _13220_/X _13223_/C VGND VGND VPWR VPWR _13227_/B sky130_fd_sc_hd__and3_4
XFILLER_87_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21436__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13587__A _11928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12491__A _12571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21987__A2 _21960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13154_ _12748_/A _13152_/X _13154_/C VGND VGND VPWR VPWR _13154_/X sky130_fd_sc_hd__and3_4
XFILLER_152_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12105_ _12105_/A _23731_/Q VGND VGND VPWR VPWR _12107_/B sky130_fd_sc_hd__or2_4
X_13085_ _13085_/A _24008_/Q VGND VGND VPWR VPWR _13086_/C sky130_fd_sc_hd__or2_4
X_17962_ _17900_/X _17961_/X _19993_/A _17900_/X VGND VGND VPWR VPWR _24497_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21739__A2 _21734_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19701_ _19441_/X _19699_/X _17875_/X _19700_/X VGND VGND VPWR VPWR _19701_/X sky130_fd_sc_hd__o22a_4
X_16913_ _16905_/A _16912_/Y _16905_/A _16912_/Y VGND VGND VPWR VPWR _16914_/A sky130_fd_sc_hd__a2bb2o_4
X_12036_ _16702_/A _12036_/B _12036_/C VGND VGND VPWR VPWR _12043_/B sky130_fd_sc_hd__and3_4
XFILLER_137_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17893_ _16943_/X _17789_/X _17014_/X _17892_/X VGND VGND VPWR VPWR _17893_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11835__A _11792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20411__A2 _20399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19632_ _19797_/A _19630_/X _19600_/X _19631_/X VGND VGND VPWR VPWR _19632_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15307__A _13952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16844_ _15521_/X _16843_/X _15521_/X _16843_/X VGND VGND VPWR VPWR _16852_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19563_ _19528_/B _19562_/X VGND VGND VPWR VPWR _19563_/X sky130_fd_sc_hd__or2_4
XANTENNA__11554__B IRQ[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16775_ _16775_/A VGND VGND VPWR VPWR _16811_/A sky130_fd_sc_hd__buf_2
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13987_ _13607_/A _24064_/Q VGND VGND VPWR VPWR _13987_/X sky130_fd_sc_hd__or2_4
XANTENNA__20867__B _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22164__A2 _22159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18514_ _17436_/C _18512_/X VGND VGND VPWR VPWR _18514_/X sky130_fd_sc_hd__or2_4
X_15726_ _12758_/A _15726_/B VGND VGND VPWR VPWR _15726_/X sky130_fd_sc_hd__or2_4
XANTENNA__17522__A _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12938_ _12976_/A _12938_/B _12937_/X VGND VGND VPWR VPWR _12946_/B sky130_fd_sc_hd__or3_4
X_19494_ _19494_/A _19705_/B VGND VGND VPWR VPWR _19548_/B sky130_fd_sc_hd__or2_4
XFILLER_46_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21911__A2 _21909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14865__B _23990_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18445_ _17250_/X _18421_/X _17250_/X _18417_/B VGND VGND VPWR VPWR _18445_/X sky130_fd_sc_hd__a2bb2o_4
X_15657_ _12693_/A _15657_/B VGND VGND VPWR VPWR _15659_/B sky130_fd_sc_hd__or2_4
X_12869_ _12869_/A _12869_/B _12869_/C VGND VGND VPWR VPWR _12874_/B sky130_fd_sc_hd__and3_4
XANTENNA__16138__A _16138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12666__A _12944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14608_ _13655_/A _14688_/B VGND VGND VPWR VPWR _14609_/C sky130_fd_sc_hd__or2_4
XFILLER_15_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18376_ _18376_/A _17530_/B VGND VGND VPWR VPWR _18379_/B sky130_fd_sc_hd__nor2_4
X_15588_ _15606_/A VGND VGND VPWR VPWR _15611_/A sky130_fd_sc_hd__buf_2
XFILLER_159_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17327_ _15185_/X VGND VGND VPWR VPWR _17327_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21675__B2 _21674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14539_ _14520_/A _24091_/Q VGND VGND VPWR VPWR _14540_/C sky130_fd_sc_hd__or2_4
XFILLER_18_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17258_ _17258_/A VGND VGND VPWR VPWR _17259_/B sky130_fd_sc_hd__inv_2
XFILLER_174_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16209_ _16216_/A _23981_/Q VGND VGND VPWR VPWR _16210_/C sky130_fd_sc_hd__or2_4
XANTENNA__13497__A _13547_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17189_ _17160_/X _17187_/X _17236_/B VGND VGND VPWR VPWR _17189_/X sky130_fd_sc_hd__o21a_4
XFILLER_143_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21219__A _21219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22910_ _19957_/A _22910_/B VGND VGND VPWR VPWR _22910_/X sky130_fd_sc_hd__or2_4
XFILLER_99_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15217__A _14663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23890_ _23728_/CLK _23890_/D VGND VGND VPWR VPWR _23890_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22841_ _15915_/Y _22836_/X _22817_/X _22840_/X VGND VGND VPWR VPWR _22842_/B sky130_fd_sc_hd__o22a_4
XFILLER_99_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22155__A2 _22147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24383__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17432__A _14261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22772_ _22749_/Y _22769_/X VGND VGND VPWR VPWR _24118_/D sky130_fd_sc_hd__and2_4
XFILLER_25_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21723_ _21546_/X _21720_/X _23692_/Q _21717_/X VGND VGND VPWR VPWR _21723_/X sky130_fd_sc_hd__o22a_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12576__A _12576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16048__A _16048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24442_ _24445_/CLK _18827_/X HRESETn VGND VGND VPWR VPWR _24442_/Q sky130_fd_sc_hd__dfrtp_4
X_21654_ _21600_/X _21620_/A _23733_/Q _21617_/A VGND VGND VPWR VPWR _23733_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20605_ _20515_/X _20604_/X _19147_/A _20522_/X VGND VGND VPWR VPWR _20605_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15887__A _15887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21666__B2 _21660_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24373_ _24422_/CLK _24373_/D HRESETn VGND VGND VPWR VPWR _24373_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_123_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21585_ _21549_/A VGND VGND VPWR VPWR _21585_/X sky130_fd_sc_hd__buf_2
X_23324_ _23880_/CLK _23324_/D VGND VGND VPWR VPWR _22346_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_165_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20536_ _20444_/X _20917_/B _20308_/X VGND VGND VPWR VPWR _20536_/X sky130_fd_sc_hd__a21o_4
XFILLER_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23255_ _23192_/CLK _23255_/D VGND VGND VPWR VPWR _15122_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21418__B2 _21381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20467_ _20380_/A _20844_/A VGND VGND VPWR VPWR _20467_/X sky130_fd_sc_hd__and2_4
XANTENNA__21969__A2 _21967_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13200__A _12362_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20626__C1 _20625_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22206_ _22141_/X _22201_/X _15563_/B _22205_/X VGND VGND VPWR VPWR _22206_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23186_ _23537_/CLK _22596_/X VGND VGND VPWR VPWR _16638_/B sky130_fd_sc_hd__dfxtp_4
X_20398_ _20234_/X VGND VGND VPWR VPWR _20398_/X sky130_fd_sc_hd__buf_2
XANTENNA__19806__B _19705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22137_ _20692_/A VGND VGND VPWR VPWR _22137_/X sky130_fd_sc_hd__buf_2
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16511__A _16362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22918__B2 _22930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22068_ _21850_/X _22067_/X _15701_/B _22064_/X VGND VGND VPWR VPWR _23492_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11655__A _15595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21019_ _24245_/Q VGND VGND VPWR VPWR _21019_/Y sky130_fd_sc_hd__inv_2
X_13910_ _14335_/A _13910_/B _13910_/C VGND VGND VPWR VPWR _13911_/C sky130_fd_sc_hd__or3_4
X_14890_ _14127_/A _14961_/B VGND VGND VPWR VPWR _14890_/X sky130_fd_sc_hd__or2_4
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_121_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR _23496_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24306__CLK _24306_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13841_ _13658_/A _13841_/B VGND VGND VPWR VPWR _13841_/X sky130_fd_sc_hd__or2_4
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13870__A _13885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13772_ _12925_/A _13772_/B VGND VGND VPWR VPWR _13774_/B sky130_fd_sc_hd__or2_4
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16560_ _16588_/A _16560_/B _16560_/C VGND VGND VPWR VPWR _16561_/C sky130_fd_sc_hd__and3_4
X_15511_ _13053_/A _15511_/B VGND VGND VPWR VPWR _15511_/X sky130_fd_sc_hd__or2_4
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12723_ _13277_/A _12723_/B VGND VGND VPWR VPWR _12725_/B sky130_fd_sc_hd__or2_4
XANTENNA__12486__A _13010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16491_ _16491_/A _16422_/B VGND VGND VPWR VPWR _16492_/C sky130_fd_sc_hd__or2_4
XFILLER_16_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18230_ _17976_/X _18049_/X _17883_/X VGND VGND VPWR VPWR _18230_/Y sky130_fd_sc_hd__o21ai_4
X_12654_ _12623_/A VGND VGND VPWR VPWR _12942_/A sky130_fd_sc_hd__buf_2
X_15442_ _15442_/A _15442_/B _15441_/X VGND VGND VPWR VPWR _15442_/X sky130_fd_sc_hd__or3_4
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11605_ _11605_/A VGND VGND VPWR VPWR _11606_/A sky130_fd_sc_hd__buf_2
XANTENNA__15797__A _12848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18161_ _17809_/X _18160_/Y _17848_/X _18133_/X VGND VGND VPWR VPWR _18161_/X sky130_fd_sc_hd__o22a_4
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12957_/A _12579_/X _12585_/C VGND VGND VPWR VPWR _12585_/X sky130_fd_sc_hd__and3_4
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15373_ _11659_/A _15300_/B VGND VGND VPWR VPWR _15373_/X sky130_fd_sc_hd__or2_4
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17112_ _12078_/X VGND VGND VPWR VPWR _17112_/X sky130_fd_sc_hd__buf_2
X_14324_ _11933_/A _14324_/B _14323_/X VGND VGND VPWR VPWR _14324_/X sky130_fd_sc_hd__or3_4
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11536_ _11536_/A _11535_/X VGND VGND VPWR VPWR _11537_/B sky130_fd_sc_hd__or2_4
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18092_ _18562_/A _18091_/Y VGND VGND VPWR VPWR _18092_/X sky130_fd_sc_hd__and2_4
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22606__B1 _12520_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17043_ _17043_/A _17481_/B VGND VGND VPWR VPWR _17044_/B sky130_fd_sc_hd__or2_4
X_14255_ _15606_/A _23647_/Q VGND VGND VPWR VPWR _14256_/C sky130_fd_sc_hd__or2_4
XFILLER_109_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13206_ _13232_/A _13204_/X _13205_/X VGND VGND VPWR VPWR _13210_/B sky130_fd_sc_hd__and3_4
X_14186_ _15324_/A VGND VGND VPWR VPWR _14191_/A sky130_fd_sc_hd__buf_2
XANTENNA__22082__B2 _22078_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22423__A _20415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13137_ _12745_/A VGND VGND VPWR VPWR _13170_/A sky130_fd_sc_hd__buf_2
XANTENNA__16421__A _16007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24320__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18994_ _18994_/A VGND VGND VPWR VPWR _18994_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13068_ _13097_/A _24040_/Q VGND VGND VPWR VPWR _13071_/B sky130_fd_sc_hd__or2_4
X_17945_ _17836_/X VGND VGND VPWR VPWR _17945_/X sky130_fd_sc_hd__buf_2
XANTENNA__22385__A2 _22383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12019_ _11984_/X _11992_/X _11999_/X _12010_/X _12018_/X VGND VGND VPWR VPWR _12019_/X
+ sky130_fd_sc_hd__a32o_4
X_17876_ _17151_/X VGND VGND VPWR VPWR _17876_/X sky130_fd_sc_hd__buf_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19615_ _19450_/A _19506_/A VGND VGND VPWR VPWR _19615_/X sky130_fd_sc_hd__or2_4
XFILLER_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16827_ _16905_/B _16826_/X _12183_/X VGND VGND VPWR VPWR _16827_/X sky130_fd_sc_hd__o21a_4
XFILLER_81_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13780__A _11813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19546_ _19546_/A _19831_/A VGND VGND VPWR VPWR _19546_/X sky130_fd_sc_hd__or2_4
X_16758_ _16757_/X _23761_/Q VGND VGND VPWR VPWR _16759_/C sky130_fd_sc_hd__or2_4
XFILLER_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15709_ _13184_/A _23812_/Q VGND VGND VPWR VPWR _15710_/C sky130_fd_sc_hd__or2_4
XFILLER_146_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21896__B2 _21892_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19477_ _24179_/Q _19457_/X _20246_/B _19454_/X VGND VGND VPWR VPWR _19477_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12396__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16689_ _16686_/X _16689_/B VGND VGND VPWR VPWR _16824_/A sky130_fd_sc_hd__or2_4
Xclkbuf_5_26_0_HCLK clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18428_ _17767_/C _17714_/X _17710_/B VGND VGND VPWR VPWR _18428_/X sky130_fd_sc_hd__o21a_4
X_18359_ _17708_/A VGND VGND VPWR VPWR _18402_/A sky130_fd_sc_hd__buf_2
XFILLER_159_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15500__A _12616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21370_ _21184_/A _21370_/B _21134_/C _21184_/D VGND VGND VPWR VPWR _21370_/X sky130_fd_sc_hd__or4_4
XANTENNA__24479__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20118__A NMI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12843__B _12842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20321_ _18891_/X _20318_/Y _20320_/X _18952_/Y _20275_/X VGND VGND VPWR VPWR _20321_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_134_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14116__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13020__A _12877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23040_ _23051_/A _23038_/Y _23040_/C VGND VGND VPWR VPWR _23040_/X sky130_fd_sc_hd__and3_4
XFILLER_31_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20252_ _18780_/X _20246_/B _20251_/X VGND VGND VPWR VPWR _20252_/X sky130_fd_sc_hd__a21o_4
XANTENNA__22073__B2 _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13955__A _13955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17427__A _17427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21820__B2 _21810_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20183_ _24460_/Q IRQ[23] _20182_/X VGND VGND VPWR VPWR _20183_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__23203__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24329__CLK _24342_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23942_ _23397_/CLK _23942_/D VGND VGND VPWR VPWR _13364_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23873_ _23649_/CLK _21403_/X VGND VGND VPWR VPWR _15638_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_151_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22128__A2 _22123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11625__D _11886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22824_ _13692_/Y _22816_/X _22818_/X _22823_/X VGND VGND VPWR VPWR _22825_/B sky130_fd_sc_hd__o22a_4
XANTENNA__17162__A _17161_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24479__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22755_ SYSTICKCLKDIV[3] VGND VGND VPWR VPWR _22755_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21706_ _21706_/A _21420_/B _21706_/C _22487_/B VGND VGND VPWR VPWR _21706_/X sky130_fd_sc_hd__or4_4
XFILLER_25_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22686_ _23124_/Q VGND VGND VPWR VPWR _22686_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22508__A _22508_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21412__A _21405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24425_ _24422_/CLK _18859_/X HRESETn VGND VGND VPWR VPWR _20541_/A sky130_fd_sc_hd__dfrtp_4
X_21637_ _21570_/X _21634_/X _23746_/Q _21631_/X VGND VGND VPWR VPWR _21637_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21639__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22300__A2 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19701__B1 _17875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12370_ _12370_/A _24012_/Q VGND VGND VPWR VPWR _12370_/X sky130_fd_sc_hd__or2_4
XFILLER_21_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24356_ _24388_/CLK _24356_/D HRESETn VGND VGND VPWR VPWR _11530_/A sky130_fd_sc_hd__dfstp_4
X_21568_ _21283_/A VGND VGND VPWR VPWR _21568_/X sky130_fd_sc_hd__buf_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23307_ _23558_/CLK _23307_/D VGND VGND VPWR VPWR _12611_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_5_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20519_ _20349_/A VGND VGND VPWR VPWR _20519_/X sky130_fd_sc_hd__buf_2
XFILLER_165_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24287_ _24287_/CLK _24287_/D HRESETn VGND VGND VPWR VPWR _24287_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_46_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR _23501_/CLK sky130_fd_sc_hd__clkbuf_1
X_21499_ _21492_/A VGND VGND VPWR VPWR _21499_/X sky130_fd_sc_hd__buf_2
XANTENNA__24149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14026__A _13705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14040_ _11698_/A _14038_/X _14040_/C VGND VGND VPWR VPWR _14041_/C sky130_fd_sc_hd__and3_4
X_23238_ _24102_/CLK _22513_/X VGND VGND VPWR VPWR _23238_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13865__A _13865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23169_ _23203_/CLK _23169_/D VGND VGND VPWR VPWR _15546_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16241__A _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15991_ _15957_/A _23406_/Q VGND VGND VPWR VPWR _15993_/B sky130_fd_sc_hd__or2_4
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22367__A2 _22362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22897__B _22896_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19768__B1 _19687_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17730_ _17730_/A _17730_/B VGND VGND VPWR VPWR _17730_/X sky130_fd_sc_hd__or2_4
X_14942_ _14973_/A _14864_/B VGND VGND VPWR VPWR _14942_/X sky130_fd_sc_hd__or2_4
XFILLER_134_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20698__A HRDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23074__A _17650_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17661_ _17661_/A VGND VGND VPWR VPWR _17661_/X sky130_fd_sc_hd__buf_2
X_14873_ _11910_/A _14871_/X _14872_/X VGND VGND VPWR VPWR _14873_/X sky130_fd_sc_hd__and3_4
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14696__A _14647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22119__A2 _22111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19400_ _19400_/A VGND VGND VPWR VPWR _19400_/Y sky130_fd_sc_hd__inv_2
X_16612_ _16646_/A _16609_/X _16611_/X VGND VGND VPWR VPWR _16612_/X sky130_fd_sc_hd__and3_4
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13824_ _15415_/A _13822_/X _13823_/X VGND VGND VPWR VPWR _13824_/X sky130_fd_sc_hd__and3_4
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17592_ _16821_/B _17913_/B _17271_/Y _17591_/X VGND VGND VPWR VPWR _17592_/X sky130_fd_sc_hd__o22a_4
XFILLER_141_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19331_ _19327_/Y _19330_/A _19327_/A _19330_/Y VGND VGND VPWR VPWR _19331_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16543_ _16534_/X _16621_/B VGND VGND VPWR VPWR _16543_/X sky130_fd_sc_hd__or2_4
X_13755_ _12650_/A _13753_/X _13755_/C VGND VGND VPWR VPWR _13756_/C sky130_fd_sc_hd__and3_4
XFILLER_44_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21878__B2 _21870_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ _13145_/A _12804_/B VGND VGND VPWR VPWR _12707_/C sky130_fd_sc_hd__or2_4
XFILLER_31_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19262_ _24306_/Q _19255_/B _19261_/Y VGND VGND VPWR VPWR _19262_/X sky130_fd_sc_hd__o21a_4
X_16474_ _16474_/A _16472_/X _16473_/X VGND VGND VPWR VPWR _16474_/X sky130_fd_sc_hd__and3_4
X_13686_ _12294_/A _13769_/B VGND VGND VPWR VPWR _13686_/X sky130_fd_sc_hd__or2_4
XANTENNA__22418__A _20377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18213_ _18020_/X _18211_/X _18065_/X _18212_/X VGND VGND VPWR VPWR _18213_/X sky130_fd_sc_hd__o22a_4
X_15425_ _15406_/A _15489_/B VGND VGND VPWR VPWR _15427_/B sky130_fd_sc_hd__or2_4
XANTENNA__21322__A _21322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12637_ _12974_/A _12514_/B VGND VGND VPWR VPWR _12637_/X sky130_fd_sc_hd__or2_4
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19193_ _19145_/X VGND VGND VPWR VPWR _19193_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12944__A _12944_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15320__A _15372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23996__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18144_ _18068_/X _18143_/X _20012_/A _18068_/X VGND VGND VPWR VPWR _24493_/D sky130_fd_sc_hd__a2bb2o_4
X_12568_ _12568_/A _12664_/B VGND VGND VPWR VPWR _12568_/X sky130_fd_sc_hd__or2_4
X_15356_ _15319_/A _23832_/Q VGND VGND VPWR VPWR _15357_/C sky130_fd_sc_hd__or2_4
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14307_ _14307_/A _14380_/B VGND VGND VPWR VPWR _14309_/B sky130_fd_sc_hd__or2_4
X_11519_ _11519_/A _11519_/B VGND VGND VPWR VPWR _11519_/X sky130_fd_sc_hd__or2_4
X_18075_ _17792_/X VGND VGND VPWR VPWR _18283_/A sky130_fd_sc_hd__buf_2
X_12499_ _12499_/A VGND VGND VPWR VPWR _12871_/A sky130_fd_sc_hd__buf_2
X_15287_ _14269_/A _24056_/Q VGND VGND VPWR VPWR _15288_/C sky130_fd_sc_hd__or2_4
XFILLER_144_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17026_ _17025_/Y VGND VGND VPWR VPWR _17026_/X sky130_fd_sc_hd__buf_2
XANTENNA__22055__B2 _22050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14238_ _15324_/A VGND VGND VPWR VPWR _14656_/A sky130_fd_sc_hd__buf_2
XANTENNA__22153__A _20859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13775__A _12623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17247__A _18320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14169_ _14169_/A _23711_/Q VGND VGND VPWR VPWR _14171_/B sky130_fd_sc_hd__or2_4
XANTENNA__16151__A _16116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21802__B2 _21767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_3_0_HCLK clkbuf_5_1_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_6_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_140_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21992__A _22007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18977_ _18963_/X _18975_/Y _18976_/Y _18968_/X VGND VGND VPWR VPWR _18977_/X sky130_fd_sc_hd__o22a_4
XFILLER_58_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20104__C _20098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17928_ _17825_/X _17178_/X _17814_/X _17206_/X VGND VGND VPWR VPWR _17928_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17859_ _17922_/A _17857_/X _17836_/X _17858_/X VGND VGND VPWR VPWR _17859_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18078__A _17801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20870_ _20864_/X _20866_/X _20867_/X HRDATA[14] _20869_/X VGND VGND VPWR VPWR _20870_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_82_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19529_ _19740_/A VGND VGND VPWR VPWR _19899_/B sky130_fd_sc_hd__buf_2
XFILLER_41_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__A2 _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13015__A _12461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22540_ _22555_/A VGND VGND VPWR VPWR _22548_/A sky130_fd_sc_hd__buf_2
X_22471_ _22471_/A VGND VGND VPWR VPWR _22471_/X sky130_fd_sc_hd__buf_2
XANTENNA__12854__A _12854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24210_ _23095_/CLK _19554_/X HRESETn VGND VGND VPWR VPWR _24210_/Q sky130_fd_sc_hd__dfrtp_4
X_21422_ _21455_/A VGND VGND VPWR VPWR _21438_/A sky130_fd_sc_hd__inv_2
X_24141_ _24137_/CLK _24141_/D HRESETn VGND VGND VPWR VPWR _24141_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21353_ _21287_/X _21348_/X _15552_/B _21352_/X VGND VGND VPWR VPWR _23905_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20304_ _20977_/A VGND VGND VPWR VPWR _20304_/X sky130_fd_sc_hd__buf_2
X_24072_ _24073_/CLK _24072_/D VGND VGND VPWR VPWR _24072_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_146_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21284_ _21283_/X _21281_/X _15865_/B _21276_/X VGND VGND VPWR VPWR _21284_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24151__CLK _24302_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13685__A _15446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23023_ _23007_/X _17681_/A _23019_/X _23022_/X VGND VGND VPWR VPWR _23024_/A sky130_fd_sc_hd__a211o_4
XANTENNA__22597__A2 _22594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20235_ _20234_/X VGND VGND VPWR VPWR _20235_/X sky130_fd_sc_hd__buf_2
XANTENNA__23719__CLK _23750_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20166_ IRQ[9] VGND VGND VPWR VPWR _20166_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20097_ NMI _20194_/A VGND VGND VPWR VPWR _20146_/A sky130_fd_sc_hd__or2_4
XFILLER_18_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23925_ _23392_/CLK _23925_/D VGND VGND VPWR VPWR _23925_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23869__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11933__A _11933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15405__A _15405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11870_ _15449_/A VGND VGND VPWR VPWR _12186_/A sky130_fd_sc_hd__buf_2
X_23856_ _24080_/CLK _23856_/D VGND VGND VPWR VPWR _16429_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22807_ _17327_/Y _22804_/X VGND VGND VPWR VPWR HWDATA[2] sky130_fd_sc_hd__nor2_4
XFILLER_77_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23787_ _23467_/CLK _21550_/X VGND VGND VPWR VPWR _23787_/Q sky130_fd_sc_hd__dfxtp_4
X_20999_ _20639_/A _20986_/X _20779_/X _20998_/Y VGND VGND VPWR VPWR _20999_/X sky130_fd_sc_hd__a211o_4
XFILLER_26_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13540_ _12949_/A VGND VGND VPWR VPWR _13540_/X sky130_fd_sc_hd__buf_2
XANTENNA__20532__A1 _20418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22738_ _22738_/A _22737_/X VGND VGND VPWR VPWR _23086_/C sky130_fd_sc_hd__and2_4
XANTENNA__20532__B2 _20510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13471_ _13467_/A _13471_/B _13471_/C VGND VGND VPWR VPWR _13475_/B sky130_fd_sc_hd__and3_4
XFILLER_164_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22669_ _22655_/A VGND VGND VPWR VPWR _22669_/X sky130_fd_sc_hd__buf_2
XFILLER_41_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12764__A _13562_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12422_ _12422_/A VGND VGND VPWR VPWR _12423_/B sky130_fd_sc_hd__inv_2
X_15210_ _15196_/X _15139_/B VGND VGND VPWR VPWR _15210_/X sky130_fd_sc_hd__or2_4
X_24408_ _24419_/CLK _18882_/X HRESETn VGND VGND VPWR VPWR _24408_/Q sky130_fd_sc_hd__dfrtp_4
X_16190_ _16210_/A _16190_/B _16189_/X VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__and3_4
XANTENNA__22285__B2 _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11576__A2 IRQ[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12353_ _13123_/A _12343_/X _12352_/X VGND VGND VPWR VPWR _12353_/X sky130_fd_sc_hd__and3_4
X_15141_ _13791_/A _15141_/B _15141_/C VGND VGND VPWR VPWR _15141_/X sky130_fd_sc_hd__and3_4
X_24339_ _24277_/CLK _19164_/X HRESETn VGND VGND VPWR VPWR _24339_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15072_ _15080_/A _23445_/Q VGND VGND VPWR VPWR _15073_/C sky130_fd_sc_hd__or2_4
X_12284_ _13276_/A _12281_/X _12283_/X VGND VGND VPWR VPWR _12284_/X sky130_fd_sc_hd__and3_4
XANTENNA__22037__B2 _22000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12525__A1 _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18900_ _18900_/A VGND VGND VPWR VPWR _18900_/X sky130_fd_sc_hd__buf_2
X_14023_ _11736_/A _14023_/B _14022_/X VGND VGND VPWR VPWR _14024_/C sky130_fd_sc_hd__and3_4
XFILLER_153_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19880_ _19819_/A _19878_/X _19859_/A _19879_/X VGND VGND VPWR VPWR _19880_/X sky130_fd_sc_hd__a211o_4
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17464__A1 _17046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18831_ _15118_/X _18796_/A _24438_/Q _18790_/A VGND VGND VPWR VPWR _24438_/D sky130_fd_sc_hd__o22a_4
XFILLER_96_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21260__A2 _21257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22701__A _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18762_ _17090_/X VGND VGND VPWR VPWR _18762_/Y sky130_fd_sc_hd__inv_2
X_15974_ _16011_/A _15972_/X _15973_/X VGND VGND VPWR VPWR _15978_/B sky130_fd_sc_hd__and3_4
XANTENNA__12004__A _12015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17713_ _16983_/A VGND VGND VPWR VPWR _18368_/A sky130_fd_sc_hd__buf_2
XFILLER_76_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14925_ _13694_/A VGND VGND VPWR VPWR _14925_/X sky130_fd_sc_hd__buf_2
X_18693_ _17801_/X _18693_/B VGND VGND VPWR VPWR _18693_/X sky130_fd_sc_hd__and2_4
X_17644_ _17915_/B _17643_/Y _17914_/B VGND VGND VPWR VPWR _17644_/X sky130_fd_sc_hd__o21a_4
X_14856_ _14096_/A _23190_/Q VGND VGND VPWR VPWR _14856_/X sky130_fd_sc_hd__or2_4
XANTENNA__20771__A1 _20635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20771__B2 _20746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11562__B IRQ[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13807_ _14311_/A _13807_/B VGND VGND VPWR VPWR _13809_/B sky130_fd_sc_hd__or2_4
X_17575_ _11608_/X _17251_/B VGND VGND VPWR VPWR _17575_/X sky130_fd_sc_hd__and2_4
XFILLER_56_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14787_ _15103_/A _14713_/B VGND VGND VPWR VPWR _14787_/X sky130_fd_sc_hd__or2_4
X_11999_ _12108_/A _11999_/B _11999_/C VGND VGND VPWR VPWR _11999_/X sky130_fd_sc_hd__or3_4
X_19314_ _24280_/Q _19228_/X _19313_/Y VGND VGND VPWR VPWR _19314_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17530__A _13567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16526_ _16526_/A _16525_/Y VGND VGND VPWR VPWR _16527_/B sky130_fd_sc_hd__or2_4
X_13738_ _15502_/A _13738_/B VGND VGND VPWR VPWR _13739_/C sky130_fd_sc_hd__or2_4
XFILLER_43_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21052__A _21045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19245_ _24296_/Q _19245_/B VGND VGND VPWR VPWR _19246_/B sky130_fd_sc_hd__and2_4
XFILLER_91_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16457_ _11714_/A VGND VGND VPWR VPWR _16490_/A sky130_fd_sc_hd__buf_2
XFILLER_31_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12674__A _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13669_ _15408_/A _13667_/X _13669_/C VGND VGND VPWR VPWR _13669_/X sky130_fd_sc_hd__and3_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15050__A _12322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15408_ _15408_/A _15408_/B _15408_/C VGND VGND VPWR VPWR _15412_/B sky130_fd_sc_hd__and3_4
XANTENNA__21079__A2 _21045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19176_ _19154_/A _19154_/B _19175_/Y VGND VGND VPWR VPWR _19176_/X sky130_fd_sc_hd__o21a_4
X_16388_ _15959_/A _16388_/B VGND VGND VPWR VPWR _16389_/C sky130_fd_sc_hd__or2_4
XANTENNA__20891__A _22471_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24174__CLK _23383_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18127_ _18126_/A _17938_/X _18126_/A _17935_/Y VGND VGND VPWR VPWR _18127_/X sky130_fd_sc_hd__a2bb2o_4
X_15339_ _15326_/A _23672_/Q VGND VGND VPWR VPWR _15339_/X sky130_fd_sc_hd__or2_4
XFILLER_172_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18058_ _18389_/A _18004_/X _18389_/A _18001_/X VGND VGND VPWR VPWR _18059_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17009_ _17009_/A _17009_/B _17008_/Y VGND VGND VPWR VPWR _17010_/B sky130_fd_sc_hd__and3_4
XFILLER_99_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_92_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR _24090_/CLK sky130_fd_sc_hd__clkbuf_1
X_20020_ _20016_/X _17675_/A _19998_/X _20019_/X VGND VGND VPWR VPWR _20020_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17455__A1 _17046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22200__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21971_ _21957_/A VGND VGND VPWR VPWR _21971_/X sky130_fd_sc_hd__buf_2
XFILLER_6_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13952__B _23264_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11753__A _11753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23710_ _23646_/CLK _21693_/X VGND VGND VPWR VPWR _13768_/B sky130_fd_sc_hd__dfxtp_4
X_20922_ _24409_/Q _20316_/X VGND VGND VPWR VPWR _20922_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12568__B _12664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853_ _21017_/A _20852_/X VGND VGND VPWR VPWR _20853_/Y sky130_fd_sc_hd__nor2_4
X_23641_ _23641_/CLK _23641_/D VGND VGND VPWR VPWR _14754_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22503__A2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23572_ _23668_/CLK _21944_/X VGND VGND VPWR VPWR _21937_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20784_ _11567_/A VGND VGND VPWR VPWR _20785_/A sky130_fd_sc_hd__inv_2
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24494__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22523_ _22461_/X _22522_/X _23231_/Q _22519_/X VGND VGND VPWR VPWR _23231_/D sky130_fd_sc_hd__o22a_4
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12584__A _12949_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16056__A _16056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22454_ _20718_/A VGND VGND VPWR VPWR _22454_/X sky130_fd_sc_hd__buf_2
XANTENNA__22267__B2 _22262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21405_ _21405_/A VGND VGND VPWR VPWR _21405_/X sky130_fd_sc_hd__buf_2
XANTENNA__15895__A _13529_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22385_ _22137_/X _22383_/X _15800_/B _22380_/X VGND VGND VPWR VPWR _23299_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17143__B1 _16242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24124_ _23416_/CLK _22793_/X HRESETn VGND VGND VPWR VPWR _22763_/A sky130_fd_sc_hd__dfrtp_4
X_21336_ _21259_/X _21334_/X _16132_/B _21331_/X VGND VGND VPWR VPWR _21336_/X sky130_fd_sc_hd__o22a_4
XFILLER_159_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22019__B2 _22014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21490__A2 _21485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20306__A _20234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24055_ _23544_/CLK _21077_/X VGND VGND VPWR VPWR _15223_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__11928__A _11928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21267_ _21266_/X _21257_/X _12789_/B _21264_/X VGND VGND VPWR VPWR _23946_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14304__A _14304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23006_ _23006_/A VGND VGND VPWR VPWR HADDR[17] sky130_fd_sc_hd__inv_2
X_20218_ _20218_/A _20218_/B _20217_/X VGND VGND VPWR VPWR _21234_/B sky130_fd_sc_hd__or3_4
XFILLER_131_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18643__B1 _18638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21198_ _21198_/A VGND VGND VPWR VPWR _21198_/X sky130_fd_sc_hd__buf_2
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20149_ _18623_/Y _18705_/X _20148_/X VGND VGND VPWR VPWR _20149_/X sky130_fd_sc_hd__o21a_4
XFILLER_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21137__A _21152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12971_ _12971_/A _24105_/Q VGND VGND VPWR VPWR _12971_/X sky130_fd_sc_hd__or2_4
XFILLER_79_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15135__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14710_ _12484_/A _14780_/B VGND VGND VPWR VPWR _14710_/X sky130_fd_sc_hd__or2_4
XFILLER_131_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23908_ _23908_/CLK _21349_/X VGND VGND VPWR VPWR _23908_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11922_ _11975_/A VGND VGND VPWR VPWR _16741_/A sky130_fd_sc_hd__buf_2
XFILLER_131_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15690_ _13300_/A _15755_/B VGND VGND VPWR VPWR _15690_/X sky130_fd_sc_hd__or2_4
XFILLER_45_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14641_ _14840_/A _14641_/B _14641_/C VGND VGND VPWR VPWR _14642_/C sky130_fd_sc_hd__or3_4
X_11853_ _11853_/A VGND VGND VPWR VPWR _11854_/A sky130_fd_sc_hd__buf_2
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23839_ _23294_/CLK _23839_/D VGND VGND VPWR VPWR _23839_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _17360_/A _17360_/B VGND VGND VPWR VPWR _17360_/X sky130_fd_sc_hd__or2_4
XANTENNA__15789__B _15789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11784_ _13400_/A VGND VGND VPWR VPWR _11784_/X sky130_fd_sc_hd__buf_2
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14572_ _15401_/A _14572_/B _14571_/X VGND VGND VPWR VPWR _14573_/C sky130_fd_sc_hd__and3_4
XPHY_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24197__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ _16192_/A _16247_/B VGND VGND VPWR VPWR _16313_/B sky130_fd_sc_hd__or2_4
XPHY_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ _13535_/A _24005_/Q VGND VGND VPWR VPWR _13524_/C sky130_fd_sc_hd__or2_4
X_17291_ _17290_/X _17292_/B VGND VGND VPWR VPWR _18651_/B sky130_fd_sc_hd__and2_4
XFILLER_159_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17382__B1 _17028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12494__A _12188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19030_ _19030_/A VGND VGND VPWR VPWR _19030_/Y sky130_fd_sc_hd__inv_2
X_16242_ _16243_/B VGND VGND VPWR VPWR _16242_/X sky130_fd_sc_hd__buf_2
X_13454_ _11865_/X _13425_/X _13434_/X _13445_/X _13453_/X VGND VGND VPWR VPWR _13454_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12405_ _12402_/X _12405_/B _12405_/C VGND VGND VPWR VPWR _12406_/C sky130_fd_sc_hd__and3_4
XFILLER_166_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13385_ _13385_/A _23974_/Q VGND VGND VPWR VPWR _13386_/C sky130_fd_sc_hd__or2_4
X_16173_ _16216_/A _16102_/B VGND VGND VPWR VPWR _16173_/X sky130_fd_sc_hd__or2_4
XFILLER_154_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17134__B1 _17132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19674__A2 _19673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15124_ _12426_/A _15122_/X _15123_/X VGND VGND VPWR VPWR _15128_/B sky130_fd_sc_hd__and3_4
XANTENNA__21481__A2 _21478_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12336_ _12336_/A VGND VGND VPWR VPWR _12337_/A sky130_fd_sc_hd__buf_2
XFILLER_114_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_16_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_16_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12267_ _13042_/A VGND VGND VPWR VPWR _12689_/A sky130_fd_sc_hd__buf_2
X_19932_ _22745_/A VGND VGND VPWR VPWR _19932_/X sky130_fd_sc_hd__buf_2
X_15055_ _15076_/A VGND VGND VPWR VPWR _15086_/A sky130_fd_sc_hd__buf_2
X_14006_ _12501_/A _14068_/B VGND VGND VPWR VPWR _14007_/C sky130_fd_sc_hd__or2_4
X_19863_ _19863_/A VGND VGND VPWR VPWR _21319_/A sky130_fd_sc_hd__buf_2
X_12198_ _12198_/A VGND VGND VPWR VPWR _12512_/A sky130_fd_sc_hd__buf_2
XFILLER_122_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18814_ _15916_/X _18810_/X _24451_/Q _18811_/X VGND VGND VPWR VPWR _18814_/X sky130_fd_sc_hd__o22a_4
X_19794_ _19742_/A _19613_/X _19662_/X VGND VGND VPWR VPWR _19803_/B sky130_fd_sc_hd__o21a_4
XFILLER_23_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18745_ _12024_/A _17075_/X VGND VGND VPWR VPWR _18745_/X sky130_fd_sc_hd__or2_4
X_15957_ _15957_/A _24046_/Q VGND VGND VPWR VPWR _15961_/B sky130_fd_sc_hd__or2_4
XFILLER_114_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12669__A _12943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18937__A1 _17290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22733__A2 _22729_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11573__A _11573_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14908_ _11928_/A _14904_/X _14907_/X VGND VGND VPWR VPWR _14908_/X sky130_fd_sc_hd__or3_4
X_18676_ _18198_/A _17998_/X VGND VGND VPWR VPWR _18676_/Y sky130_fd_sc_hd__nor2_4
X_15888_ _13531_/A _15826_/B VGND VGND VPWR VPWR _15890_/B sky130_fd_sc_hd__or2_4
XFILLER_23_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20886__A _20885_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17627_ _17624_/Y _17626_/Y _17341_/B VGND VGND VPWR VPWR _17627_/X sky130_fd_sc_hd__o21a_4
X_14839_ _14647_/X _14839_/B _14839_/C VGND VGND VPWR VPWR _14839_/X sky130_fd_sc_hd__and3_4
XFILLER_52_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18356__A _18019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17558_ _17047_/A _17557_/X _17050_/X VGND VGND VPWR VPWR _17558_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22497__B2 _22491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16509_ _16166_/X _16446_/B VGND VGND VPWR VPWR _16510_/C sky130_fd_sc_hd__or2_4
XANTENNA__12985__A1 _12914_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17489_ _17600_/D VGND VGND VPWR VPWR _17490_/D sky130_fd_sc_hd__inv_2
X_19228_ _19228_/A _19227_/X VGND VGND VPWR VPWR _19228_/X sky130_fd_sc_hd__and2_4
XANTENNA__22249__B2 _22248_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21510__A _21489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19159_ _19159_/A _19159_/B VGND VGND VPWR VPWR _19160_/B sky130_fd_sc_hd__and2_4
XANTENNA__16604__A _11686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22170_ _22169_/X _22123_/A _23445_/Q _22106_/A VGND VGND VPWR VPWR _23445_/D sky130_fd_sc_hd__o22a_4
XFILLER_133_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21121_ _20841_/X _21118_/X _24029_/Q _21115_/X VGND VGND VPWR VPWR _21121_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19915__A _18774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14124__A _13981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17428__A1 _17425_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21052_ _21045_/A VGND VGND VPWR VPWR _21052_/X sky130_fd_sc_hd__buf_2
XFILLER_132_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17428__B2 _17427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20003_ _20003_/A VGND VGND VPWR VPWR _20003_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13963__A _13990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13682__B _13765_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12579__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22724__A2 _22722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21954_ _21826_/X _21953_/X _23566_/Q _21950_/X VGND VGND VPWR VPWR _21954_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ _20425_/A _20904_/X _19231_/A _20758_/X VGND VGND VPWR VPWR _20905_/X sky130_fd_sc_hd__o22a_4
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21885_ _21024_/A VGND VGND VPWR VPWR _21885_/X sky130_fd_sc_hd__buf_2
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14794__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17170__A _17169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23624_ _24073_/CLK _21842_/X VGND VGND VPWR VPWR _23624_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20639_/A _20824_/X _20779_/X _20835_/Y VGND VGND VPWR VPWR _20836_/X sky130_fd_sc_hd__a211o_4
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23555_ _23650_/CLK _23555_/D VGND VGND VPWR VPWR _15807_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15402__B _15465_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20767_ _20857_/A _20767_/B VGND VGND VPWR VPWR _20767_/Y sky130_fd_sc_hd__nand2_4
XFILLER_39_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21160__B2 _21159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__A _13251_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22506_ _22432_/X _22501_/X _12671_/B _22505_/X VGND VGND VPWR VPWR _22506_/X sky130_fd_sc_hd__o22a_4
XFILLER_156_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23486_ _23997_/CLK _22076_/X VGND VGND VPWR VPWR _13772_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_168_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20698_ HRDATA[13] _20697_/X VGND VGND VPWR VPWR _20700_/B sky130_fd_sc_hd__or2_4
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14018__B _23264_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22437_ _20558_/A VGND VGND VPWR VPWR _22437_/X sky130_fd_sc_hd__buf_2
XFILLER_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13170_ _13170_/A _13170_/B _13169_/X VGND VGND VPWR VPWR _13170_/X sky130_fd_sc_hd__and3_4
XFILLER_136_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22368_ _22108_/X _22362_/X _16260_/B _22366_/X VGND VGND VPWR VPWR _22368_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21463__A2 _21462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22660__B2 _22655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12121_ _12164_/A _23763_/Q VGND VGND VPWR VPWR _12121_/X sky130_fd_sc_hd__or2_4
X_24107_ _23558_/CLK _20511_/X VGND VGND VPWR VPWR _12669_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__11658__A _14772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21319_ _21319_/A VGND VGND VPWR VPWR _21320_/C sky130_fd_sc_hd__buf_2
X_22299_ _22129_/X _22294_/X _23366_/Q _22298_/X VGND VGND VPWR VPWR _22299_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14034__A _11680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24038_ _24102_/CLK _21109_/X VGND VGND VPWR VPWR _13286_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21215__A2 _21212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12052_ _12041_/A _12128_/B VGND VGND VPWR VPWR _12052_/X sky130_fd_sc_hd__or2_4
XFILLER_172_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17419__B2 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22251__A _22244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20423__B1 _20235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16860_ _15656_/X _16842_/X _15656_/X _16842_/X VGND VGND VPWR VPWR _16860_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20974__A1 _18717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15811_ _12854_/A _15866_/B VGND VGND VPWR VPWR _15811_/X sky130_fd_sc_hd__or2_4
X_16791_ _16791_/A _23633_/Q VGND VGND VPWR VPWR _16791_/X sky130_fd_sc_hd__or2_4
XANTENNA__12489__A _12869_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18919__A1 _17172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18530_ _18499_/X _18526_/X _18527_/X _18529_/X VGND VGND VPWR VPWR _18530_/X sky130_fd_sc_hd__o22a_4
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15742_ _15741_/X _23684_/Q VGND VGND VPWR VPWR _15742_/X sky130_fd_sc_hd__or2_4
X_12954_ _12954_/A _12950_/X _12954_/C VGND VGND VPWR VPWR _12962_/B sky130_fd_sc_hd__or3_4
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11905_ _11904_/X VGND VGND VPWR VPWR _11905_/X sky130_fd_sc_hd__buf_2
XANTENNA__23082__A _23081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18461_ _18461_/A _17375_/A VGND VGND VPWR VPWR _18462_/D sky130_fd_sc_hd__and2_4
X_15673_ _13170_/A _15673_/B _15672_/X VGND VGND VPWR VPWR _15677_/B sky130_fd_sc_hd__and3_4
XFILLER_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12885_ _12885_/A _23977_/Q VGND VGND VPWR VPWR _12886_/C sky130_fd_sc_hd__or2_4
XFILLER_46_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_7_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17412_ _17412_/A _17412_/B VGND VGND VPWR VPWR _17412_/X sky130_fd_sc_hd__and2_4
X_14624_ _14834_/A _23354_/Q VGND VGND VPWR VPWR _14624_/X sky130_fd_sc_hd__or2_4
X_11836_ _11836_/A _23892_/Q VGND VGND VPWR VPWR _11837_/C sky130_fd_sc_hd__or2_4
XANTENNA__22479__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18392_ _17499_/Y _18391_/X VGND VGND VPWR VPWR _18392_/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17343_ _11592_/X _17357_/B _17414_/A _12891_/A _17342_/Y VGND VGND VPWR VPWR _17343_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14555_ _12427_/A _14553_/X _14554_/X VGND VGND VPWR VPWR _14555_/X sky130_fd_sc_hd__and3_4
XPHY_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11767_ _16031_/A VGND VGND VPWR VPWR _16048_/A sky130_fd_sc_hd__buf_2
XANTENNA__21151__B2 _21145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13506_ _12644_/A VGND VGND VPWR VPWR _13535_/A sky130_fd_sc_hd__buf_2
XFILLER_158_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17274_ _17274_/A VGND VGND VPWR VPWR _17276_/A sky130_fd_sc_hd__inv_2
X_14486_ _12410_/A _14484_/X _14485_/X VGND VGND VPWR VPWR _14490_/B sky130_fd_sc_hd__and3_4
XANTENNA__22426__A _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11698_ _11698_/A VGND VGND VPWR VPWR _12604_/A sky130_fd_sc_hd__buf_2
X_19013_ _24394_/Q VGND VGND VPWR VPWR _19013_/Y sky130_fd_sc_hd__inv_2
X_16225_ _16185_/A _16223_/X _16224_/X VGND VGND VPWR VPWR _16229_/B sky130_fd_sc_hd__and3_4
X_13437_ _13431_/X _24005_/Q VGND VGND VPWR VPWR _13438_/C sky130_fd_sc_hd__or2_4
XFILLER_158_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16156_ _16156_/A _16226_/B VGND VGND VPWR VPWR _16158_/B sky130_fd_sc_hd__or2_4
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21454__A2 _21448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13368_ _13387_/A VGND VGND VPWR VPWR _13378_/A sky130_fd_sc_hd__buf_2
XANTENNA__12671__B _12671_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15107_ _15095_/A _23477_/Q VGND VGND VPWR VPWR _15107_/X sky130_fd_sc_hd__or2_4
X_12319_ _11856_/A _11630_/A _12263_/X _12264_/X _12318_/X VGND VGND VPWR VPWR _12320_/A
+ sky130_fd_sc_hd__a32o_4
X_16087_ _16016_/Y _16085_/X VGND VGND VPWR VPWR _16088_/A sky130_fd_sc_hd__or2_4
X_13299_ _12516_/A _13295_/X _13299_/C VGND VGND VPWR VPWR _13299_/X sky130_fd_sc_hd__or3_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24212__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21206__A2 _21205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19915_ _18774_/X VGND VGND VPWR VPWR _19915_/X sky130_fd_sc_hd__buf_2
X_15038_ _13606_/A _15038_/B VGND VGND VPWR VPWR _15039_/C sky130_fd_sc_hd__or2_4
XFILLER_102_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22403__B2 _22366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22161__A _20937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13783__A _13692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19846_ _21603_/A VGND VGND VPWR VPWR _21134_/A sky130_fd_sc_hd__buf_2
XFILLER_68_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17830__A1 _17813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16989_ _16989_/A _16989_/B VGND VGND VPWR VPWR _18189_/A sky130_fd_sc_hd__or2_4
X_19777_ _19777_/A VGND VGND VPWR VPWR _19777_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24362__CLK _24357_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22706__A2 _22701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18728_ _17108_/X _17346_/B VGND VGND VPWR VPWR _18731_/A sky130_fd_sc_hd__or2_4
XANTENNA__20717__A1 _24226_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18659_ _16973_/X VGND VGND VPWR VPWR _18661_/A sky130_fd_sc_hd__inv_2
XFILLER_97_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17702__B _17473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21390__B2 _21388_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21670_ _21677_/A VGND VGND VPWR VPWR _21670_/X sky130_fd_sc_hd__buf_2
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20621_ _20620_/X VGND VGND VPWR VPWR _20621_/Y sky130_fd_sc_hd__inv_2
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21142__B2 _21138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13023__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23340_ _23204_/CLK _23340_/D VGND VGND VPWR VPWR _12374_/B sky130_fd_sc_hd__dfxtp_4
X_20552_ _18272_/X _20446_/X _20538_/X _20551_/Y VGND VGND VPWR VPWR _20552_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17897__A1 _16935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21693__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22890__A1 _16452_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21240__A _21239_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23271_ _24039_/CLK _23271_/D VGND VGND VPWR VPWR _23271_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20483_ _20438_/A _20482_/X VGND VGND VPWR VPWR _20483_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__16334__A _11727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22222_ _11827_/B VGND VGND VPWR VPWR _22222_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24343__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22642__B2 _22641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22153_ _20859_/A VGND VGND VPWR VPWR _22153_/X sky130_fd_sc_hd__buf_2
XFILLER_160_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21104_ _21104_/A VGND VGND VPWR VPWR _21104_/X sky130_fd_sc_hd__buf_2
X_22084_ _21879_/X _22081_/X _23480_/Q _22078_/X VGND VGND VPWR VPWR _22084_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22071__A _22057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14789__A _15081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_62_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21035_ _21042_/A VGND VGND VPWR VPWR _21035_/X sky130_fd_sc_hd__buf_2
XANTENNA__13693__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17165__A _13266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17821__A1 _17816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22986_ _22978_/X _22986_/B _22986_/C VGND VGND VPWR VPWR _22986_/X sky130_fd_sc_hd__and3_4
XFILLER_167_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21937_ _21937_/A VGND VGND VPWR VPWR _21937_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11941__A _11941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15413__A _14325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12670_ _12670_/A _12668_/X _12669_/X VGND VGND VPWR VPWR _12674_/B sky130_fd_sc_hd__and3_4
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21868_ _21867_/X _21863_/X _23613_/Q _21858_/X VGND VGND VPWR VPWR _23613_/D sky130_fd_sc_hd__o22a_4
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ _23864_/CLK _23607_/D VGND VGND VPWR VPWR _15222_/B sky130_fd_sc_hd__dfxtp_4
X_11621_ _12473_/A VGND VGND VPWR VPWR _12188_/A sky130_fd_sc_hd__buf_2
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20819_ _20819_/A VGND VGND VPWR VPWR _20819_/X sky130_fd_sc_hd__buf_2
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21799_ _21589_/X _21798_/X _14601_/B _21795_/X VGND VGND VPWR VPWR _23642_/D sky130_fd_sc_hd__o22a_4
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ _12410_/A _14340_/B _14340_/C VGND VGND VPWR VPWR _14340_/X sky130_fd_sc_hd__and3_4
X_23538_ _23537_/CLK _23538_/D VGND VGND VPWR VPWR _23538_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ _24439_/Q IRQ[2] VGND VGND VPWR VPWR _11552_/Y sky130_fd_sc_hd__nand2_4
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14271_ _12427_/A _14271_/B _14271_/C VGND VGND VPWR VPWR _14271_/X sky130_fd_sc_hd__and3_4
X_23469_ _23501_/CLK _23469_/D VGND VGND VPWR VPWR _16196_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12772__A _12976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16010_ _16009_/X _16010_/B VGND VGND VPWR VPWR _16011_/C sky130_fd_sc_hd__or2_4
X_13222_ _13253_/A _24007_/Q VGND VGND VPWR VPWR _13223_/C sky130_fd_sc_hd__or2_4
XFILLER_171_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21436__A2 _21434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22633__B2 _22598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13153_ _12702_/A _23591_/Q VGND VGND VPWR VPWR _13154_/C sky130_fd_sc_hd__or2_4
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12104_ _11951_/X _12104_/B _12103_/X VGND VGND VPWR VPWR _12104_/X sky130_fd_sc_hd__and3_4
X_13084_ _13097_/A _23688_/Q VGND VGND VPWR VPWR _13086_/B sky130_fd_sc_hd__or2_4
XANTENNA__23077__A _23076_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17961_ _16935_/X _17958_/X _17653_/X _17960_/X VGND VGND VPWR VPWR _17961_/X sky130_fd_sc_hd__o22a_4
XFILLER_97_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14699__A _15649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12035_ _16691_/A _23539_/Q VGND VGND VPWR VPWR _12036_/C sky130_fd_sc_hd__or2_4
X_19700_ _19700_/A VGND VGND VPWR VPWR _19700_/X sky130_fd_sc_hd__buf_2
X_16912_ _16911_/X VGND VGND VPWR VPWR _16912_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17892_ _17791_/X _17804_/Y _17886_/X _17888_/Y _17891_/X VGND VGND VPWR VPWR _17892_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20213__B _22039_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20947__B2 _20282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19631_ _19589_/X _19619_/A _19596_/X VGND VGND VPWR VPWR _19631_/X sky130_fd_sc_hd__o21a_4
X_16843_ _15656_/X _16842_/X _15654_/X VGND VGND VPWR VPWR _16843_/X sky130_fd_sc_hd__o21a_4
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14211__B _23455_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13108__A _12962_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19562_ _19849_/B _19649_/A VGND VGND VPWR VPWR _19562_/X sky130_fd_sc_hd__or2_4
XANTENNA__17803__A _17793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16774_ _16791_/A _16774_/B VGND VGND VPWR VPWR _16774_/X sky130_fd_sc_hd__or2_4
X_13986_ _13642_/A _23616_/Q VGND VGND VPWR VPWR _13988_/B sky130_fd_sc_hd__or2_4
XFILLER_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18513_ _17436_/C _18512_/X VGND VGND VPWR VPWR _18513_/Y sky130_fd_sc_hd__nand2_4
X_15725_ _13091_/A _15721_/X _15724_/X VGND VGND VPWR VPWR _15733_/B sky130_fd_sc_hd__or3_4
X_12937_ _12975_/A _12937_/B _12936_/X VGND VGND VPWR VPWR _12937_/X sky130_fd_sc_hd__and3_4
X_19493_ _19493_/A VGND VGND VPWR VPWR _19705_/B sky130_fd_sc_hd__buf_2
XANTENNA__17522__B _17522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12947__A _12641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16419__A _11971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11851__A _11671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18444_ _18198_/X _18343_/B _18265_/X _18443_/X VGND VGND VPWR VPWR _18444_/X sky130_fd_sc_hd__a211o_4
XFILLER_61_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15656_ _15582_/X _15653_/X _15655_/Y VGND VGND VPWR VPWR _15656_/X sky130_fd_sc_hd__a21o_4
X_12868_ _12868_/A _24009_/Q VGND VGND VPWR VPWR _12869_/C sky130_fd_sc_hd__or2_4
XFILLER_61_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14607_ _13652_/A _14686_/B VGND VGND VPWR VPWR _14607_/X sky130_fd_sc_hd__or2_4
X_11819_ _11762_/X _11817_/X _11818_/X VGND VGND VPWR VPWR _11819_/X sky130_fd_sc_hd__and3_4
X_18375_ _18483_/A _18290_/A VGND VGND VPWR VPWR _18375_/X sky130_fd_sc_hd__or2_4
X_15587_ _15610_/A _15525_/B VGND VGND VPWR VPWR _15587_/X sky130_fd_sc_hd__or2_4
X_12799_ _13563_/A _12791_/X _12798_/X VGND VGND VPWR VPWR _12799_/X sky130_fd_sc_hd__or3_4
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21124__B2 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22321__B1 _23349_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17326_ _17324_/X _17326_/B VGND VGND VPWR VPWR _18689_/A sky130_fd_sc_hd__and2_4
XANTENNA__21675__A2 _21670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14538_ _14519_/A _23483_/Q VGND VGND VPWR VPWR _14540_/B sky130_fd_sc_hd__or2_4
XANTENNA__22872__A1 _17273_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_2_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_2_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22156__A _22471_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14881__B _23958_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17343__A3 _17414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17257_ _17255_/X _17256_/B VGND VGND VPWR VPWR _17258_/A sky130_fd_sc_hd__or2_4
X_14469_ _12498_/A _14469_/B VGND VGND VPWR VPWR _14469_/X sky130_fd_sc_hd__or2_4
XFILLER_31_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16208_ _16215_/A _16132_/B VGND VGND VPWR VPWR _16208_/X sky130_fd_sc_hd__or2_4
XFILLER_174_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21995__A _21991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17188_ _17188_/A _17187_/X VGND VGND VPWR VPWR _17236_/B sky130_fd_sc_hd__or2_4
XANTENNA__22624__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23602__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16139_ _16108_/A _16139_/B VGND VGND VPWR VPWR _16139_/X sky130_fd_sc_hd__or2_4
XFILLER_102_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19829_ _19732_/X _19822_/X _19828_/X _18780_/X _19512_/X VGND VGND VPWR VPWR _24193_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14121__B _23551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13018__A _12878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22840_ _20700_/A _14483_/Y VGND VGND VPWR VPWR _22840_/X sky130_fd_sc_hd__or2_4
XFILLER_83_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13960__B _23200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22771_ SYSTICKCLKDIV[0] _22749_/Y _22770_/Y VGND VGND VPWR VPWR _24117_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21363__A1 _21304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12857__A _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21363__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15233__A _14663_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21722_ _21544_/X _21720_/X _16199_/B _21717_/X VGND VGND VPWR VPWR _21722_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21653_ _21598_/X _21648_/X _23734_/Q _21617_/A VGND VGND VPWR VPWR _23734_/D sky130_fd_sc_hd__o22a_4
X_24441_ _24445_/CLK _24441_/D HRESETn VGND VGND VPWR VPWR _20923_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24258__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20604_ _20516_/X _20603_/X _24358_/Q _20475_/X VGND VGND VPWR VPWR _20604_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21666__A2 _21663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21584_ _20860_/A VGND VGND VPWR VPWR _21584_/X sky130_fd_sc_hd__buf_2
XFILLER_21_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22863__A1 _14767_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24372_ _24397_/CLK _24372_/D HRESETn VGND VGND VPWR VPWR _11544_/C sky130_fd_sc_hd__dfstp_4
XFILLER_149_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14791__B _14717_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23323_ _23323_/CLK _23323_/D VGND VGND VPWR VPWR _23323_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13688__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20535_ _18597_/Y VGND VGND VPWR VPWR _20535_/X sky130_fd_sc_hd__buf_2
XANTENNA__20874__B1 _20866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21418__A2 _21391_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20466_ _20231_/A VGND VGND VPWR VPWR _20466_/X sky130_fd_sc_hd__buf_2
X_23254_ _23192_/CLK _23254_/D VGND VGND VPWR VPWR _14912_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23282__CLK _23537_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20626__B1 _20538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22205_ _22176_/A VGND VGND VPWR VPWR _22205_/X sky130_fd_sc_hd__buf_2
X_23185_ _23281_/CLK _23185_/D VGND VGND VPWR VPWR _16774_/B sky130_fd_sc_hd__dfxtp_4
X_20397_ _20302_/X _20395_/X _16436_/B _20396_/X VGND VGND VPWR VPWR _24112_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19492__B1 HRDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22136_ _22134_/X _22135_/X _15682_/B _22130_/X VGND VGND VPWR VPWR _23460_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11936__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22067_ _22060_/A VGND VGND VPWR VPWR _22067_/X sky130_fd_sc_hd__buf_2
XFILLER_102_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14312__A _12485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21018_ _18774_/X _20342_/X _20662_/X _21017_/Y VGND VGND VPWR VPWR _21018_/X sky130_fd_sc_hd__a211o_4
XFILLER_48_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14031__B _23296_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13840_ _15404_/A _13838_/X _13840_/C VGND VGND VPWR VPWR _13844_/B sky130_fd_sc_hd__and3_4
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18438__B _17448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21145__A _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13771_ _12578_/A _13767_/X _13770_/X VGND VGND VPWR VPWR _13771_/X sky130_fd_sc_hd__or3_4
XANTENNA__12767__A _12766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22969_ _22946_/X _18500_/A _22959_/X _22968_/X VGND VGND VPWR VPWR _22969_/X sky130_fd_sc_hd__a211o_4
XFILLER_56_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16239__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21354__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11671__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15510_ _12635_/A _15508_/X _15509_/X VGND VGND VPWR VPWR _15510_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_69_0_HCLK clkbuf_6_34_0_HCLK/X VGND VGND VPWR VPWR _24184_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15143__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12722_ _12722_/A _12720_/X _12721_/X VGND VGND VPWR VPWR _12722_/X sky130_fd_sc_hd__and3_4
X_16490_ _16490_/A _16421_/B VGND VGND VPWR VPWR _16490_/X sky130_fd_sc_hd__or2_4
XFILLER_31_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15441_ _12300_/A _15439_/X _15441_/C VGND VGND VPWR VPWR _15441_/X sky130_fd_sc_hd__and3_4
X_12653_ _12941_/A _12651_/X _12653_/C VGND VGND VPWR VPWR _12653_/X sky130_fd_sc_hd__and3_4
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14982__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21106__B2 _21101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18160_ _17833_/X _18158_/X _17811_/X _18159_/X VGND VGND VPWR VPWR _18160_/Y sky130_fd_sc_hd__a22oi_4
X_11604_ _11604_/A VGND VGND VPWR VPWR _11605_/A sky130_fd_sc_hd__buf_2
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22854__A1 _15117_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15372_ _15372_/A _15372_/B _15372_/C VGND VGND VPWR VPWR _15376_/B sky130_fd_sc_hd__and3_4
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12949_/A _12584_/B VGND VGND VPWR VPWR _12585_/C sky130_fd_sc_hd__or2_4
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17111_ _18198_/A VGND VGND VPWR VPWR _17111_/X sky130_fd_sc_hd__buf_2
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _11879_/A _14321_/X _14323_/C VGND VGND VPWR VPWR _14323_/X sky130_fd_sc_hd__and3_4
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11535_ _11535_/A _19018_/A VGND VGND VPWR VPWR _11535_/X sky130_fd_sc_hd__or2_4
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18091_ _17875_/X _18090_/X _17883_/X VGND VGND VPWR VPWR _18091_/Y sky130_fd_sc_hd__o21ai_4
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17042_ _17297_/A VGND VGND VPWR VPWR _17043_/A sky130_fd_sc_hd__inv_2
XFILLER_7_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14254_ _14254_/A _23231_/Q VGND VGND VPWR VPWR _14254_/X sky130_fd_sc_hd__or2_4
XANTENNA__22606__B2 _22605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13205_ _13205_/A _23783_/Q VGND VGND VPWR VPWR _13205_/X sky130_fd_sc_hd__or2_4
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19483__B1 HRDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14185_ _14616_/A _14185_/B _14184_/X VGND VGND VPWR VPWR _14192_/B sky130_fd_sc_hd__and3_4
XANTENNA__22082__A2 _22081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16702__A _16702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12007__A _12105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13136_ _12722_/A _13134_/X _13135_/X VGND VGND VPWR VPWR _13136_/X sky130_fd_sc_hd__and3_4
XFILLER_174_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20224__A _20510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18993_ _18959_/A VGND VGND VPWR VPWR _18993_/X sky130_fd_sc_hd__buf_2
XFILLER_155_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14847__A1 _14767_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11846__A _11836_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13067_ _13067_/A VGND VGND VPWR VPWR _13097_/A sky130_fd_sc_hd__buf_2
X_17944_ _17869_/X VGND VGND VPWR VPWR _17944_/X sky130_fd_sc_hd__buf_2
XANTENNA__14222__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19786__A1 _19788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12018_ _11867_/X _12018_/B VGND VGND VPWR VPWR _12018_/X sky130_fd_sc_hd__and2_4
XFILLER_66_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11565__B IRQ[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17875_ _17874_/X VGND VGND VPWR VPWR _17875_/X sky130_fd_sc_hd__buf_2
XFILLER_93_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21593__B2 _21585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19614_ _19613_/X _19604_/Y VGND VGND VPWR VPWR _19614_/X sky130_fd_sc_hd__and2_4
XANTENNA__17533__A _13262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16826_ _16533_/X _16824_/X _16825_/Y VGND VGND VPWR VPWR _16826_/X sky130_fd_sc_hd__o21a_4
XFILLER_54_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16757_ _11772_/X VGND VGND VPWR VPWR _16757_/X sky130_fd_sc_hd__buf_2
X_19545_ _19545_/A _19545_/B VGND VGND VPWR VPWR _19831_/A sky130_fd_sc_hd__or2_4
XFILLER_94_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13969_ _12468_/A _13969_/B _13969_/C VGND VGND VPWR VPWR _13973_/B sky130_fd_sc_hd__and3_4
XANTENNA__12677__A _12979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15708_ _12240_/A _23108_/Q VGND VGND VPWR VPWR _15708_/X sky130_fd_sc_hd__or2_4
XFILLER_0_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15053__A _14773_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21896__A2 _21895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19476_ _19806_/A _19475_/Y VGND VGND VPWR VPWR _19476_/X sky130_fd_sc_hd__or2_4
XANTENNA__24400__CLK _23281_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16688_ _16688_/A VGND VGND VPWR VPWR _16689_/B sky130_fd_sc_hd__inv_2
XANTENNA__20894__A _20772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18427_ _18330_/X _18404_/X _18373_/X _18426_/X VGND VGND VPWR VPWR _18427_/X sky130_fd_sc_hd__o22a_4
X_15639_ _13886_/A _15639_/B _15638_/X VGND VGND VPWR VPWR _15639_/X sky130_fd_sc_hd__and3_4
XANTENNA__14892__A _14114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18358_ _17903_/A _22990_/B VGND VGND VPWR VPWR _18358_/X sky130_fd_sc_hd__or2_4
XFILLER_148_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17309_ _17308_/X VGND VGND VPWR VPWR _17310_/B sky130_fd_sc_hd__inv_2
XFILLER_30_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18289_ _17975_/X _18285_/Y _18089_/X _18288_/Y VGND VGND VPWR VPWR _18289_/X sky130_fd_sc_hd__a211o_4
XFILLER_174_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13301__A _13301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20320_ _20320_/A _20450_/B VGND VGND VPWR VPWR _20320_/X sky130_fd_sc_hd__or2_4
XFILLER_147_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20251_ _20251_/A VGND VGND VPWR VPWR _20251_/X sky130_fd_sc_hd__buf_2
XFILLER_127_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22073__A2 _22067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16612__A _16646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21820__A2 _21815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20182_ _20182_/A _20181_/Y VGND VGND VPWR VPWR _20182_/X sky130_fd_sc_hd__or2_4
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11756__A _11755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15228__A _14771_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23941_ _23557_/CLK _23941_/D VGND VGND VPWR VPWR _13512_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_130_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23872_ _23649_/CLK _23872_/D VGND VGND VPWR VPWR _23872_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22823_ _22819_/X _15117_/Y VGND VGND VPWR VPWR _22823_/X sky130_fd_sc_hd__or2_4
XFILLER_84_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12587__A _12587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21336__B2 _21331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22754_ SYSTICKCLKDIV[3] _22781_/A SYSTICKCLKDIV[2] _22753_/Y VGND VGND VPWR VPWR
+ _22754_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15015__A1 _14012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21705_ _21705_/A VGND VGND VPWR VPWR _21705_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22685_ _22484_/X _22658_/A _23125_/Q _22648_/A VGND VGND VPWR VPWR _22685_/X sky130_fd_sc_hd__o22a_4
X_24424_ _23347_/CLK _18860_/X HRESETn VGND VGND VPWR VPWR _24424_/Q sky130_fd_sc_hd__dfrtp_4
X_21636_ _21568_/X _21634_/X _15854_/B _21631_/X VGND VGND VPWR VPWR _23747_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21639__A2 _21634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24355_ _24388_/CLK _24355_/D HRESETn VGND VGND VPWR VPWR _19053_/A sky130_fd_sc_hd__dfstp_4
XFILLER_60_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21567_ _21565_/X _21566_/X _23780_/Q _21561_/X VGND VGND VPWR VPWR _23780_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14307__A _14307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13211__A _11682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23306_ _23404_/CLK _23306_/D VGND VGND VPWR VPWR _12785_/B sky130_fd_sc_hd__dfxtp_4
X_20518_ _20470_/X _20517_/X _24394_/Q _20429_/X VGND VGND VPWR VPWR _20518_/X sky130_fd_sc_hd__o22a_4
X_21498_ _21278_/X _21492_/X _13477_/B _21496_/X VGND VGND VPWR VPWR _23813_/D sky130_fd_sc_hd__o22a_4
XFILLER_158_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24286_ _24287_/CLK _19302_/X HRESETn VGND VGND VPWR VPWR _19235_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_158_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14026__B _23776_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23237_ _23397_/CLK _22514_/X VGND VGND VPWR VPWR _23237_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20449_ _11575_/A VGND VGND VPWR VPWR _20450_/A sky130_fd_sc_hd__inv_2
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16522__A _16521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23168_ _23203_/CLK _23168_/D VGND VGND VPWR VPWR _23168_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11666__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22119_ _22117_/X _22111_/X _23467_/Q _22118_/X VGND VGND VPWR VPWR _22119_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15138__A _14277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15990_ _15961_/A _15990_/B _15990_/C VGND VGND VPWR VPWR _15994_/B sky130_fd_sc_hd__and3_4
X_23099_ _23515_/CLK _23099_/D VGND VGND VPWR VPWR _14531_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14941_ _14783_/X _14935_/X _14940_/X VGND VGND VPWR VPWR _14941_/X sky130_fd_sc_hd__or3_4
XFILLER_75_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14977__A _15076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17660_ _17660_/A _17660_/B VGND VGND VPWR VPWR _17661_/A sky130_fd_sc_hd__or2_4
XANTENNA__17353__A _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23074__B _23079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14872_ _11895_/X _14934_/B VGND VGND VPWR VPWR _14872_/X sky130_fd_sc_hd__or2_4
XFILLER_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16451__B1 _11608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16611_ _16611_/A _23538_/Q VGND VGND VPWR VPWR _16611_/X sky130_fd_sc_hd__or2_4
X_13823_ _13823_/A _13897_/B VGND VGND VPWR VPWR _13823_/X sky130_fd_sc_hd__or2_4
X_17591_ _17546_/Y _17583_/X _17590_/X VGND VGND VPWR VPWR _17591_/X sky130_fd_sc_hd__o21a_4
X_19330_ _19330_/A VGND VGND VPWR VPWR _19330_/Y sky130_fd_sc_hd__inv_2
X_16542_ _12108_/A _16542_/B _16542_/C VGND VGND VPWR VPWR _16542_/X sky130_fd_sc_hd__or3_4
X_13754_ _12927_/A _24062_/Q VGND VGND VPWR VPWR _13755_/C sky130_fd_sc_hd__or2_4
XFILLER_62_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21878__A2 _21875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12705_ _12735_/A _12803_/B VGND VGND VPWR VPWR _12707_/B sky130_fd_sc_hd__or2_4
X_19261_ _19256_/B VGND VGND VPWR VPWR _19261_/Y sky130_fd_sc_hd__inv_2
X_16473_ _16491_/A _16413_/B VGND VGND VPWR VPWR _16473_/X sky130_fd_sc_hd__or2_4
XANTENNA__19940__B2 _20512_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13685_ _15446_/A _13768_/B VGND VGND VPWR VPWR _13687_/B sky130_fd_sc_hd__or2_4
X_18212_ _17770_/Y _18182_/X _17770_/Y _18182_/X VGND VGND VPWR VPWR _18212_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15424_ _13657_/A _15424_/B _15424_/C VGND VGND VPWR VPWR _15428_/B sky130_fd_sc_hd__and3_4
X_12636_ _12973_/A _23339_/Q VGND VGND VPWR VPWR _12638_/B sky130_fd_sc_hd__or2_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22827__A1 _17425_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19192_ _24325_/Q _19145_/X _19191_/Y VGND VGND VPWR VPWR _24325_/D sky130_fd_sc_hd__o21a_4
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ _18020_/X _18141_/X _18065_/X _18142_/X VGND VGND VPWR VPWR _18143_/X sky130_fd_sc_hd__o22a_4
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _15318_/A _23128_/Q VGND VGND VPWR VPWR _15357_/B sky130_fd_sc_hd__or2_4
XFILLER_54_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12567_ _11915_/A VGND VGND VPWR VPWR _12570_/A sky130_fd_sc_hd__buf_2
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14217__A _14201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13121__A _13099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14306_ _12445_/A _14304_/X _14306_/C VGND VGND VPWR VPWR _14310_/B sky130_fd_sc_hd__and3_4
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11518_ _11518_/A _11518_/B VGND VGND VPWR VPWR _11519_/B sky130_fd_sc_hd__or2_4
X_18074_ _18150_/A _17572_/X VGND VGND VPWR VPWR _18074_/X sky130_fd_sc_hd__or2_4
X_15286_ _15267_/A _15351_/B VGND VGND VPWR VPWR _15286_/X sky130_fd_sc_hd__or2_4
X_12498_ _12498_/A VGND VGND VPWR VPWR _12499_/A sky130_fd_sc_hd__buf_2
XFILLER_89_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17025_ _17025_/A VGND VGND VPWR VPWR _17025_/Y sky130_fd_sc_hd__inv_2
X_14237_ _14616_/A _14237_/B _14237_/C VGND VGND VPWR VPWR _14242_/B sky130_fd_sc_hd__and3_4
XANTENNA__22055__A2 _22053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14168_ _15007_/A VGND VGND VPWR VPWR _14169_/A sky130_fd_sc_hd__buf_2
XANTENNA__17247__B _17246_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13119_ _12758_/A _13035_/B VGND VGND VPWR VPWR _13119_/X sky130_fd_sc_hd__or2_4
XFILLER_140_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18976_ _24400_/Q VGND VGND VPWR VPWR _18976_/Y sky130_fd_sc_hd__inv_2
X_14099_ _14103_/A _14099_/B _14098_/X VGND VGND VPWR VPWR _14099_/X sky130_fd_sc_hd__and3_4
XFILLER_98_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17927_ _17825_/X _17167_/X _17230_/X _17175_/X VGND VGND VPWR VPWR _17927_/X sky130_fd_sc_hd__o22a_4
XFILLER_152_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13791__A _13791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17234__A2 _17187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17858_ _17837_/X _17208_/X _17838_/X _17211_/X VGND VGND VPWR VPWR _17858_/X sky130_fd_sc_hd__o22a_4
XFILLER_61_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16809_ _16606_/A _16805_/X _16808_/X VGND VGND VPWR VPWR _16809_/X sky130_fd_sc_hd__or3_4
XFILLER_81_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17789_ _17010_/B _17788_/Y _17011_/Y VGND VGND VPWR VPWR _17789_/X sky130_fd_sc_hd__o21a_4
XFILLER_19_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19528_ _19528_/A _19528_/B VGND VGND VPWR VPWR _19740_/A sky130_fd_sc_hd__or2_4
XANTENNA__12200__A _12569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_52_0_HCLK clkbuf_7_53_0_HCLK/A VGND VGND VPWR VPWR _23204_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_62_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21513__A _21506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19459_ HRDATA[1] VGND VGND VPWR VPWR _19459_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18094__A _18538_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16607__A _11705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22470_ _22468_/X _22462_/X _14337_/B _22469_/X VGND VGND VPWR VPWR _23260_/D sky130_fd_sc_hd__o22a_4
XFILLER_33_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21421_ _21420_/X VGND VGND VPWR VPWR _21455_/A sky130_fd_sc_hd__buf_2
XANTENNA__19918__A _19438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13031__A _12911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24140_ _24137_/CLK _20087_/Y HRESETn VGND VGND VPWR VPWR _24140_/Q sky130_fd_sc_hd__dfrtp_4
X_21352_ _21338_/A VGND VGND VPWR VPWR _21352_/X sky130_fd_sc_hd__buf_2
XANTENNA__19637__B HRDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20303_ _20226_/X VGND VGND VPWR VPWR _20977_/A sky130_fd_sc_hd__buf_2
XFILLER_163_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24071_ _24039_/CLK _24071_/D VGND VGND VPWR VPWR _24071_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21283_ _21283_/A VGND VGND VPWR VPWR _21283_/X sky130_fd_sc_hd__buf_2
XANTENNA__17438__A _13947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12870__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20234_ _16915_/C _18779_/X _20233_/Y VGND VGND VPWR VPWR _20234_/X sky130_fd_sc_hd__o21a_4
X_23022_ _23008_/X _23020_/X _23022_/C VGND VGND VPWR VPWR _23022_/X sky130_fd_sc_hd__and3_4
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20165_ _24446_/Q VGND VGND VPWR VPWR _20165_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23320__CLK _23416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24446__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20096_ _11635_/A _20095_/X VGND VGND VPWR VPWR _20194_/A sky130_fd_sc_hd__nor2_4
XFILLER_76_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21557__B2 _21549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22754__B1 SYSTICKCLKDIV[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17173__A _17172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23924_ _23668_/CLK _21325_/X VGND VGND VPWR VPWR _21317_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23855_ _23983_/CLK _21433_/X VGND VGND VPWR VPWR _16287_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22506__B1 _12671_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22806_ _15117_/Y _22804_/X VGND VGND VPWR VPWR HWDATA[1] sky130_fd_sc_hd__nor2_4
XFILLER_72_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23786_ _23467_/CLK _21552_/X VGND VGND VPWR VPWR _23786_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22519__A _22505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20998_ _20997_/X VGND VGND VPWR VPWR _20998_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21423__A _21438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22737_ _22737_/A _18576_/B _20598_/B VGND VGND VPWR VPWR _22737_/X sky130_fd_sc_hd__and3_4
XFILLER_53_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16517__A _16163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13470_ _13443_/A _13470_/B VGND VGND VPWR VPWR _13471_/C sky130_fd_sc_hd__or2_4
XFILLER_125_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22668_ _22454_/X _22665_/X _15493_/B _22662_/X VGND VGND VPWR VPWR _23138_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12421_ _12320_/Y _12418_/X VGND VGND VPWR VPWR _12422_/A sky130_fd_sc_hd__or2_4
XFILLER_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24407_ _24419_/CLK _24407_/D HRESETn VGND VGND VPWR VPWR _24407_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21619_ _21539_/X _21613_/X _16253_/B _21617_/X VGND VGND VPWR VPWR _23759_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22285__A2 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22599_ _22420_/X _22594_/X _16415_/B _22598_/X VGND VGND VPWR VPWR _22599_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14037__A _13719_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15140_ _15294_/A _15211_/B VGND VGND VPWR VPWR _15141_/C sky130_fd_sc_hd__or2_4
X_12352_ _11755_/X _12352_/B _12351_/X VGND VGND VPWR VPWR _12352_/X sky130_fd_sc_hd__or3_4
X_24338_ _24277_/CLK _24338_/D HRESETn VGND VGND VPWR VPWR _19159_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13876__A _14386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15071_ _15095_/A _23157_/Q VGND VGND VPWR VPWR _15073_/B sky130_fd_sc_hd__or2_4
XANTENNA__22037__A2 _22010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12283_ _13139_/A _12393_/B VGND VGND VPWR VPWR _12283_/X sky130_fd_sc_hd__or2_4
XANTENNA__12780__A _13067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24269_ _24495_/CLK _24269_/D HRESETn VGND VGND VPWR VPWR _24269_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23069__B _23079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16252__A _16099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14022_ _13705_/A _23744_/Q VGND VGND VPWR VPWR _14022_/X sky130_fd_sc_hd__or2_4
XFILLER_88_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21796__A1 _21584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21796__B2 _21795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18830_ _15251_/A _18824_/X _24439_/Q _18825_/X VGND VGND VPWR VPWR _24439_/D sky130_fd_sc_hd__o22a_4
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23085__A _20216_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15973_ _11903_/X _16039_/B VGND VGND VPWR VPWR _15973_/X sky130_fd_sc_hd__or2_4
X_18761_ _18220_/A _18176_/A _17626_/Y _18758_/X VGND VGND VPWR VPWR _18773_/B sky130_fd_sc_hd__a211o_4
X_17712_ _17712_/A _17710_/A VGND VGND VPWR VPWR _17767_/A sky130_fd_sc_hd__or2_4
X_14924_ _14916_/X _14922_/X _14923_/X VGND VGND VPWR VPWR _14924_/X sky130_fd_sc_hd__and3_4
XANTENNA__17083__A _17188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18692_ _18518_/X _17324_/X _18335_/A VGND VGND VPWR VPWR _18692_/X sky130_fd_sc_hd__a21o_4
XFILLER_152_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17643_ _17642_/X VGND VGND VPWR VPWR _17643_/Y sky130_fd_sc_hd__inv_2
X_14855_ _13662_/A _14851_/X _14854_/X VGND VGND VPWR VPWR _14855_/X sky130_fd_sc_hd__or3_4
XFILLER_64_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13806_ _15398_/A _13801_/X _13805_/X VGND VGND VPWR VPWR _13806_/X sky130_fd_sc_hd__or3_4
X_17574_ _16162_/X VGND VGND VPWR VPWR _17574_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23963__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14786_ _14786_/A VGND VGND VPWR VPWR _15081_/A sky130_fd_sc_hd__buf_2
XANTENNA__18177__B1 _18176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11998_ _11963_/A _11996_/X _11997_/X VGND VGND VPWR VPWR _11999_/C sky130_fd_sc_hd__and3_4
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19313_ _19313_/A VGND VGND VPWR VPWR _19313_/Y sky130_fd_sc_hd__inv_2
X_16525_ _16525_/A VGND VGND VPWR VPWR _16525_/Y sky130_fd_sc_hd__inv_2
X_13737_ _12600_/A VGND VGND VPWR VPWR _15502_/A sky130_fd_sc_hd__buf_2
Xclkbuf_6_39_0_HCLK clkbuf_6_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_79_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12955__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15331__A _15377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16456_ _13377_/A VGND VGND VPWR VPWR _16474_/A sky130_fd_sc_hd__buf_2
X_19244_ _24295_/Q _19244_/B VGND VGND VPWR VPWR _19245_/B sky130_fd_sc_hd__and2_4
X_13668_ _13632_/A _13758_/B VGND VGND VPWR VPWR _13669_/C sky130_fd_sc_hd__or2_4
X_15407_ _13632_/A _15478_/B VGND VGND VPWR VPWR _15408_/C sky130_fd_sc_hd__or2_4
XANTENNA__24319__CLK _24287_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12619_ _12632_/A _12619_/B VGND VGND VPWR VPWR _12619_/X sky130_fd_sc_hd__or2_4
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19175_ _19155_/B VGND VGND VPWR VPWR _19175_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15050__B _23253_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16387_ _15956_/A _16387_/B VGND VGND VPWR VPWR _16389_/B sky130_fd_sc_hd__or2_4
XFILLER_129_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13599_ _13957_/A VGND VGND VPWR VPWR _14296_/A sky130_fd_sc_hd__buf_2
XFILLER_129_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18126_ _18126_/A _17932_/Y VGND VGND VPWR VPWR _18126_/X sky130_fd_sc_hd__or2_4
X_15338_ _11752_/A _15338_/B _15337_/X VGND VGND VPWR VPWR _15338_/X sky130_fd_sc_hd__or3_4
XANTENNA__13786__A _11928_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18057_ _18538_/A VGND VGND VPWR VPWR _18389_/A sky130_fd_sc_hd__buf_2
XANTENNA__12690__A _12690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15269_ _15269_/A _15267_/X _15268_/X VGND VGND VPWR VPWR _15269_/X sky130_fd_sc_hd__and3_4
XFILLER_145_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24469__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17008_ _17008_/A VGND VGND VPWR VPWR _17008_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21787__B2 _21781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19473__A HRDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18959_ _18959_/A VGND VGND VPWR VPWR _18959_/X sky130_fd_sc_hd__buf_2
XFILLER_6_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22200__A2 _22194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21970_ _21855_/X _21967_/X _15481_/B _21964_/X VGND VGND VPWR VPWR _23554_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14410__A _12576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20921_ _20863_/A _20919_/X _20920_/X VGND VGND VPWR VPWR _20921_/X sky130_fd_sc_hd__a21o_4
XFILLER_54_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13026__A _12506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23640_ _23770_/CLK _23640_/D VGND VGND VPWR VPWR _23640_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20852_ _20754_/X _20851_/X _19137_/A _20761_/X VGND VGND VPWR VPWR _20852_/X sky130_fd_sc_hd__o22a_4
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19904__A1 _19576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21243__A _21528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23571_ _23764_/CLK _21947_/X VGND VGND VPWR VPWR _23571_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12865__A _12889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20783_ _24415_/Q _20617_/B VGND VGND VPWR VPWR _20783_/Y sky130_fd_sc_hd__nand2_4
XFILLER_168_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16337__A _13414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21711__B2 _21710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22522_ _22489_/A VGND VGND VPWR VPWR _22522_/X sky130_fd_sc_hd__buf_2
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12584__B _12584_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22453_ _22452_/X _22450_/X _15789_/B _22445_/X VGND VGND VPWR VPWR _23267_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22267__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21404_ _21290_/X _21398_/X _23872_/Q _21402_/X VGND VGND VPWR VPWR _23872_/D sky130_fd_sc_hd__o22a_4
X_22384_ _22134_/X _22383_/X _15668_/B _22380_/X VGND VGND VPWR VPWR _23300_/D sky130_fd_sc_hd__o22a_4
XFILLER_157_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22074__A _22041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24123_ _23416_/CLK _24123_/D HRESETn VGND VGND VPWR VPWR _22766_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13696__A _13696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21335_ _21256_/X _21334_/X _16054_/B _21331_/X VGND VGND VPWR VPWR _23918_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22019__A2 _22017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16072__A _16048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24054_ _23544_/CLK _21078_/X VGND VGND VPWR VPWR _14884_/B sky130_fd_sc_hd__dfxtp_4
X_21266_ _20531_/A VGND VGND VPWR VPWR _21266_/X sky130_fd_sc_hd__buf_2
XFILLER_2_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22802__A _22799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21778__B2 _21774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23005_ _22977_/X _16986_/A _22989_/X _23004_/X VGND VGND VPWR VPWR _23006_/A sky130_fd_sc_hd__a211o_4
XFILLER_2_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20217_ _16937_/X _17033_/A _17017_/B _20217_/D VGND VGND VPWR VPWR _20217_/X sky130_fd_sc_hd__and4_4
XANTENNA__18643__A1 _17793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21197_ _20416_/X _21191_/X _16280_/B _21195_/X VGND VGND VPWR VPWR _23983_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12105__A _12105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20148_ _20196_/A _20147_/X VGND VGND VPWR VPWR _20148_/X sky130_fd_sc_hd__or2_4
X_12970_ _12970_/A _23497_/Q VGND VGND VPWR VPWR _12972_/B sky130_fd_sc_hd__or2_4
X_20079_ _19960_/X VGND VGND VPWR VPWR _20079_/X sky130_fd_sc_hd__buf_2
XANTENNA__20738__C1 _20737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23907_ _23939_/CLK _21350_/X VGND VGND VPWR VPWR _15819_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_79_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11921_ _11891_/X VGND VGND VPWR VPWR _11975_/A sky130_fd_sc_hd__buf_2
XFILLER_46_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14640_ _14685_/A _14640_/B _14639_/X VGND VGND VPWR VPWR _14641_/C sky130_fd_sc_hd__and3_4
X_11852_ _11603_/A VGND VGND VPWR VPWR _11853_/A sky130_fd_sc_hd__inv_2
X_23838_ _23582_/CLK _21457_/X VGND VGND VPWR VPWR _13758_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14974__B _14895_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _15423_/A _23546_/Q VGND VGND VPWR VPWR _14571_/X sky130_fd_sc_hd__or2_4
XPHY_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _13092_/A VGND VGND VPWR VPWR _13400_/A sky130_fd_sc_hd__buf_2
X_23769_ _23770_/CLK _23769_/D VGND VGND VPWR VPWR _14788_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20505__A2 _20443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16310_ _13367_/A VGND VGND VPWR VPWR _16313_/A sky130_fd_sc_hd__buf_2
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21702__B2 _21667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13522_ _13534_/A _23685_/Q VGND VGND VPWR VPWR _13524_/B sky130_fd_sc_hd__or2_4
XANTENNA__15151__A _13954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17290_ _14700_/X VGND VGND VPWR VPWR _17290_/X sky130_fd_sc_hd__buf_2
XPHY_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17382__A1 _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17382__B2 _17381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16241_ _16240_/X VGND VGND VPWR VPWR _16243_/B sky130_fd_sc_hd__inv_2
X_13453_ _13453_/A _13452_/X VGND VGND VPWR VPWR _13453_/X sky130_fd_sc_hd__and2_4
XFILLER_16_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14990__A _14171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12404_ _15851_/A _12314_/B VGND VGND VPWR VPWR _12405_/C sky130_fd_sc_hd__or2_4
XANTENNA__21466__B1 _15227_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16172_ _13397_/A VGND VGND VPWR VPWR _16216_/A sky130_fd_sc_hd__buf_2
XFILLER_142_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13384_ _13384_/A _13309_/B VGND VGND VPWR VPWR _13384_/X sky130_fd_sc_hd__or2_4
XFILLER_126_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17134__A1 _15252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15123_ _11898_/A _15123_/B VGND VGND VPWR VPWR _15123_/X sky130_fd_sc_hd__or2_4
XANTENNA__17078__A _11643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12335_ _15324_/A VGND VGND VPWR VPWR _12336_/A sky130_fd_sc_hd__buf_2
XFILLER_127_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18882__A1 _15380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19931_ _19920_/X VGND VGND VPWR VPWR _19931_/X sky130_fd_sc_hd__buf_2
X_15054_ _15075_/A _23349_/Q VGND VGND VPWR VPWR _15054_/X sky130_fd_sc_hd__or2_4
XFILLER_99_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12266_ _12266_/A VGND VGND VPWR VPWR _12726_/A sky130_fd_sc_hd__buf_2
XFILLER_135_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22712__A _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14214__B _23679_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21769__B2 _21767_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14005_ _12474_/A _23104_/Q VGND VGND VPWR VPWR _14007_/B sky130_fd_sc_hd__or2_4
XANTENNA__18634__A1 _17109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19862_ _19842_/A _19861_/X _19788_/A VGND VGND VPWR VPWR _19862_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__17806__A _17805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12015__A _12015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12197_ _15444_/A VGND VGND VPWR VPWR _12198_/A sky130_fd_sc_hd__buf_2
XFILLER_68_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18813_ _15784_/X _18810_/X _20159_/A _18811_/X VGND VGND VPWR VPWR _24452_/D sky130_fd_sc_hd__o22a_4
X_19793_ _19696_/X _19791_/Y _22737_/A _19573_/A VGND VGND VPWR VPWR _19793_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22718__B1 _15501_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11854__A _11854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18744_ _18744_/A _17108_/X VGND VGND VPWR VPWR _18744_/X sky130_fd_sc_hd__or2_4
X_15956_ _15956_/A VGND VGND VPWR VPWR _15957_/A sky130_fd_sc_hd__buf_2
XFILLER_37_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12669__B _12669_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14907_ _13955_/A _14907_/B _14907_/C VGND VGND VPWR VPWR _14907_/X sky130_fd_sc_hd__and3_4
XANTENNA__11573__B IRQ[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15887_ _15887_/A _15883_/X _15887_/C VGND VGND VPWR VPWR _15887_/X sky130_fd_sc_hd__or3_4
X_18675_ _17316_/X _18675_/B VGND VGND VPWR VPWR _18675_/X sky130_fd_sc_hd__or2_4
XFILLER_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17541__A _12678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17626_ _17626_/A VGND VGND VPWR VPWR _17626_/Y sky130_fd_sc_hd__inv_2
X_14838_ _14658_/A _14754_/B VGND VGND VPWR VPWR _14839_/C sky130_fd_sc_hd__or2_4
XANTENNA__14884__B _14884_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22159__A _22147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24141__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17557_ _11611_/B _17035_/A VGND VGND VPWR VPWR _17557_/X sky130_fd_sc_hd__and2_4
X_14769_ _14769_/A VGND VGND VPWR VPWR _15106_/A sky130_fd_sc_hd__buf_2
XANTENNA__22497__A2 _22494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12685__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15061__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16508_ _16164_/X _16445_/B VGND VGND VPWR VPWR _16510_/B sky130_fd_sc_hd__or2_4
XFILLER_108_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12985__A2 _12982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17488_ _17486_/Y _17487_/X VGND VGND VPWR VPWR _17600_/D sky130_fd_sc_hd__or2_4
XFILLER_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15996__A _15969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19227_ _24278_/Q _19321_/A VGND VGND VPWR VPWR _19227_/X sky130_fd_sc_hd__and2_4
XANTENNA__22249__A2 _22244_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16439_ _16101_/A _16439_/B VGND VGND VPWR VPWR _16440_/C sky130_fd_sc_hd__or2_4
XFILLER_34_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24291__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19158_ _19158_/A _19158_/B VGND VGND VPWR VPWR _19159_/B sky130_fd_sc_hd__and2_4
XFILLER_121_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18109_ _17903_/A VGND VGND VPWR VPWR _18111_/A sky130_fd_sc_hd__buf_2
XFILLER_145_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18873__A1 _14261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19089_ _19087_/Y _19088_/Y _11524_/B VGND VGND VPWR VPWR _19089_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14405__A _14512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21120_ _20819_/X _21118_/X _24030_/Q _21115_/X VGND VGND VPWR VPWR _24030_/D sky130_fd_sc_hd__o22a_4
XFILLER_132_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22622__A _22622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21051_ _20531_/X _21045_/X _24074_/Q _21049_/X VGND VGND VPWR VPWR _21051_/X sky130_fd_sc_hd__o22a_4
XFILLER_154_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20002_ _20001_/X VGND VGND VPWR VPWR _20002_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13963__B _24032_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21238__A _21238_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19931__A _19920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15236__A _14201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12579__B _12579_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22185__B2 _22184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21953_ _21960_/A VGND VGND VPWR VPWR _21953_/X sky130_fd_sc_hd__buf_2
XFILLER_54_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21932__B2 _21927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20904_ _20703_/X _20903_/X _24378_/Q _18893_/A VGND VGND VPWR VPWR _20904_/X sky130_fd_sc_hd__o22a_4
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21884_ _21883_/X _21875_/X _23606_/Q _21809_/X VGND VGND VPWR VPWR _23606_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24366__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _24039_/CLK _21844_/X VGND VGND VPWR VPWR _23623_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ _20834_/X VGND VGND VPWR VPWR _20835_/Y sky130_fd_sc_hd__inv_2
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12595__A _12659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_22_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_23554_ _23587_/CLK _23554_/D VGND VGND VPWR VPWR _15481_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20766_ _20695_/X _20752_/Y _20764_/X _20765_/Y _20714_/X VGND VGND VPWR VPWR _20767_/B
+ sky130_fd_sc_hd__a32o_4
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21160__A2 _21155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22505_ _22505_/A VGND VGND VPWR VPWR _22505_/X sky130_fd_sc_hd__buf_2
XFILLER_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23485_ _23678_/CLK _22077_/X VGND VGND VPWR VPWR _13845_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20697_ _20697_/A VGND VGND VPWR VPWR _20697_/X sky130_fd_sc_hd__buf_2
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22436_ _22435_/X _22426_/X _12759_/B _22433_/X VGND VGND VPWR VPWR _23274_/D sky130_fd_sc_hd__o22a_4
XFILLER_109_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21999__B2 _21993_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11939__A _16138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22660__A2 _22658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22367_ _22105_/X _22362_/X _16398_/B _22366_/X VGND VGND VPWR VPWR _22367_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14315__A _13656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24106_ _23558_/CLK _24106_/D VGND VGND VPWR VPWR _24106_/Q sky130_fd_sc_hd__dfxtp_4
X_12120_ _16080_/A VGND VGND VPWR VPWR _12164_/A sky130_fd_sc_hd__buf_2
X_21318_ _21028_/A VGND VGND VPWR VPWR _21420_/B sky130_fd_sc_hd__buf_2
X_22298_ _22291_/A VGND VGND VPWR VPWR _22298_/X sky130_fd_sc_hd__buf_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24037_ _23493_/CLK _21110_/X VGND VGND VPWR VPWR _24037_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12051_ _12051_/A _24051_/Q VGND VGND VPWR VPWR _12053_/B sky130_fd_sc_hd__or2_4
X_21249_ _21534_/A VGND VGND VPWR VPWR _21249_/X sky130_fd_sc_hd__buf_2
XFILLER_132_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21148__A _21155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11674__A _11674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15810_ _12852_/A _15865_/B VGND VGND VPWR VPWR _15810_/X sky130_fd_sc_hd__or2_4
XANTENNA__15146__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16790_ _16647_/A _16790_/B _16790_/C VGND VGND VPWR VPWR _16794_/B sky130_fd_sc_hd__and3_4
XFILLER_19_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14050__A _11674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19577__C1 _19576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15741_ _13067_/A VGND VGND VPWR VPWR _15741_/X sky130_fd_sc_hd__buf_2
X_12953_ _12953_/A _12953_/B _12952_/X VGND VGND VPWR VPWR _12954_/C sky130_fd_sc_hd__and3_4
XANTENNA__24164__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14985__A _14169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_104_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR _24039_/CLK sky130_fd_sc_hd__clkbuf_1
X_11904_ _11903_/X VGND VGND VPWR VPWR _11904_/X sky130_fd_sc_hd__buf_2
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15672_ _13139_/A _15744_/B VGND VGND VPWR VPWR _15672_/X sky130_fd_sc_hd__or2_4
XFILLER_2_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18460_ _17798_/A _17374_/A VGND VGND VPWR VPWR _18460_/X sky130_fd_sc_hd__and2_4
X_12884_ _12884_/A _23913_/Q VGND VGND VPWR VPWR _12884_/X sky130_fd_sc_hd__or2_4
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17411_ _17153_/A _17439_/B VGND VGND VPWR VPWR _17412_/B sky130_fd_sc_hd__or2_4
X_14623_ _14623_/A VGND VGND VPWR VPWR _14834_/A sky130_fd_sc_hd__buf_2
X_11835_ _11792_/X _21655_/A VGND VGND VPWR VPWR _11837_/B sky130_fd_sc_hd__or2_4
X_18391_ _17594_/X _17638_/Y _18320_/A _17452_/X VGND VGND VPWR VPWR _18391_/X sky130_fd_sc_hd__o22a_4
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17297_/B VGND VGND VPWR VPWR _17342_/Y sky130_fd_sc_hd__inv_2
XPHY_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14270_/A _23514_/Q VGND VGND VPWR VPWR _14554_/X sky130_fd_sc_hd__or2_4
XPHY_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11704_/X VGND VGND VPWR VPWR _11834_/A sky130_fd_sc_hd__buf_2
XANTENNA__21151__A2 _21148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14209__B _23167_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13505_ _13534_/A _24037_/Q VGND VGND VPWR VPWR _13505_/X sky130_fd_sc_hd__or2_4
XFILLER_147_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17273_ _14334_/X VGND VGND VPWR VPWR _17273_/Y sky130_fd_sc_hd__inv_2
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _12362_/A _14485_/B VGND VGND VPWR VPWR _14485_/X sky130_fd_sc_hd__or2_4
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18192__A _18310_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11697_ _11697_/A VGND VGND VPWR VPWR _11698_/A sky130_fd_sc_hd__buf_2
XANTENNA__24314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16224_ _16231_/A _16224_/B VGND VGND VPWR VPWR _16224_/X sky130_fd_sc_hd__or2_4
XANTENNA__21439__B1 _12549_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19012_ _11536_/A _11535_/X _19005_/Y VGND VGND VPWR VPWR _19012_/Y sky130_fd_sc_hd__a21oi_4
X_13436_ _13462_/A _23685_/Q VGND VGND VPWR VPWR _13438_/B sky130_fd_sc_hd__or2_4
XANTENNA__20227__A _20226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22100__B2 _22094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16155_ _16155_/A _16153_/X _16155_/C VGND VGND VPWR VPWR _16159_/B sky130_fd_sc_hd__and3_4
XANTENNA__11849__A _11686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13367_ _13367_/A VGND VGND VPWR VPWR _13413_/A sky130_fd_sc_hd__buf_2
XANTENNA__18855__A1 _12678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14225__A _14225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15106_ _15106_/A _15102_/X _15106_/C VGND VGND VPWR VPWR _15114_/B sky130_fd_sc_hd__or3_4
X_12318_ _12882_/A _12275_/X _12285_/X _12308_/X _12317_/X VGND VGND VPWR VPWR _12318_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_114_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16086_ _16016_/Y _16085_/X VGND VGND VPWR VPWR _16086_/X sky130_fd_sc_hd__and2_4
X_13298_ _13321_/A _13296_/X _13297_/X VGND VGND VPWR VPWR _13299_/C sky130_fd_sc_hd__and3_4
XFILLER_154_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22442__A _20595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19914_ _20867_/A VGND VGND VPWR VPWR _21007_/A sky130_fd_sc_hd__buf_2
X_15037_ _13974_/A _23093_/Q VGND VGND VPWR VPWR _15039_/B sky130_fd_sc_hd__or2_4
X_12249_ _14450_/A VGND VGND VPWR VPWR _13016_/A sky130_fd_sc_hd__buf_2
XANTENNA__22403__A2 _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19845_ _17296_/A VGND VGND VPWR VPWR _21603_/A sky130_fd_sc_hd__buf_2
XANTENNA__13783__B _13781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19751__A _19539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19776_ _19705_/B _19787_/B VGND VGND VPWR VPWR _19776_/X sky130_fd_sc_hd__and2_4
X_16988_ _16988_/A _16988_/B VGND VGND VPWR VPWR _16989_/B sky130_fd_sc_hd__or2_4
XFILLER_37_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18727_ _18022_/X _17005_/X _18698_/B VGND VGND VPWR VPWR _18727_/X sky130_fd_sc_hd__o21a_4
XFILLER_37_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20112__D _20124_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15939_ _11903_/X VGND VGND VPWR VPWR _15982_/A sky130_fd_sc_hd__buf_2
XFILLER_114_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14895__A _14131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21914__B2 _21913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18658_ _18657_/X VGND VGND VPWR VPWR _18658_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21390__A2 _21384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18791__B1 _24468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17609_ _18415_/A _18415_/B _17387_/A _17609_/D VGND VGND VPWR VPWR _17636_/A sky130_fd_sc_hd__or4_4
X_18589_ _18589_/A VGND VGND VPWR VPWR _18589_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13304__A _13304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20620_ _20447_/X _20617_/Y _20619_/X _19043_/Y _20495_/X VGND VGND VPWR VPWR _20620_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21142__A2 _21141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21521__A _21134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20551_ _20501_/A _20550_/X VGND VGND VPWR VPWR _20551_/Y sky130_fd_sc_hd__nor2_4
X_23270_ _24039_/CLK _22446_/X VGND VGND VPWR VPWR _13273_/B sky130_fd_sc_hd__dfxtp_4
X_20482_ _20466_/X _20468_/Y _20479_/X _20480_/Y _20481_/X VGND VGND VPWR VPWR _20482_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_20_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22221_ _22169_/X _22194_/A _23413_/Q _22184_/A VGND VGND VPWR VPWR _23413_/D sky130_fd_sc_hd__o22a_4
XFILLER_146_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18846__A1 _17255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20653__A1 _18426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22152_ _22151_/X _22147_/X _13901_/B _22142_/X VGND VGND VPWR VPWR _23453_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21103_ _20531_/X _21097_/X _24042_/Q _21101_/X VGND VGND VPWR VPWR _24042_/D sky130_fd_sc_hd__o22a_4
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17446__A _17170_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22083_ _21877_/X _22081_/X _14834_/B _22078_/X VGND VGND VPWR VPWR _22083_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21034_ _21049_/A VGND VGND VPWR VPWR _21042_/A sky130_fd_sc_hd__buf_2
XFILLER_120_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24187__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20600__A _20847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22985_ _18448_/X _22973_/B VGND VGND VPWR VPWR _22986_/C sky130_fd_sc_hd__or2_4
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21905__B2 _21899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21936_ _21885_/X _21909_/A _23573_/Q _21899_/A VGND VGND VPWR VPWR _23573_/D sky130_fd_sc_hd__o22a_4
XFILLER_167_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15413__B _15470_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21867_ _20841_/A VGND VGND VPWR VPWR _21867_/X sky130_fd_sc_hd__buf_2
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23511_/CLK _23606_/D VGND VGND VPWR VPWR _23606_/Q sky130_fd_sc_hd__dfxtp_4
X_11620_ _13792_/A VGND VGND VPWR VPWR _12473_/A sky130_fd_sc_hd__buf_2
XFILLER_70_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20818_ _20818_/A VGND VGND VPWR VPWR _20819_/A sky130_fd_sc_hd__buf_2
XFILLER_11_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17337__A1 _15117_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21798_ _21791_/A VGND VGND VPWR VPWR _21798_/X sky130_fd_sc_hd__buf_2
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14029__B _24032_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21431__A _21431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23537_ _23537_/CLK _21999_/X VGND VGND VPWR VPWR _23537_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _24437_/Q IRQ[0] VGND VGND VPWR VPWR _11551_/X sky130_fd_sc_hd__and2_4
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20749_ HRDATA[11] _20843_/B VGND VGND VPWR VPWR _20751_/B sky130_fd_sc_hd__or2_4
XFILLER_11_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _14270_/A _14339_/B VGND VGND VPWR VPWR _14271_/C sky130_fd_sc_hd__or2_4
X_23468_ _23852_/CLK _22116_/X VGND VGND VPWR VPWR _12259_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13221_ _12362_/A VGND VGND VPWR VPWR _13253_/A sky130_fd_sc_hd__buf_2
XANTENNA__11669__A _12979_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22419_ _22418_/X _22414_/X _16751_/B _22409_/X VGND VGND VPWR VPWR _23281_/D sky130_fd_sc_hd__o22a_4
XFILLER_137_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22633__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23399_ _23303_/CLK _23399_/D VGND VGND VPWR VPWR _13240_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13152_ _13152_/A _23943_/Q VGND VGND VPWR VPWR _13152_/X sky130_fd_sc_hd__or2_4
XFILLER_124_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_29_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR _24397_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_151_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22262__A _22226_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12103_ _12103_/A _23827_/Q VGND VGND VPWR VPWR _12103_/X sky130_fd_sc_hd__or2_4
XANTENNA__13884__A _13884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13083_ _13100_/A _13083_/B _13082_/X VGND VGND VPWR VPWR _13092_/B sky130_fd_sc_hd__or3_4
X_17960_ _17779_/X _17959_/X _17779_/X _17959_/X VGND VGND VPWR VPWR _17960_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12034_ _16594_/A VGND VGND VPWR VPWR _16691_/A sky130_fd_sc_hd__buf_2
X_16911_ _12025_/A _16904_/Y _16911_/C _16911_/D VGND VGND VPWR VPWR _16911_/X sky130_fd_sc_hd__or4_4
XFILLER_104_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17891_ _17260_/A _17887_/X _17890_/X VGND VGND VPWR VPWR _17891_/X sky130_fd_sc_hd__o21a_4
XFILLER_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19630_ _19537_/B _19622_/B VGND VGND VPWR VPWR _19630_/X sky130_fd_sc_hd__and2_4
X_16842_ _15391_/X _16842_/B VGND VGND VPWR VPWR _16842_/X sky130_fd_sc_hd__and2_4
XFILLER_111_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19561_ _19450_/A _19507_/B VGND VGND VPWR VPWR _19649_/A sky130_fd_sc_hd__or2_4
XFILLER_77_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13985_ _13985_/A _13983_/X _13985_/C VGND VGND VPWR VPWR _13989_/B sky130_fd_sc_hd__and3_4
X_16773_ _16608_/A VGND VGND VPWR VPWR _16791_/A sky130_fd_sc_hd__buf_2
XANTENNA__20510__A _20510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18187__A _16941_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18512_ _18413_/X _17429_/X _18508_/X _18467_/X _18511_/Y VGND VGND VPWR VPWR _18512_/X
+ sky130_fd_sc_hd__a32o_4
X_12936_ _12943_/A _23465_/Q VGND VGND VPWR VPWR _12936_/X sky130_fd_sc_hd__or2_4
X_15724_ _12766_/X _15722_/X _15724_/C VGND VGND VPWR VPWR _15724_/X sky130_fd_sc_hd__and3_4
XANTENNA__15604__A _13866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19492_ _19480_/A _19491_/X HRDATA[10] _19442_/X VGND VGND VPWR VPWR _19493_/A sky130_fd_sc_hd__o22a_4
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15323__B _23768_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18443_ _18389_/A _18443_/B VGND VGND VPWR VPWR _18443_/X sky130_fd_sc_hd__and2_4
X_12867_ _12867_/A _23689_/Q VGND VGND VPWR VPWR _12869_/B sky130_fd_sc_hd__or2_4
X_15655_ _15654_/X VGND VGND VPWR VPWR _15655_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13124__A _12676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14606_ _13593_/A _14604_/X _14605_/X VGND VGND VPWR VPWR _14606_/X sky130_fd_sc_hd__and3_4
X_11818_ _12156_/A _21183_/A VGND VGND VPWR VPWR _11818_/X sky130_fd_sc_hd__or2_4
X_18374_ _18517_/A VGND VGND VPWR VPWR _18483_/A sky130_fd_sc_hd__buf_2
X_15586_ _13866_/A VGND VGND VPWR VPWR _15610_/A sky130_fd_sc_hd__buf_2
X_12798_ _13343_/A _12798_/B _12798_/C VGND VGND VPWR VPWR _12798_/X sky130_fd_sc_hd__and3_4
XANTENNA__22437__A _20558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18525__B1 _18516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21341__A _21341_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22321__B2 _22284_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14537_ _14372_/A _14533_/X _14536_/X VGND VGND VPWR VPWR _14537_/X sky130_fd_sc_hd__or3_4
XFILLER_109_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17325_ _15380_/A _17323_/Y VGND VGND VPWR VPWR _17326_/B sky130_fd_sc_hd__or2_4
XFILLER_144_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20332__B1 _20714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11749_ _11694_/X _11732_/X _11749_/C VGND VGND VPWR VPWR _11749_/X sky130_fd_sc_hd__or3_4
XFILLER_109_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ _11915_/A _14466_/X _14468_/C VGND VGND VPWR VPWR _14472_/B sky130_fd_sc_hd__and3_4
X_17256_ _17255_/X _17256_/B VGND VGND VPWR VPWR _17256_/X sky130_fd_sc_hd__and2_4
XFILLER_174_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16207_ _13383_/A _16207_/B _16207_/C VGND VGND VPWR VPWR _16239_/B sky130_fd_sc_hd__or3_4
X_13419_ _13455_/A _23269_/Q VGND VGND VPWR VPWR _13419_/X sky130_fd_sc_hd__or2_4
XFILLER_31_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18828__A1 _14844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17187_ _12024_/A _17144_/A _18744_/A _17146_/A VGND VGND VPWR VPWR _17187_/X sky130_fd_sc_hd__o22a_4
X_14399_ _14369_/A _14399_/B VGND VGND VPWR VPWR _14399_/X sky130_fd_sc_hd__or2_4
X_16138_ _16138_/A _16138_/B _16138_/C VGND VGND VPWR VPWR _16138_/X sky130_fd_sc_hd__or3_4
XFILLER_127_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17500__A1 _16768_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22172__A _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13794__A _13952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16069_ _16057_/A _23118_/Q VGND VGND VPWR VPWR _16071_/B sky130_fd_sc_hd__or2_4
XANTENNA__17266__A _16819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16170__A _13408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22388__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21060__B2 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19828_ _19781_/A _19787_/A _19828_/C _19828_/D VGND VGND VPWR VPWR _19828_/X sky130_fd_sc_hd__or4_4
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12203__A _13042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19759_ _19746_/X _19755_/X _19556_/X _19758_/X VGND VGND VPWR VPWR _19759_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20420__A _20895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22770_ _22769_/X VGND VGND VPWR VPWR _22770_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21363__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22560__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21721_ _21541_/X _21720_/X _23694_/Q _21717_/X VGND VGND VPWR VPWR _21721_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13034__A _12570_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24440_ _24445_/CLK _18829_/X HRESETn VGND VGND VPWR VPWR _24440_/Q sky130_fd_sc_hd__dfrtp_4
X_21652_ _21596_/X _21648_/X _23735_/Q _21617_/A VGND VGND VPWR VPWR _23735_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20603_ _20425_/X _20602_/X _24294_/Q _20519_/X VGND VGND VPWR VPWR _20603_/X sky130_fd_sc_hd__o22a_4
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24371_ _24397_/CLK _18955_/Y HRESETn VGND VGND VPWR VPWR _11544_/D sky130_fd_sc_hd__dfstp_4
XANTENNA__12873__A _12873_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21583_ _21582_/X _21578_/X _23773_/Q _21573_/X VGND VGND VPWR VPWR _21583_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16345__A _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23322_ _23294_/CLK _23322_/D VGND VGND VPWR VPWR _14570_/B sky130_fd_sc_hd__dfxtp_4
X_20534_ _20895_/A VGND VGND VPWR VPWR _20534_/X sky130_fd_sc_hd__buf_2
XFILLER_20_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23253_ _23904_/CLK _23253_/D VGND VGND VPWR VPWR _23253_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18819__A1 _17161_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20465_ _20418_/X _20464_/X _24109_/Q _20396_/X VGND VGND VPWR VPWR _20465_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22204_ _22139_/X _22201_/X _15497_/B _22198_/X VGND VGND VPWR VPWR _23426_/D sky130_fd_sc_hd__o22a_4
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20626__A1 _18394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23184_ _23728_/CLK _22599_/X VGND VGND VPWR VPWR _16415_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_165_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20396_ _20396_/A VGND VGND VPWR VPWR _20396_/X sky130_fd_sc_hd__buf_2
X_22135_ _22123_/A VGND VGND VPWR VPWR _22135_/X sky130_fd_sc_hd__buf_2
XFILLER_106_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16080__A _16080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22379__B2 _22373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22066_ _21848_/X _22060_/X _13469_/B _22064_/X VGND VGND VPWR VPWR _23493_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22810__A _17284_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21051__B2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21017_ _21017_/A _21016_/X VGND VGND VPWR VPWR _21017_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__12113__A _16079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21426__A _21455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13770_ _12635_/A _13768_/X _13769_/X VGND VGND VPWR VPWR _13770_/X sky130_fd_sc_hd__and3_4
X_22968_ _22947_/X _22966_/Y _22967_/X VGND VGND VPWR VPWR _22968_/X sky130_fd_sc_hd__and3_4
XANTENNA__21354__A2 _21348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12721_ _12721_/A _23978_/Q VGND VGND VPWR VPWR _12721_/X sky130_fd_sc_hd__or2_4
XFILLER_43_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21919_ _21855_/X _21916_/X _15471_/B _21913_/X VGND VGND VPWR VPWR _23586_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20562__B1 _20306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22899_ _12112_/Y _22885_/X _19909_/X _22898_/X VGND VGND VPWR VPWR _22899_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15440_ _13676_/A _15512_/B VGND VGND VPWR VPWR _15441_/C sky130_fd_sc_hd__or2_4
X_12652_ _12644_/A _12549_/B VGND VGND VPWR VPWR _12653_/C sky130_fd_sc_hd__or2_4
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24202__CLK _24182_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21106__A2 _21104_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22303__B2 _22298_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _11603_/A VGND VGND VPWR VPWR _11604_/A sky130_fd_sc_hd__buf_2
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _13704_/A _24088_/Q VGND VGND VPWR VPWR _15372_/C sky130_fd_sc_hd__or2_4
X_12583_ _12583_/A VGND VGND VPWR VPWR _12949_/A sky130_fd_sc_hd__buf_2
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16255__A _16159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12783__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14322_ _12198_/A _23644_/Q VGND VGND VPWR VPWR _14323_/C sky130_fd_sc_hd__or2_4
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17110_ _17109_/X VGND VGND VPWR VPWR _18198_/A sky130_fd_sc_hd__buf_2
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11534_ _24360_/Q _11533_/X VGND VGND VPWR VPWR _19018_/A sky130_fd_sc_hd__or2_4
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18090_ _17877_/X _17203_/X _17880_/X VGND VGND VPWR VPWR _18090_/X sky130_fd_sc_hd__o21a_4
XFILLER_157_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17041_ _17039_/A VGND VGND VPWR VPWR _17357_/B sky130_fd_sc_hd__inv_2
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ _14656_/A _14251_/X _14252_/X VGND VGND VPWR VPWR _14253_/X sky130_fd_sc_hd__and3_4
XANTENNA__22606__A2 _22601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19566__A HRDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13204_ _13230_/A _13204_/B VGND VGND VPWR VPWR _13204_/X sky130_fd_sc_hd__or2_4
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14184_ _14196_/A _23519_/Q VGND VGND VPWR VPWR _14184_/X sky130_fd_sc_hd__or2_4
XFILLER_125_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13135_ _12721_/A _23783_/Q VGND VGND VPWR VPWR _13135_/X sky130_fd_sc_hd__or2_4
X_18992_ _18978_/X _18991_/X _18978_/X _24366_/Q VGND VGND VPWR VPWR _24366_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14847__A2 _14844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13066_ _13096_/A _13066_/B _13066_/C VGND VGND VPWR VPWR _13072_/B sky130_fd_sc_hd__and3_4
X_17943_ _17943_/A VGND VGND VPWR VPWR _17943_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13119__A _12758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12017_ _16145_/A _12013_/X _12017_/C VGND VGND VPWR VPWR _12018_/B sky130_fd_sc_hd__or3_4
X_17874_ _17873_/X VGND VGND VPWR VPWR _17874_/X sky130_fd_sc_hd__buf_2
XANTENNA__12023__A _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19613_ _19532_/A VGND VGND VPWR VPWR _19613_/X sky130_fd_sc_hd__buf_2
X_16825_ _16686_/X _16822_/Y _16688_/A VGND VGND VPWR VPWR _16825_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__17533__B _17522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12958__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11862__A _13689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19544_ _19888_/B _19629_/A VGND VGND VPWR VPWR _19816_/B sky130_fd_sc_hd__or2_4
XANTENNA__15334__A _15372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16756_ _16755_/X _16756_/B VGND VGND VPWR VPWR _16756_/X sky130_fd_sc_hd__or2_4
XFILLER_65_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13968_ _12502_/A _24000_/Q VGND VGND VPWR VPWR _13969_/C sky130_fd_sc_hd__or2_4
XFILLER_62_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18746__B1 _17816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22542__B2 _22541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15707_ _13306_/A _15703_/X _15707_/C VGND VGND VPWR VPWR _15707_/X sky130_fd_sc_hd__or3_4
XANTENNA__11581__B IRQ[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12919_ _12644_/A _12919_/B VGND VGND VPWR VPWR _12919_/X sky130_fd_sc_hd__or2_4
X_19475_ _20246_/B _19518_/A _19474_/X HRDATA[15] VGND VGND VPWR VPWR _19475_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13899_ _13888_/A VGND VGND VPWR VPWR _14390_/A sky130_fd_sc_hd__buf_2
X_16687_ _16687_/A _16685_/X VGND VGND VPWR VPWR _16688_/A sky130_fd_sc_hd__or2_4
X_18426_ _18405_/X _18410_/Y _18412_/X _18424_/X _18425_/Y VGND VGND VPWR VPWR _18426_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_22_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15638_ _13885_/A _15638_/B VGND VGND VPWR VPWR _15638_/X sky130_fd_sc_hd__or2_4
X_18357_ _17906_/B VGND VGND VPWR VPWR _22990_/B sky130_fd_sc_hd__inv_2
XANTENNA__12693__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15569_ _12435_/A _15569_/B VGND VGND VPWR VPWR _15569_/X sky130_fd_sc_hd__or2_4
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19710__A2 _19848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17308_ _14412_/X _17308_/B VGND VGND VPWR VPWR _17308_/X sky130_fd_sc_hd__or2_4
X_18288_ _18288_/A _18287_/X VGND VGND VPWR VPWR _18288_/Y sky130_fd_sc_hd__nor2_4
XFILLER_30_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22058__B1 _12668_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17239_ _17236_/B VGND VGND VPWR VPWR _17240_/B sky130_fd_sc_hd__inv_2
XFILLER_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20250_ _20308_/A VGND VGND VPWR VPWR _20251_/A sky130_fd_sc_hd__buf_2
XFILLER_157_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17708__B _17381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20415__A _20415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20181_ _24458_/Q IRQ[21] _20180_/X VGND VGND VPWR VPWR _20181_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_7_12_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR _24422_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__14413__A _14412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_75_0_HCLK clkbuf_7_74_0_HCLK/A VGND VGND VPWR VPWR _23392_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_130_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13029__A _12513_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23940_ _23908_/CLK _23940_/D VGND VGND VPWR VPWR _23940_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24488__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23871_ _23101_/CLK _23871_/D VGND VGND VPWR VPWR _23871_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12868__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11772__A _16049_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22822_ _22814_/X _22822_/B VGND VGND VPWR VPWR HWDATA[8] sky130_fd_sc_hd__nor2_4
XFILLER_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24225__CLK _24137_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21336__A2 _21334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22533__B2 _22498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22753_ _22753_/A VGND VGND VPWR VPWR _22753_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21704_ _21600_/X _21677_/A _23701_/Q _21667_/A VGND VGND VPWR VPWR _23701_/D sky130_fd_sc_hd__o22a_4
X_22684_ _22482_/X _22679_/X _14958_/B _22648_/A VGND VGND VPWR VPWR _22684_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24375__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24423_ _24422_/CLK _24423_/D HRESETn VGND VGND VPWR VPWR _20579_/A sky130_fd_sc_hd__dfrtp_4
X_21635_ _21565_/X _21634_/X _23748_/Q _21631_/X VGND VGND VPWR VPWR _23748_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22297__B1 _13199_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13699__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24354_ _24388_/CLK _24354_/D HRESETn VGND VGND VPWR VPWR _11528_/A sky130_fd_sc_hd__dfstp_4
X_21566_ _21542_/A VGND VGND VPWR VPWR _21566_/X sky130_fd_sc_hd__buf_2
XFILLER_21_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22805__A _15048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23305_ _23561_/CLK _22377_/X VGND VGND VPWR VPWR _23305_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20517_ _24426_/Q _20427_/X _24458_/Q _20471_/X VGND VGND VPWR VPWR _20517_/X sky130_fd_sc_hd__o22a_4
X_24285_ _24292_/CLK _24285_/D HRESETn VGND VGND VPWR VPWR _19234_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21497_ _21275_/X _21492_/X _23814_/Q _21496_/X VGND VGND VPWR VPWR _21497_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12108__A _12108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23236_ _23303_/CLK _22516_/X VGND VGND VPWR VPWR _15704_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_10_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20448_ _20448_/A _20318_/B VGND VGND VPWR VPWR _20448_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__20325__A _20267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15419__A _11932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11947__A _11943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21272__B2 _21264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23167_ _23229_/CLK _22623_/X VGND VGND VPWR VPWR _23167_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_133_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20379_ _20302_/X _20378_/X _24113_/Q _20225_/X VGND VGND VPWR VPWR _24113_/D sky130_fd_sc_hd__o22a_4
X_22118_ _22118_/A VGND VGND VPWR VPWR _22118_/X sky130_fd_sc_hd__buf_2
X_23098_ _23098_/CLK _23098_/D VGND VGND VPWR VPWR _14604_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22049_ _21819_/X _22046_/X _23505_/Q _22043_/X VGND VGND VPWR VPWR _22049_/X sky130_fd_sc_hd__o22a_4
X_14940_ _14925_/X _14940_/B _14939_/X VGND VGND VPWR VPWR _14940_/X sky130_fd_sc_hd__and3_4
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14871_ _12473_/A _14871_/B VGND VGND VPWR VPWR _14871_/X sky130_fd_sc_hd__or2_4
XFILLER_21_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16451__A1 _11858_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11682__A _11682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16610_ _16775_/A VGND VGND VPWR VPWR _16611_/A sky130_fd_sc_hd__buf_2
X_13822_ _14325_/A _13896_/B VGND VGND VPWR VPWR _13822_/X sky130_fd_sc_hd__or2_4
X_17590_ _17120_/Y _17968_/B _17583_/A _17589_/X VGND VGND VPWR VPWR _17590_/X sky130_fd_sc_hd__o22a_4
XFILLER_169_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22524__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13753_ _13753_/A _23614_/Q VGND VGND VPWR VPWR _13753_/X sky130_fd_sc_hd__or2_4
X_16541_ _12001_/X _16541_/B _16541_/C VGND VGND VPWR VPWR _16542_/C sky130_fd_sc_hd__and3_4
XFILLER_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12704_ _12704_/A _12704_/B _12703_/X VGND VGND VPWR VPWR _12708_/B sky130_fd_sc_hd__and3_4
XANTENNA__13017__A1 _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19260_ _24307_/Q _19256_/B _19258_/Y VGND VGND VPWR VPWR _24307_/D sky130_fd_sc_hd__o21a_4
X_16472_ _16490_/A _16412_/B VGND VGND VPWR VPWR _16472_/X sky130_fd_sc_hd__or2_4
X_13684_ _12299_/A _13684_/B _13684_/C VGND VGND VPWR VPWR _13684_/X sky130_fd_sc_hd__and3_4
XFILLER_44_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18211_ _18187_/X _19400_/A _18033_/X _18210_/X VGND VGND VPWR VPWR _18211_/X sky130_fd_sc_hd__o22a_4
X_12635_ _12635_/A VGND VGND VPWR VPWR _12944_/A sky130_fd_sc_hd__buf_2
X_15423_ _15423_/A _15487_/B VGND VGND VPWR VPWR _15424_/C sky130_fd_sc_hd__or2_4
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14765__A1 _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19191_ _19146_/X VGND VGND VPWR VPWR _19191_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18142_ _18013_/C _18013_/B _18013_/C _18013_/B VGND VGND VPWR VPWR _18142_/X sky130_fd_sc_hd__a2bb2o_4
X_15354_ _11752_/A _15354_/B _15354_/C VGND VGND VPWR VPWR _15362_/B sky130_fd_sc_hd__or3_4
X_12566_ _12493_/A _12566_/B _12566_/C VGND VGND VPWR VPWR _12571_/B sky130_fd_sc_hd__and3_4
XFILLER_15_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22715__A _22708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14305_ _15393_/A _23964_/Q VGND VGND VPWR VPWR _14306_/C sky130_fd_sc_hd__or2_4
X_11517_ _11516_/X VGND VGND VPWR VPWR _11518_/B sky130_fd_sc_hd__inv_2
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18073_ _18072_/X VGND VGND VPWR VPWR _18073_/Y sky130_fd_sc_hd__inv_2
X_15285_ _14149_/A _15285_/B _15284_/X VGND VGND VPWR VPWR _15289_/B sky130_fd_sc_hd__and3_4
X_12497_ _12497_/A VGND VGND VPWR VPWR _12498_/A sky130_fd_sc_hd__buf_2
XANTENNA__12018__A _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16713__A _16713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17024_ _17024_/A VGND VGND VPWR VPWR _17024_/X sky130_fd_sc_hd__buf_2
X_14236_ _14665_/A _23839_/Q VGND VGND VPWR VPWR _14237_/C sky130_fd_sc_hd__or2_4
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20235__A _20234_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11857__A _11857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14167_ _12425_/A _14167_/B _14167_/C VGND VGND VPWR VPWR _14167_/X sky130_fd_sc_hd__and3_4
XANTENNA__15329__A _13695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22460__B1 _23264_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13118_ _13096_/A _13118_/B _13118_/C VGND VGND VPWR VPWR _13122_/B sky130_fd_sc_hd__and3_4
X_18975_ _24368_/Q _11542_/B _18948_/B VGND VGND VPWR VPWR _18975_/Y sky130_fd_sc_hd__a21oi_4
X_14098_ _14138_/A _23743_/Q VGND VGND VPWR VPWR _14098_/X sky130_fd_sc_hd__or2_4
XANTENNA__22450__A _22438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13049_ _13049_/A VGND VGND VPWR VPWR _13049_/Y sky130_fd_sc_hd__inv_2
X_17926_ _17878_/A VGND VGND VPWR VPWR _18126_/A sky130_fd_sc_hd__buf_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24248__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21066__A _21033_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17857_ _17837_/X _17205_/X _17838_/X _17207_/X VGND VGND VPWR VPWR _17857_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12688__A _11881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16808_ _16656_/A _16806_/X _16807_/X VGND VGND VPWR VPWR _16808_/X sky130_fd_sc_hd__and3_4
XFILLER_82_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17788_ _24160_/Q _17008_/Y _16999_/B VGND VGND VPWR VPWR _17788_/Y sky130_fd_sc_hd__o21ai_4
X_19527_ _19624_/A VGND VGND VPWR VPWR _19528_/A sky130_fd_sc_hd__inv_2
XANTENNA__15999__A _15998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16739_ _12061_/A _16737_/X _16738_/X VGND VGND VPWR VPWR _16739_/X sky130_fd_sc_hd__and3_4
XANTENNA__18375__A _18483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19458_ _24165_/Q _19454_/X HRDATA[17] _19457_/X VGND VGND VPWR VPWR _19458_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__17942__A1 _17875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18409_ _18409_/A _18409_/B _18409_/C _18408_/X VGND VGND VPWR VPWR _18409_/X sky130_fd_sc_hd__or4_4
XANTENNA__15511__B _15511_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19389_ _19377_/A VGND VGND VPWR VPWR _19389_/X sky130_fd_sc_hd__buf_2
X_21420_ _21184_/A _21420_/B _21134_/C _21134_/D VGND VGND VPWR VPWR _21420_/X sky130_fd_sc_hd__or4_4
XFILLER_72_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19695__A1 _19797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14127__B _23935_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21351_ _21285_/X _21348_/X _23906_/Q _21345_/X VGND VGND VPWR VPWR _23906_/D sky130_fd_sc_hd__o22a_4
XFILLER_120_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20302_ _20533_/A VGND VGND VPWR VPWR _20302_/X sky130_fd_sc_hd__buf_2
XFILLER_107_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24070_ _24102_/CLK _24070_/D VGND VGND VPWR VPWR _24070_/Q sky130_fd_sc_hd__dfxtp_4
X_21282_ _21280_/X _21281_/X _23940_/Q _21276_/X VGND VGND VPWR VPWR _23940_/D sky130_fd_sc_hd__o22a_4
XFILLER_162_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13192__B1 _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23021_ _18272_/X _23003_/B VGND VGND VPWR VPWR _23022_/C sky130_fd_sc_hd__or2_4
X_20233_ _20217_/D VGND VGND VPWR VPWR _20233_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15239__A _12336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14143__A _12287_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20164_ IRQ[11] VGND VGND VPWR VPWR _20164_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17454__A _12097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20095_ _17820_/X _17817_/X _18887_/X _20095_/D VGND VGND VPWR VPWR _20095_/X sky130_fd_sc_hd__or4_4
XANTENNA__21557__A2 _21554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23923_ _23764_/CLK _23923_/D VGND VGND VPWR VPWR _23923_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12598__A _12925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_5_0_HCLK clkbuf_6_2_0_HCLK/X VGND VGND VPWR VPWR _24294_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_45_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23854_ _24078_/CLK _23854_/D VGND VGND VPWR VPWR _15989_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22506__B2 _22505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22805_ _15048_/X _22804_/X VGND VGND VPWR VPWR HWDATA[0] sky130_fd_sc_hd__nor2_4
X_23785_ _23561_/CLK _23785_/D VGND VGND VPWR VPWR _23785_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20517__B1 _24458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20997_ _22846_/B _20313_/X _20780_/X _20996_/Y VGND VGND VPWR VPWR _20997_/X sky130_fd_sc_hd__a211o_4
XANTENNA__19383__B1 _18148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15702__A _13304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22736_ _22945_/A HREADY VGND VGND VPWR VPWR _22736_/X sky130_fd_sc_hd__and2_4
XFILLER_53_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23765__CLK _23904_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22667_ _22452_/X _22665_/X _15826_/B _22662_/X VGND VGND VPWR VPWR _23139_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14318__A _15406_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12420_ _12320_/Y _12419_/X VGND VGND VPWR VPWR _12423_/A sky130_fd_sc_hd__and2_4
X_24406_ _24422_/CLK _24406_/D HRESETn VGND VGND VPWR VPWR _24406_/Q sky130_fd_sc_hd__dfrtp_4
X_21618_ _21536_/X _21613_/X _16391_/B _21617_/X VGND VGND VPWR VPWR _23760_/D sky130_fd_sc_hd__o22a_4
XFILLER_139_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22598_ _22598_/A VGND VGND VPWR VPWR _22598_/X sky130_fd_sc_hd__buf_2
XFILLER_139_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12351_ _12387_/A _12349_/X _12350_/X VGND VGND VPWR VPWR _12351_/X sky130_fd_sc_hd__and3_4
X_24337_ _24277_/CLK _24337_/D HRESETn VGND VGND VPWR VPWR _19158_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21493__B2 _21489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21549_ _21549_/A VGND VGND VPWR VPWR _21549_/X sky130_fd_sc_hd__buf_2
XFILLER_166_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15070_ _14773_/A VGND VGND VPWR VPWR _15095_/A sky130_fd_sc_hd__buf_2
X_12282_ _12311_/A VGND VGND VPWR VPWR _13139_/A sky130_fd_sc_hd__buf_2
X_24268_ _24495_/CLK _24268_/D HRESETn VGND VGND VPWR VPWR _24268_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20055__A _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20048__A2 _20031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14021_ _13700_/A _23360_/Q VGND VGND VPWR VPWR _14023_/B sky130_fd_sc_hd__or2_4
XFILLER_88_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11677__A _13530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19989__A2 _19983_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15149__A _14988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23219_ _23379_/CLK _23219_/D VGND VGND VPWR VPWR _12124_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23145__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24199_ _23671_/CLK _19772_/Y HRESETn VGND VGND VPWR VPWR _11664_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14053__A _13705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21796__A2 _21791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14988__A _14988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24339__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17364__A _15653_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13892__A _14385_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18760_ _18757_/X _18759_/X _18506_/A VGND VGND VPWR VPWR _18773_/A sky130_fd_sc_hd__a21o_4
X_15972_ _11889_/X _16038_/B VGND VGND VPWR VPWR _15972_/X sky130_fd_sc_hd__or2_4
XANTENNA__23085__B _23084_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17711_ _17711_/A VGND VGND VPWR VPWR _17712_/A sky130_fd_sc_hd__inv_2
X_14923_ _14919_/A _23766_/Q VGND VGND VPWR VPWR _14923_/X sky130_fd_sc_hd__or2_4
X_18691_ _17975_/X _17943_/Y _17944_/X _18690_/Y VGND VGND VPWR VPWR _18691_/X sky130_fd_sc_hd__a211o_4
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17642_ _17642_/A _17642_/B _17642_/C VGND VGND VPWR VPWR _17642_/X sky130_fd_sc_hd__and3_4
XFILLER_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14854_ _14094_/A _14852_/X _14854_/C VGND VGND VPWR VPWR _14854_/X sky130_fd_sc_hd__and3_4
XFILLER_91_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13805_ _12445_/A _13803_/X _13805_/C VGND VGND VPWR VPWR _13805_/X sky130_fd_sc_hd__and3_4
X_17573_ _17572_/X VGND VGND VPWR VPWR _18099_/A sky130_fd_sc_hd__inv_2
X_14785_ _13717_/A VGND VGND VPWR VPWR _14786_/A sky130_fd_sc_hd__buf_2
XFILLER_63_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11997_ _12103_/A _11828_/B VGND VGND VPWR VPWR _11997_/X sky130_fd_sc_hd__or2_4
X_19312_ _19230_/A _19313_/A _19311_/Y VGND VGND VPWR VPWR _24281_/D sky130_fd_sc_hd__o21a_4
X_16524_ _16452_/Y _16521_/X VGND VGND VPWR VPWR _16525_/A sky130_fd_sc_hd__or2_4
X_13736_ _13744_/A _13736_/B VGND VGND VPWR VPWR _13736_/X sky130_fd_sc_hd__or2_4
XANTENNA__21181__B1 _23990_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19243_ _24294_/Q _19243_/B VGND VGND VPWR VPWR _19244_/B sky130_fd_sc_hd__and2_4
X_16455_ _11702_/X _16455_/B _16455_/C VGND VGND VPWR VPWR _16455_/X sky130_fd_sc_hd__and3_4
X_13667_ _15406_/A _13757_/B VGND VGND VPWR VPWR _13667_/X sky130_fd_sc_hd__or2_4
XANTENNA__13132__A _13276_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15406_ _15406_/A _15477_/B VGND VGND VPWR VPWR _15408_/B sky130_fd_sc_hd__or2_4
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12618_ _12646_/A _12618_/B VGND VGND VPWR VPWR _12618_/X sky130_fd_sc_hd__or2_4
X_19174_ _19155_/A _19155_/B _19173_/Y VGND VGND VPWR VPWR _19174_/X sky130_fd_sc_hd__o21a_4
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13598_ _12450_/X VGND VGND VPWR VPWR _13957_/A sky130_fd_sc_hd__buf_2
X_16386_ _16309_/X _16383_/X _16385_/Y VGND VGND VPWR VPWR _16527_/A sky130_fd_sc_hd__a21o_4
XANTENNA__22445__A _22433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18125_ _17810_/X _18125_/B VGND VGND VPWR VPWR _18125_/X sky130_fd_sc_hd__or2_4
X_12549_ _12895_/A _12549_/B VGND VGND VPWR VPWR _12549_/X sky130_fd_sc_hd__or2_4
XANTENNA__21484__B2 _21482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15337_ _11697_/A _15337_/B _15337_/C VGND VGND VPWR VPWR _15337_/X sky130_fd_sc_hd__and3_4
XANTENNA__22681__B1 _14743_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12971__A _12971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18056_ _17111_/X _18653_/B _17224_/X _18055_/X VGND VGND VPWR VPWR _18056_/X sky130_fd_sc_hd__a211o_4
X_15268_ _14269_/A _23992_/Q VGND VGND VPWR VPWR _15268_/X sky130_fd_sc_hd__or2_4
X_17007_ _17905_/A _17906_/B _17906_/C _16994_/B VGND VGND VPWR VPWR _17009_/B sky130_fd_sc_hd__or4_4
XANTENNA__19754__A _19705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14910__A1 _15281_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14219_ _14248_/A _23551_/Q VGND VGND VPWR VPWR _14220_/C sky130_fd_sc_hd__or2_4
XANTENNA__15059__A _12322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15199_ _15198_/X _15136_/B VGND VGND VPWR VPWR _15199_/X sky130_fd_sc_hd__or2_4
XANTENNA__21787__A2 _21784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22180__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14898__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17274__A _17274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18958_ _18957_/X VGND VGND VPWR VPWR _18959_/A sky130_fd_sc_hd__buf_2
XFILLER_112_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17909_ _17909_/A VGND VGND VPWR VPWR _17909_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18889_ _17817_/X _18889_/B _18888_/X VGND VGND VPWR VPWR _20274_/A sky130_fd_sc_hd__or3_4
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13307__A _13307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20920_ _19756_/Y _20873_/A _20917_/B _20843_/B VGND VGND VPWR VPWR _20920_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21524__A _21549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20851_ _20755_/X _20850_/X _11522_/A _20708_/X VGND VGND VPWR VPWR _20851_/X sky130_fd_sc_hd__o22a_4
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15522__A _15439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23570_ _23204_/CLK _21948_/X VGND VGND VPWR VPWR _23570_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20782_ _20315_/A VGND VGND VPWR VPWR _20782_/X sky130_fd_sc_hd__buf_2
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22521_ _22459_/X _22515_/X _23232_/Q _22519_/X VGND VGND VPWR VPWR _22521_/X sky130_fd_sc_hd__o22a_4
XFILLER_161_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14138__A _14138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18833__A _12061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13042__A _13042_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22452_ _20692_/A VGND VGND VPWR VPWR _22452_/X sky130_fd_sc_hd__buf_2
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21403_ _21287_/X _21398_/X _15638_/B _21402_/X VGND VGND VPWR VPWR _21403_/X sky130_fd_sc_hd__o22a_4
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22383_ _22376_/A VGND VGND VPWR VPWR _22383_/X sky130_fd_sc_hd__buf_2
XANTENNA__23168__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12881__A _12881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16353__A _13414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24122_ _23416_/CLK _24122_/D HRESETn VGND VGND VPWR VPWR _22784_/A sky130_fd_sc_hd__dfrtp_4
X_21334_ _21341_/A VGND VGND VPWR VPWR _21334_/X sky130_fd_sc_hd__buf_2
XANTENNA__15154__A1 _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21227__B2 _21223_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24053_ _23203_/CLK _21079_/X VGND VGND VPWR VPWR _24053_/Q sky130_fd_sc_hd__dfxtp_4
X_21265_ _21263_/X _21257_/X _12618_/B _21264_/X VGND VGND VPWR VPWR _23947_/D sky130_fd_sc_hd__o22a_4
XFILLER_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24389__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21778__A2 _21777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23004_ _22978_/X _23001_/Y _23004_/C VGND VGND VPWR VPWR _23004_/X sky130_fd_sc_hd__and3_4
X_20216_ _22798_/A _11647_/B _16936_/X _20216_/D VGND VGND VPWR VPWR _20217_/D sky130_fd_sc_hd__or4_4
XFILLER_131_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21196_ _20395_/X _21191_/X _16422_/B _21195_/X VGND VGND VPWR VPWR _23984_/D sky130_fd_sc_hd__o22a_4
XFILLER_173_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20147_ _11636_/A _20147_/B VGND VGND VPWR VPWR _20147_/X sky130_fd_sc_hd__and2_4
XFILLER_104_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_45_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14601__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22727__A1 _20860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22727__B2 _22726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15416__B _15473_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20738__B1 _20538_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20078_ _20077_/X VGND VGND VPWR VPWR _24142_/D sky130_fd_sc_hd__inv_2
XFILLER_46_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13217__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23906_ _23587_/CLK _23906_/D VGND VGND VPWR VPWR _23906_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11920_ _16148_/A VGND VGND VPWR VPWR _16713_/A sky130_fd_sc_hd__buf_2
XFILLER_100_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21434__A _21441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11851_ _11671_/X _11809_/X _11850_/X VGND VGND VPWR VPWR _11851_/X sky130_fd_sc_hd__and3_4
XFILLER_79_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23837_ _23518_/CLK _23837_/D VGND VGND VPWR VPWR _13839_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15432__A _12191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11960__A _11960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _15395_/A _14570_/B VGND VGND VPWR VPWR _14572_/B sky130_fd_sc_hd__or2_4
XPHY_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _12354_/A VGND VGND VPWR VPWR _13092_/A sky130_fd_sc_hd__buf_2
X_23768_ _23770_/CLK _21595_/X VGND VGND VPWR VPWR _23768_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0_0_HCLK clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _12957_/A VGND VGND VPWR VPWR _13521_/X sky130_fd_sc_hd__buf_2
XPHY_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22719_ _22705_/A VGND VGND VPWR VPWR _22719_/X sky130_fd_sc_hd__buf_2
XPHY_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23699_ _23760_/CLK _21714_/X VGND VGND VPWR VPWR _23699_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14048__A _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13452_ _12890_/A _13448_/X _13452_/C VGND VGND VPWR VPWR _13452_/X sky130_fd_sc_hd__or3_4
X_16240_ _16239_/X VGND VGND VPWR VPWR _16240_/X sky130_fd_sc_hd__buf_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22265__A _22258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ _12373_/X _23724_/Q VGND VGND VPWR VPWR _12405_/B sky130_fd_sc_hd__or2_4
XANTENNA__13887__A _15595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16171_ _16215_/A _23373_/Q VGND VGND VPWR VPWR _16171_/X sky130_fd_sc_hd__or2_4
X_13383_ _13383_/A _13363_/X _13383_/C VGND VGND VPWR VPWR _13417_/B sky130_fd_sc_hd__or3_4
XANTENNA__21466__B2 _21431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12791__A _12773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ _13717_/A VGND VGND VPWR VPWR _15324_/A sky130_fd_sc_hd__buf_2
XFILLER_51_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15122_ _14140_/A _15122_/B VGND VGND VPWR VPWR _15122_/X sky130_fd_sc_hd__or2_4
XANTENNA__17078__B _17077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_127_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR _24073_/CLK sky130_fd_sc_hd__clkbuf_1
X_19930_ _19921_/X _24175_/Q _19925_/X _20380_/B VGND VGND VPWR VPWR _24175_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20216__C _16936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15053_ _14773_/A VGND VGND VPWR VPWR _15075_/A sky130_fd_sc_hd__buf_2
XANTENNA__21218__B2 _21216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12265_ _13016_/A VGND VGND VPWR VPWR _12882_/A sky130_fd_sc_hd__buf_2
XFILLER_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21769__A2 _21763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14004_ _12287_/A _13999_/X _14004_/C VGND VGND VPWR VPWR _14004_/X sky130_fd_sc_hd__or3_4
XANTENNA_clkbuf_3_6_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21609__A _21624_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19861_ _19612_/A _19895_/C VGND VGND VPWR VPWR _19861_/X sky130_fd_sc_hd__or2_4
XFILLER_134_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12196_ _13630_/A VGND VGND VPWR VPWR _15444_/A sky130_fd_sc_hd__buf_2
XANTENNA__24173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18812_ _13567_/X _18810_/X _24453_/Q _18811_/X VGND VGND VPWR VPWR _18812_/X sky130_fd_sc_hd__o22a_4
XFILLER_150_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19792_ HRDATA[16] VGND VGND VPWR VPWR _22737_/A sky130_fd_sc_hd__buf_2
XFILLER_95_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22718__B2 _22712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18743_ _18667_/X _18742_/X _24470_/Q _18667_/X VGND VGND VPWR VPWR _18743_/X sky130_fd_sc_hd__a2bb2o_4
X_15955_ _13462_/A VGND VGND VPWR VPWR _15956_/A sky130_fd_sc_hd__buf_2
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14230__B _23615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13127__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14906_ _14155_/A _23862_/Q VGND VGND VPWR VPWR _14907_/C sky130_fd_sc_hd__or2_4
XFILLER_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18674_ _18674_/A _18674_/B _18674_/C VGND VGND VPWR VPWR _18675_/B sky130_fd_sc_hd__and3_4
X_15886_ _13521_/X _15884_/X _15885_/X VGND VGND VPWR VPWR _15887_/C sky130_fd_sc_hd__and3_4
X_17625_ _18744_/A _17346_/B VGND VGND VPWR VPWR _17626_/A sky130_fd_sc_hd__or2_4
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14837_ _14657_/A _14753_/B VGND VGND VPWR VPWR _14839_/B sky130_fd_sc_hd__or2_4
XANTENNA__12966__A _12942_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11870__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15342__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17556_ _16309_/X VGND VGND VPWR VPWR _17556_/Y sky130_fd_sc_hd__inv_2
X_14768_ _15321_/A VGND VGND VPWR VPWR _14769_/A sky130_fd_sc_hd__buf_2
XFILLER_32_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16507_ _16507_/A _16505_/X _16507_/C VGND VGND VPWR VPWR _16511_/B sky130_fd_sc_hd__and3_4
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13719_ _13719_/A VGND VGND VPWR VPWR _13720_/A sky130_fd_sc_hd__buf_2
XANTENNA__20901__B1 _20512_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17487_ _12680_/X _17487_/B VGND VGND VPWR VPWR _17487_/X sky130_fd_sc_hd__and2_4
XFILLER_147_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14699_ _15649_/A _14699_/B _14699_/C VGND VGND VPWR VPWR _14699_/X sky130_fd_sc_hd__or3_4
XFILLER_60_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19226_ _24129_/Q _19226_/B VGND VGND VPWR VPWR _19321_/A sky130_fd_sc_hd__and2_4
X_16438_ _16112_/A _16438_/B VGND VGND VPWR VPWR _16440_/B sky130_fd_sc_hd__or2_4
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22175__A _22208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19157_ _24336_/Q _19157_/B VGND VGND VPWR VPWR _19158_/B sky130_fd_sc_hd__and2_4
XANTENNA__21457__B2 _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16369_ _16362_/X _16365_/X _16369_/C VGND VGND VPWR VPWR _16369_/X sky130_fd_sc_hd__or3_4
XFILLER_117_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18108_ _24155_/Q _18111_/C _16994_/B VGND VGND VPWR VPWR _23043_/B sky130_fd_sc_hd__o21a_4
XFILLER_173_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19088_ _11523_/B VGND VGND VPWR VPWR _19088_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22903__A _22884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18039_ _18674_/A _18039_/B VGND VGND VPWR VPWR _18042_/C sky130_fd_sc_hd__nor2_4
XANTENNA__12206__A _12687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16901__A _16901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21050_ _20509_/X _21045_/X _12647_/B _21049_/X VGND VGND VPWR VPWR _21050_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20001_ _19992_/X _17904_/X _19998_/X _20000_/X VGND VGND VPWR VPWR _20001_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15517__A _15517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14421__A _14421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22709__B2 _22705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14140__B _23615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22185__A2 _22180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19586__B1 HRDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13037__A _11881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21952_ _21824_/X _21946_/X _16267_/B _21950_/X VGND VGND VPWR VPWR _23567_/D sky130_fd_sc_hd__o22a_4
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21932__A2 _21930_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20903_ _24410_/Q _20427_/A _24442_/Q _20704_/X VGND VGND VPWR VPWR _20903_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21883_ _21313_/A VGND VGND VPWR VPWR _21883_/X sky130_fd_sc_hd__buf_2
XANTENNA__12876__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11780__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23622_ _24102_/CLK _23622_/D VGND VGND VPWR VPWR _13388_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20834_ _18590_/X _20675_/X _20780_/X _20833_/Y VGND VGND VPWR VPWR _20834_/X sky130_fd_sc_hd__a211o_4
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18010__B1 _18009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21696__A1 _21584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23553_ _23744_/CLK _23553_/D VGND VGND VPWR VPWR _15540_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21696__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20765_ _20765_/A VGND VGND VPWR VPWR _20765_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22504_ _22430_/X _22501_/X _12303_/B _22498_/X VGND VGND VPWR VPWR _23244_/D sky130_fd_sc_hd__o22a_4
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23484_ _23323_/CLK _22079_/X VGND VGND VPWR VPWR _23484_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20696_ _20845_/A VGND VGND VPWR VPWR _20700_/A sky130_fd_sc_hd__buf_2
XFILLER_126_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22435_ _20530_/A VGND VGND VPWR VPWR _22435_/X sky130_fd_sc_hd__buf_2
XFILLER_109_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16083__A _16187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21999__A2 _21996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22366_ _22366_/A VGND VGND VPWR VPWR _22366_/X sky130_fd_sc_hd__buf_2
XANTENNA__22813__A _22799_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24105_ _23337_/CLK _20560_/X VGND VGND VPWR VPWR _24105_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21317_ _21317_/A VGND VGND VPWR VPWR _21317_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22297_ _22127_/X _22294_/X _13199_/B _22291_/X VGND VGND VPWR VPWR _23367_/D sky130_fd_sc_hd__o22a_4
XFILLER_11_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23953__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24036_ _23908_/CLK _24036_/D VGND VGND VPWR VPWR _24036_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12050_ _16744_/A VGND VGND VPWR VPWR _12051_/A sky130_fd_sc_hd__buf_2
X_21248_ _21247_/X _21245_/X _23954_/Q _21240_/X VGND VGND VPWR VPWR _23954_/D sky130_fd_sc_hd__o22a_4
XFILLER_117_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14331__A _14331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21179_ _20959_/X _21176_/X _23992_/Q _21173_/X VGND VGND VPWR VPWR _21179_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24309__CLK _24342_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15146__B _15146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15740_ _11755_/X _15736_/X _15739_/X VGND VGND VPWR VPWR _15740_/X sky130_fd_sc_hd__or3_4
XFILLER_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12952_ _12940_/A _24073_/Q VGND VGND VPWR VPWR _12952_/X sky130_fd_sc_hd__or2_4
XANTENNA__20187__A1 _24464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14985__B _23253_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11903_ _13427_/A VGND VGND VPWR VPWR _11903_/X sky130_fd_sc_hd__buf_2
X_15671_ _13300_/A _23684_/Q VGND VGND VPWR VPWR _15673_/B sky130_fd_sc_hd__or2_4
X_12883_ _13483_/A _12857_/X _12866_/X _12874_/X _12882_/X VGND VGND VPWR VPWR _12883_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12786__A _13343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19329__B1 _17048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11690__A _11689_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17410_ _17410_/A VGND VGND VPWR VPWR _17439_/B sky130_fd_sc_hd__inv_2
X_14622_ _14656_/A VGND VGND VPWR VPWR _14693_/A sky130_fd_sc_hd__buf_2
X_11834_ _11834_/A _11834_/B _11833_/X VGND VGND VPWR VPWR _11838_/B sky130_fd_sc_hd__and3_4
XFILLER_45_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18390_ _18198_/X _18411_/B _18265_/X _18389_/X VGND VGND VPWR VPWR _18390_/X sky130_fd_sc_hd__a211o_4
XFILLER_73_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17341_/A _17341_/B VGND VGND VPWR VPWR _17341_/X sky130_fd_sc_hd__and2_4
XFILLER_92_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21687__B2 _21681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14553_ _12434_/A _14618_/B VGND VGND VPWR VPWR _14553_/X sky130_fd_sc_hd__or2_4
X_11765_ _11762_/X _11763_/X _11765_/C VGND VGND VPWR VPWR _11765_/X sky130_fd_sc_hd__and3_4
XPHY_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _12651_/A VGND VGND VPWR VPWR _13534_/A sky130_fd_sc_hd__buf_2
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17272_ _14412_/X VGND VGND VPWR VPWR _17272_/X sky130_fd_sc_hd__buf_2
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14484_ _12372_/A _14484_/B VGND VGND VPWR VPWR _14484_/X sky130_fd_sc_hd__or2_4
X_11696_ _13694_/A VGND VGND VPWR VPWR _11697_/A sky130_fd_sc_hd__buf_2
XANTENNA__20508__A _22117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19011_ _18993_/X _19008_/X _19010_/X _19004_/A VGND VGND VPWR VPWR _24363_/D sky130_fd_sc_hd__a2bb2o_4
X_16223_ _16181_/X _23117_/Q VGND VGND VPWR VPWR _16223_/X sky130_fd_sc_hd__or2_4
X_13435_ _12889_/A VGND VGND VPWR VPWR _13474_/A sky130_fd_sc_hd__buf_2
XANTENNA__21439__B2 _21438_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22100__A2 _22099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13366_ _13410_/A _13366_/B _13366_/C VGND VGND VPWR VPWR _13366_/X sky130_fd_sc_hd__and3_4
X_16154_ _16157_/A _16224_/B VGND VGND VPWR VPWR _16155_/C sky130_fd_sc_hd__or2_4
XFILLER_155_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15105_ _15081_/A _15105_/B _15105_/C VGND VGND VPWR VPWR _15106_/C sky130_fd_sc_hd__and3_4
X_12317_ _11864_/A _12316_/X VGND VGND VPWR VPWR _12317_/X sky130_fd_sc_hd__and2_4
X_13297_ _13320_/A _13297_/B VGND VGND VPWR VPWR _13297_/X sky130_fd_sc_hd__or2_4
X_16085_ _11671_/X _16085_/B _16085_/C VGND VGND VPWR VPWR _16085_/X sky130_fd_sc_hd__and3_4
X_19913_ _19913_/A VGND VGND VPWR VPWR _20867_/A sky130_fd_sc_hd__buf_2
X_15036_ _11931_/A _15036_/B _15036_/C VGND VGND VPWR VPWR _15036_/X sky130_fd_sc_hd__or3_4
X_12248_ _11967_/A VGND VGND VPWR VPWR _14450_/A sky130_fd_sc_hd__buf_2
XANTENNA__11865__A _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24372__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19844_ _19890_/B _19843_/X VGND VGND VPWR VPWR _19844_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__20414__A2 _20304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15337__A _11697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21611__B2 _21610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12179_ _11671_/X _12147_/X _12178_/X VGND VGND VPWR VPWR _12180_/A sky130_fd_sc_hd__and3_4
XFILLER_25_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14241__A _14656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19775_ _19773_/X _19518_/X _19774_/X _19638_/X VGND VGND VPWR VPWR _19775_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15056__B _23733_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16987_ _16987_/A _16986_/X VGND VGND VPWR VPWR _16988_/B sky130_fd_sc_hd__or2_4
XFILLER_27_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19568__B1 _19519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20897__B _20339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18726_ _18625_/X _20155_/A _20154_/A _18624_/X VGND VGND VPWR VPWR _24471_/D sky130_fd_sc_hd__o22a_4
X_15938_ _15944_/A _23278_/Q VGND VGND VPWR VPWR _15941_/B sky130_fd_sc_hd__or2_4
XFILLER_49_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21914__A2 _21909_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14895__B _14895_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18657_ _18506_/X _18649_/Y _18650_/X _18009_/X _18656_/X VGND VGND VPWR VPWR _18657_/X
+ sky130_fd_sc_hd__a32o_4
X_15869_ _13546_/A _15869_/B VGND VGND VPWR VPWR _15870_/C sky130_fd_sc_hd__or2_4
XANTENNA__12696__A _12696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16168__A _16163_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18791__A1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15072__A _15080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17608_ _17607_/X VGND VGND VPWR VPWR _17637_/B sky130_fd_sc_hd__inv_2
XFILLER_24_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18588_ _18557_/A _18586_/X _17792_/X _18587_/X VGND VGND VPWR VPWR _18589_/A sky130_fd_sc_hd__a211o_4
XANTENNA__21127__B1 _14716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10_0_HCLK_A clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17539_ _17539_/A _17467_/B VGND VGND VPWR VPWR _17539_/X sky130_fd_sc_hd__or2_4
XANTENNA__21678__B2 _21674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18543__A1 _18467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18383__A _17187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15800__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20550_ _20539_/X _20548_/X _24329_/Q _20549_/X VGND VGND VPWR VPWR _20550_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21521__B _21370_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_9_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__20418__A _20533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19209_ _19138_/B VGND VGND VPWR VPWR _19209_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22627__B1 _14362_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20481_ _20255_/A VGND VGND VPWR VPWR _20481_/X sky130_fd_sc_hd__buf_2
XANTENNA__14416__A _14334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22220_ _22167_/X _22215_/X _14891_/B _22184_/A VGND VGND VPWR VPWR _23414_/D sky130_fd_sc_hd__o22a_4
XFILLER_164_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22151_ _20840_/A VGND VGND VPWR VPWR _22151_/X sky130_fd_sc_hd__buf_2
XFILLER_156_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21102_ _20509_/X _21097_/X _12608_/B _21101_/X VGND VGND VPWR VPWR _24043_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_7_110_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR _23493_/CLK sky130_fd_sc_hd__clkbuf_1
X_22082_ _21874_/X _22081_/X _14597_/B _22078_/X VGND VGND VPWR VPWR _22082_/X sky130_fd_sc_hd__o22a_4
XFILLER_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21033_ _21033_/A VGND VGND VPWR VPWR _21049_/A sky130_fd_sc_hd__inv_2
XANTENNA__15247__A _13882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13990__A _13990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22984_ _22961_/A _22984_/B VGND VGND VPWR VPWR _22986_/B sky130_fd_sc_hd__nand2_4
XANTENNA__21366__B1 _15155_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21905__A2 _21902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21935_ _21883_/X _21930_/X _14934_/B _21899_/A VGND VGND VPWR VPWR _23574_/D sky130_fd_sc_hd__o22a_4
XFILLER_167_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21866_ _21865_/X _21863_/X _23614_/Q _21858_/X VGND VGND VPWR VPWR _21866_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22808__A _17319_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _24222_/Q _20773_/X _20816_/Y VGND VGND VPWR VPWR _20818_/A sky130_fd_sc_hd__o21a_4
XANTENNA__21712__A _21741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23605_ _23617_/CLK _21886_/X VGND VGND VPWR VPWR _23605_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21669__B2 _21667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19389__A _19377_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21797_ _21587_/X _21791_/X _14470_/B _21795_/X VGND VGND VPWR VPWR _21797_/X sky130_fd_sc_hd__o22a_4
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19731__B1 _17813_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _24438_/Q IRQ[1] VGND VGND VPWR VPWR _11550_/X sky130_fd_sc_hd__and2_4
X_23536_ _23662_/CLK _22001_/X VGND VGND VPWR VPWR _16388_/B sky130_fd_sc_hd__dfxtp_4
X_20748_ _20697_/A VGND VGND VPWR VPWR _20843_/B sky130_fd_sc_hd__buf_2
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23467_ _23467_/CLK _22119_/X VGND VGND VPWR VPWR _23467_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22618__B1 _15473_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20679_ _20679_/A _20494_/B VGND VGND VPWR VPWR _20679_/X sky130_fd_sc_hd__or2_4
XFILLER_149_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14326__A _13655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13220_ _13220_/A _23687_/Q VGND VGND VPWR VPWR _13220_/X sky130_fd_sc_hd__or2_4
XANTENNA__13230__A _13230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18298__B1 _18176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22418_ _20377_/A VGND VGND VPWR VPWR _22418_/X sky130_fd_sc_hd__buf_2
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23398_ _24102_/CLK _22249_/X VGND VGND VPWR VPWR _23398_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22543__A _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13151_ _13338_/A _13151_/B _13150_/X VGND VGND VPWR VPWR _13151_/X sky130_fd_sc_hd__or3_4
X_22349_ _14723_/B VGND VGND VPWR VPWR _23321_/D sky130_fd_sc_hd__buf_2
XANTENNA__16541__A _12001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12102_ _12102_/A _23123_/Q VGND VGND VPWR VPWR _12104_/B sky130_fd_sc_hd__or2_4
XFILLER_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13082_ _13099_/A _13079_/X _13082_/C VGND VGND VPWR VPWR _13082_/X sky130_fd_sc_hd__and3_4
XANTENNA__21159__A _21152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13884__B _13807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24131__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11685__A _11684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24019_ _23889_/CLK _24019_/D VGND VGND VPWR VPWR _24019_/Q sky130_fd_sc_hd__dfxtp_4
X_12033_ _11905_/X VGND VGND VPWR VPWR _16594_/A sky130_fd_sc_hd__buf_2
XFILLER_78_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16910_ _16910_/A VGND VGND VPWR VPWR _16911_/D sky130_fd_sc_hd__inv_2
XANTENNA__15157__A _14272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17890_ _18409_/A VGND VGND VPWR VPWR _17890_/X sky130_fd_sc_hd__buf_2
XANTENNA__14061__A _13696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16841_ _13269_/X _16841_/B VGND VGND VPWR VPWR _16896_/A sky130_fd_sc_hd__or2_4
XFILLER_38_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14996__A _13952_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_15_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_78_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19560_ _19560_/A VGND VGND VPWR VPWR _19849_/B sky130_fd_sc_hd__buf_2
X_16772_ _16759_/A _16772_/B _16772_/C VGND VGND VPWR VPWR _16778_/B sky130_fd_sc_hd__and3_4
XANTENNA__24281__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13984_ _13964_/A _23968_/Q VGND VGND VPWR VPWR _13985_/C sky130_fd_sc_hd__or2_4
XFILLER_92_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18511_ _17435_/Y _18510_/X _17441_/X VGND VGND VPWR VPWR _18511_/Y sky130_fd_sc_hd__o21ai_4
X_15723_ _12783_/X _23748_/Q VGND VGND VPWR VPWR _15724_/C sky130_fd_sc_hd__or2_4
X_12935_ _12942_/A _12935_/B VGND VGND VPWR VPWR _12937_/B sky130_fd_sc_hd__or2_4
X_19491_ _24174_/Q _19455_/Y HRDATA[26] _19452_/X VGND VGND VPWR VPWR _19491_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13405__A _13379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18442_ _18441_/X VGND VGND VPWR VPWR _18442_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15654_ _15582_/X _15652_/Y VGND VGND VPWR VPWR _15654_/X sky130_fd_sc_hd__or2_4
X_12866_ _12866_/A _12861_/X _12866_/C VGND VGND VPWR VPWR _12866_/X sky130_fd_sc_hd__or3_4
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14605_ _12484_/A _14684_/B VGND VGND VPWR VPWR _14605_/X sky130_fd_sc_hd__or2_4
X_18373_ _18032_/X VGND VGND VPWR VPWR _18373_/X sky130_fd_sc_hd__buf_2
X_11817_ _11717_/X _21317_/A VGND VGND VPWR VPWR _11817_/X sky130_fd_sc_hd__or2_4
X_15585_ _14647_/X _15585_/B _15585_/C VGND VGND VPWR VPWR _15585_/X sky130_fd_sc_hd__and3_4
XFILLER_159_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12834_/A _12797_/B VGND VGND VPWR VPWR _12798_/C sky130_fd_sc_hd__or2_4
XANTENNA__16716__A _16595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22321__A2 _22294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17324_ _15382_/B _17324_/B VGND VGND VPWR VPWR _17324_/X sky130_fd_sc_hd__or2_4
XANTENNA__15620__A _15620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _13752_/A _14536_/B _14535_/X VGND VGND VPWR VPWR _14536_/X sky130_fd_sc_hd__and3_4
XFILLER_18_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20332__A1 _20306_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11748_ _12168_/A _11745_/X _11748_/C VGND VGND VPWR VPWR _11749_/C sky130_fd_sc_hd__and3_4
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17255_ _16685_/X VGND VGND VPWR VPWR _17255_/X sky130_fd_sc_hd__buf_2
XFILLER_146_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14467_ _12540_/A _24091_/Q VGND VGND VPWR VPWR _14468_/C sky130_fd_sc_hd__or2_4
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11679_ _15377_/A VGND VGND VPWR VPWR _11680_/A sky130_fd_sc_hd__buf_2
XFILLER_174_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16206_ _16222_/A _16198_/X _16206_/C VGND VGND VPWR VPWR _16207_/C sky130_fd_sc_hd__and3_4
X_13418_ _13342_/Y _13417_/X VGND VGND VPWR VPWR _13582_/A sky130_fd_sc_hd__and2_4
XFILLER_128_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22085__B2 _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17186_ _15116_/X VGND VGND VPWR VPWR _18744_/A sky130_fd_sc_hd__inv_2
XFILLER_31_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14398_ _14383_/A _14396_/X _14398_/C VGND VGND VPWR VPWR _14398_/X sky130_fd_sc_hd__and3_4
XANTENNA__12573__A1 _13453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16137_ _16110_/A _16135_/X _16136_/X VGND VGND VPWR VPWR _16138_/C sky130_fd_sc_hd__and3_4
XANTENNA__17547__A _17274_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13349_ _13349_/A VGND VGND VPWR VPWR _13410_/A sky130_fd_sc_hd__buf_2
XANTENNA__21832__B2 _21822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16068_ _16222_/A _16068_/B _16068_/C VGND VGND VPWR VPWR _16068_/X sky130_fd_sc_hd__and3_4
XFILLER_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11595__A _11595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22388__A2 _22383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15019_ _15000_/A _23605_/Q VGND VGND VPWR VPWR _15019_/X sky130_fd_sc_hd__or2_4
XFILLER_68_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22900__B _22899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17264__A1 _17261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21060__A2 _21059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19827_ _19899_/A _19826_/X VGND VGND VPWR VPWR _19828_/D sky130_fd_sc_hd__nor2_4
XFILLER_69_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19758_ _19696_/X _19756_/Y _20917_/B _19573_/A VGND VGND VPWR VPWR _19758_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18709_ _18709_/A _18709_/B VGND VGND VPWR VPWR _18709_/X sky130_fd_sc_hd__or2_4
X_19689_ _19819_/A _19689_/B VGND VGND VPWR VPWR _19689_/X sky130_fd_sc_hd__and2_4
XFILLER_25_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13315__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21720_ _21727_/A VGND VGND VPWR VPWR _21720_/X sky130_fd_sc_hd__buf_2
XANTENNA__22560__A2 _22558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21651_ _21594_/X _21648_/X _23736_/Q _21645_/X VGND VGND VPWR VPWR _21651_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_35_0_HCLK clkbuf_7_34_0_HCLK/A VGND VGND VPWR VPWR _23119_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_33_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15530__A _12258_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20602_ _20470_/X _20601_/X _24390_/Q _20429_/X VGND VGND VPWR VPWR _20602_/X sky130_fd_sc_hd__o22a_4
X_24370_ _24397_/CLK _18970_/X HRESETn VGND VGND VPWR VPWR _24370_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA_clkbuf_4_9_0_HCLK_A clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_98_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR _23303_/CLK sky130_fd_sc_hd__clkbuf_1
X_21582_ _20841_/A VGND VGND VPWR VPWR _21582_/X sky130_fd_sc_hd__buf_2
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23321_ _23391_/CLK _23321_/D VGND VGND VPWR VPWR _14723_/B sky130_fd_sc_hd__dfxtp_4
X_20533_ _20533_/A VGND VGND VPWR VPWR _20533_/X sky130_fd_sc_hd__buf_2
XFILLER_137_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14146__A _14003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22076__A1 _21865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23252_ _23476_/CLK _22492_/X VGND VGND VPWR VPWR _11845_/B sky130_fd_sc_hd__dfxtp_4
X_20464_ _20464_/A VGND VGND VPWR VPWR _20464_/X sky130_fd_sc_hd__buf_2
XFILLER_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22076__B2 _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24154__CLK _24302_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22203_ _22137_/X _22201_/X _15830_/B _22198_/X VGND VGND VPWR VPWR _22203_/X sky130_fd_sc_hd__o22a_4
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21823__B2 _21822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23183_ _23119_/CLK _22600_/X VGND VGND VPWR VPWR _16273_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16361__A _11784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20395_ _21821_/A VGND VGND VPWR VPWR _20395_/X sky130_fd_sc_hd__buf_2
XFILLER_118_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_HCLK clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22134_ _20658_/A VGND VGND VPWR VPWR _22134_/X sky130_fd_sc_hd__buf_2
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22379__A2 _22376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22065_ _21845_/X _22060_/X _23494_/Q _22064_/X VGND VGND VPWR VPWR _22065_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21016_ _20343_/A _21015_/X _24309_/Q _20352_/A VGND VGND VPWR VPWR _21016_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21051__A2 _21045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21339__B1 _12533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22967_ _18525_/X _22938_/B VGND VGND VPWR VPWR _22967_/X sky130_fd_sc_hd__or2_4
XANTENNA__18755__A1 _17100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13225__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12720_ _12689_/A _12809_/B VGND VGND VPWR VPWR _12720_/X sky130_fd_sc_hd__or2_4
XANTENNA__17920__A _17919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21918_ _21853_/X _21916_/X _15866_/B _21913_/X VGND VGND VPWR VPWR _21918_/X sky130_fd_sc_hd__o22a_4
X_22898_ _19915_/X _22840_/X _15915_/Y _20665_/X VGND VGND VPWR VPWR _22898_/X sky130_fd_sc_hd__o22a_4
XFILLER_167_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12651_ _12651_/A _12548_/B VGND VGND VPWR VPWR _12651_/X sky130_fd_sc_hd__or2_4
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21849_ _21848_/X _21839_/X _23621_/Q _21846_/X VGND VGND VPWR VPWR _23621_/D sky130_fd_sc_hd__o22a_4
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16536__A _12106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22303__A2 _22301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15440__A _13676_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11602_ _17091_/A _11590_/X _11598_/X _17078_/C VGND VGND VPWR VPWR _11635_/A sky130_fd_sc_hd__or4_4
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12582_ _12600_/A VGND VGND VPWR VPWR _12583_/A sky130_fd_sc_hd__buf_2
X_15370_ _13699_/A _23480_/Q VGND VGND VPWR VPWR _15372_/B sky130_fd_sc_hd__or2_4
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ _12191_/A _14406_/B VGND VGND VPWR VPWR _14321_/X sky130_fd_sc_hd__or2_4
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _24359_/Q _19030_/A VGND VGND VPWR VPWR _11533_/X sky130_fd_sc_hd__or2_4
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23519_ _23582_/CLK _22025_/X VGND VGND VPWR VPWR _23519_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17191__B1 _14549_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24499_ _24472_/CLK _17787_/X HRESETn VGND VGND VPWR VPWR _24499_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ _17297_/A _17039_/X VGND VGND VPWR VPWR _17040_/X sky130_fd_sc_hd__and2_4
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14252_ _14240_/A _24095_/Q VGND VGND VPWR VPWR _14252_/X sky130_fd_sc_hd__or2_4
XFILLER_143_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13203_ _13251_/A _13197_/X _13202_/X VGND VGND VPWR VPWR _13211_/B sky130_fd_sc_hd__or3_4
XANTENNA__13895__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14183_ _14226_/A VGND VGND VPWR VPWR _14196_/A sky130_fd_sc_hd__buf_2
XANTENNA__16271__A _16099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17494__A1 _17491_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13134_ _12696_/A _13204_/B VGND VGND VPWR VPWR _13134_/X sky130_fd_sc_hd__or2_4
XFILLER_3_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18991_ _18987_/X _18988_/Y _18989_/Y _18990_/X VGND VGND VPWR VPWR _18991_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17494__B2 _17493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13065_ _13095_/A _23784_/Q VGND VGND VPWR VPWR _13066_/C sky130_fd_sc_hd__or2_4
X_17942_ _17875_/X _17931_/X _17848_/X _17941_/X VGND VGND VPWR VPWR _17943_/A sky130_fd_sc_hd__o22a_4
XFILLER_112_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12016_ _12001_/A _12016_/B _12016_/C VGND VGND VPWR VPWR _12017_/C sky130_fd_sc_hd__and3_4
XANTENNA__21617__A _21617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17873_ _11610_/X VGND VGND VPWR VPWR _17873_/X sky130_fd_sc_hd__buf_2
XFILLER_61_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19612_ _19612_/A VGND VGND VPWR VPWR _19781_/A sky130_fd_sc_hd__buf_2
X_16824_ _16824_/A _16823_/X VGND VGND VPWR VPWR _16824_/X sky130_fd_sc_hd__or2_4
XANTENNA__15615__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20240__B HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19543_ _19480_/X _19542_/X HRDATA[6] _19484_/X VGND VGND VPWR VPWR _19629_/A sky130_fd_sc_hd__o22a_4
X_16755_ _11768_/X VGND VGND VPWR VPWR _16755_/X sky130_fd_sc_hd__buf_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13967_ _13642_/A _23680_/Q VGND VGND VPWR VPWR _13969_/B sky130_fd_sc_hd__or2_4
XANTENNA__18746__A1 _17817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15706_ _12741_/A _15706_/B _15706_/C VGND VGND VPWR VPWR _15707_/C sky130_fd_sc_hd__and3_4
XANTENNA__13135__A _12721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24027__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12918_ _12651_/A _23369_/Q VGND VGND VPWR VPWR _12918_/X sky130_fd_sc_hd__or2_4
X_19474_ _19438_/B VGND VGND VPWR VPWR _19474_/X sky130_fd_sc_hd__buf_2
XFILLER_61_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16686_ _16687_/A _16685_/X VGND VGND VPWR VPWR _16686_/X sky130_fd_sc_hd__and2_4
X_13898_ _14375_/A _13896_/X _13898_/C VGND VGND VPWR VPWR _13898_/X sky130_fd_sc_hd__and3_4
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18425_ _17387_/Y _18424_/B _18176_/X VGND VGND VPWR VPWR _18425_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21352__A _21338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15637_ _13884_/A _23713_/Q VGND VGND VPWR VPWR _15639_/B sky130_fd_sc_hd__or2_4
X_12849_ _12440_/A _12847_/X _12848_/X VGND VGND VPWR VPWR _12849_/X sky130_fd_sc_hd__and3_4
XANTENNA__15350__A _15372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18356_ _18019_/X VGND VGND VPWR VPWR _18356_/X sky130_fd_sc_hd__buf_2
X_15568_ _14431_/A _15566_/X _15568_/C VGND VGND VPWR VPWR _15568_/X sky130_fd_sc_hd__and3_4
XANTENNA__24177__CLK _24184_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17307_ _17272_/X _17308_/B VGND VGND VPWR VPWR _17307_/X sky130_fd_sc_hd__and2_4
X_14519_ _14519_/A _14455_/B VGND VGND VPWR VPWR _14521_/B sky130_fd_sc_hd__or2_4
XFILLER_30_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19757__A HRDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18287_ _17809_/X _18286_/X _17848_/X _17949_/X VGND VGND VPWR VPWR _18287_/X sky130_fd_sc_hd__o22a_4
X_15499_ _12578_/A _15495_/X _15498_/X VGND VGND VPWR VPWR _15499_/X sky130_fd_sc_hd__or3_4
XFILLER_147_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17238_ _17112_/X VGND VGND VPWR VPWR _17823_/A sky130_fd_sc_hd__buf_2
XANTENNA__22058__B2 _22057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17169_ _15517_/X VGND VGND VPWR VPWR _17169_/X sky130_fd_sc_hd__buf_2
XANTENNA__16181__A _13378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20180_ _20180_/A _20179_/Y VGND VGND VPWR VPWR _20180_/X sky130_fd_sc_hd__or2_4
XFILLER_170_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22911__A _22910_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21018__C1 _21017_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12214__A _15439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23870_ _23101_/CLK _21407_/X VGND VGND VPWR VPWR _13769_/B sky130_fd_sc_hd__dfxtp_4
X_22821_ _17397_/Y _22816_/X _22818_/X _22820_/X VGND VGND VPWR VPWR _22822_/B sky130_fd_sc_hd__o22a_4
XANTENNA__13045__A _13045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22752_ _24121_/Q VGND VGND VPWR VPWR _22781_/A sky130_fd_sc_hd__inv_2
XFILLER_164_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22358__A _22358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21703_ _21598_/X _21698_/X _23702_/Q _21667_/A VGND VGND VPWR VPWR _23702_/D sky130_fd_sc_hd__o22a_4
X_22683_ _22480_/X _22679_/X _15162_/B _22648_/A VGND VGND VPWR VPWR _23127_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12884__A _12884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21634_ _21620_/A VGND VGND VPWR VPWR _21634_/X sky130_fd_sc_hd__buf_2
X_24422_ _24422_/CLK _24422_/D HRESETn VGND VGND VPWR VPWR _24422_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22297__B2 _22291_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21565_ _21280_/A VGND VGND VPWR VPWR _21565_/X sky130_fd_sc_hd__buf_2
X_24353_ _24388_/CLK _24353_/D HRESETn VGND VGND VPWR VPWR _19063_/A sky130_fd_sc_hd__dfstp_4
XFILLER_139_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23544__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23304_ _23496_/CLK _22378_/X VGND VGND VPWR VPWR _12999_/B sky130_fd_sc_hd__dfxtp_4
X_20516_ _20344_/A VGND VGND VPWR VPWR _20516_/X sky130_fd_sc_hd__buf_2
XANTENNA__22049__B2 _22043_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24284_ _24292_/CLK _24284_/D HRESETn VGND VGND VPWR VPWR _24284_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21496_ _21489_/A VGND VGND VPWR VPWR _21496_/X sky130_fd_sc_hd__buf_2
XANTENNA__22093__A _22118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16920__B1 _16915_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23235_ _23303_/CLK _23235_/D VGND VGND VPWR VPWR _15836_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20447_ _20447_/A VGND VGND VPWR VPWR _20447_/X sky130_fd_sc_hd__buf_2
XANTENNA__16091__A _15969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14604__A _13596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21272__A2 _21269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23166_ _23229_/CLK _22624_/X VGND VGND VPWR VPWR _13736_/B sky130_fd_sc_hd__dfxtp_4
X_20378_ _21534_/A VGND VGND VPWR VPWR _20378_/X sky130_fd_sc_hd__buf_2
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22117_ _22117_/A VGND VGND VPWR VPWR _22117_/X sky130_fd_sc_hd__buf_2
XFILLER_69_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23097_ _24090_/CLK _22731_/X VGND VGND VPWR VPWR _14827_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_79_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22048_ _21817_/X _22046_/X _23506_/Q _22043_/X VGND VGND VPWR VPWR _23506_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18425__B1 _18176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22221__B2 _22184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11963__A _11963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14870_ _14991_/A _14866_/X _14869_/X VGND VGND VPWR VPWR _14870_/X sky130_fd_sc_hd__or3_4
XFILLER_60_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16451__A2 _11631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13821_ _15412_/A _13821_/B _13820_/X VGND VGND VPWR VPWR _13821_/X sky130_fd_sc_hd__or3_4
XFILLER_91_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23999_ _23997_/CLK _23999_/D VGND VGND VPWR VPWR _23999_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16540_ _16539_/X _23762_/Q VGND VGND VPWR VPWR _16541_/C sky130_fd_sc_hd__or2_4
X_13752_ _13752_/A _13750_/X _13752_/C VGND VGND VPWR VPWR _13756_/B sky130_fd_sc_hd__and3_4
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24198__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12703_ _13279_/A _24010_/Q VGND VGND VPWR VPWR _12703_/X sky130_fd_sc_hd__or2_4
XANTENNA__17400__A1 _17397_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16471_ _11684_/X _16462_/X _16470_/X VGND VGND VPWR VPWR _16471_/X sky130_fd_sc_hd__and3_4
XANTENNA__17400__B2 _17399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12794__A _12833_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13683_ _15447_/A _13766_/B VGND VGND VPWR VPWR _13684_/C sky130_fd_sc_hd__or2_4
XFILLER_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24127__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18210_ _18192_/X _18197_/Y _18205_/X _18208_/X _18209_/Y VGND VGND VPWR VPWR _18210_/X
+ sky130_fd_sc_hd__a32o_4
X_15422_ _12477_/A _23906_/Q VGND VGND VPWR VPWR _15424_/B sky130_fd_sc_hd__or2_4
XANTENNA__15170__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12634_ _12634_/A VGND VGND VPWR VPWR _12635_/A sky130_fd_sc_hd__buf_2
XFILLER_19_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19190_ _19147_/A _19146_/X _19189_/Y VGND VGND VPWR VPWR _24326_/D sky130_fd_sc_hd__o21a_4
XFILLER_169_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22288__B2 _22284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18141_ _17963_/X _18112_/X _18033_/X _18140_/X VGND VGND VPWR VPWR _18141_/X sky130_fd_sc_hd__o22a_4
XFILLER_129_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15353_ _13695_/A _15351_/X _15352_/X VGND VGND VPWR VPWR _15354_/C sky130_fd_sc_hd__and3_4
X_12565_ _12513_/A _12565_/B VGND VGND VPWR VPWR _12566_/C sky130_fd_sc_hd__or2_4
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_81_0_HCLK clkbuf_6_40_0_HCLK/X VGND VGND VPWR VPWR _23991_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ _14304_/A _14376_/B VGND VGND VPWR VPWR _14304_/X sky130_fd_sc_hd__or2_4
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18072_ _18022_/X _18024_/X _18070_/Y _18027_/X _23049_/B VGND VGND VPWR VPWR _18072_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ _11516_/A _11515_/Y VGND VGND VPWR VPWR _11516_/X sky130_fd_sc_hd__and2_4
XFILLER_11_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15284_ _15257_/A _23960_/Q VGND VGND VPWR VPWR _15284_/X sky130_fd_sc_hd__or2_4
X_12496_ _13666_/A VGND VGND VPWR VPWR _12497_/A sky130_fd_sc_hd__buf_2
XFILLER_116_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17023_ _17022_/X VGND VGND VPWR VPWR _17024_/A sky130_fd_sc_hd__buf_2
X_14235_ _14235_/A _23135_/Q VGND VGND VPWR VPWR _14237_/B sky130_fd_sc_hd__or2_4
XFILLER_171_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14514__A _11781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14166_ _14131_/A _23807_/Q VGND VGND VPWR VPWR _14167_/C sky130_fd_sc_hd__or2_4
XANTENNA__22460__B2 _22457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13117_ _13089_/A _24104_/Q VGND VGND VPWR VPWR _13118_/C sky130_fd_sc_hd__or2_4
X_18974_ _18959_/X _18973_/X _18959_/X _24369_/Q VGND VGND VPWR VPWR _24369_/D sky130_fd_sc_hd__a2bb2o_4
X_14097_ _14137_/A _23359_/Q VGND VGND VPWR VPWR _14099_/B sky130_fd_sc_hd__or2_4
XFILLER_98_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13048_ _11856_/A _11629_/A _13017_/X _12264_/X _13047_/X VGND VGND VPWR VPWR _13049_/A
+ sky130_fd_sc_hd__a32o_4
X_17925_ _17813_/X _17921_/Y _17824_/X _17924_/Y VGND VGND VPWR VPWR _17925_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12969__A _12945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11873__A _12857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15345__A _15369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17856_ _17227_/X VGND VGND VPWR VPWR _17856_/X sky130_fd_sc_hd__buf_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16807_ _16611_/A _23889_/Q VGND VGND VPWR VPWR _16807_/X sky130_fd_sc_hd__or2_4
X_17787_ _11642_/X _17786_/X _24499_/Q _11642_/X VGND VGND VPWR VPWR _17787_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14999_ _15022_/A _14995_/X _14999_/C VGND VGND VPWR VPWR _14999_/X sky130_fd_sc_hd__or3_4
XFILLER_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19526_ _19624_/B _19682_/A VGND VGND VPWR VPWR _19550_/B sky130_fd_sc_hd__or2_4
X_16738_ _12064_/X _23665_/Q VGND VGND VPWR VPWR _16738_/X sky130_fd_sc_hd__or2_4
XFILLER_35_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19457_ _19457_/A VGND VGND VPWR VPWR _19457_/X sky130_fd_sc_hd__buf_2
XFILLER_62_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16669_ _16676_/A _23122_/Q VGND VGND VPWR VPWR _16671_/B sky130_fd_sc_hd__or2_4
XANTENNA__16176__A _13398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15080__A _15080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18408_ _18282_/A _17384_/X VGND VGND VPWR VPWR _18408_/X sky130_fd_sc_hd__and2_4
X_19388_ _19381_/X _17012_/X _19381_/X _24243_/Q VGND VGND VPWR VPWR _24243_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21810__A _21809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18339_ _17227_/X _18083_/Y _17833_/A _18085_/X VGND VGND VPWR VPWR _18339_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12209__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21350_ _21283_/X _21348_/X _15819_/B _21345_/X VGND VGND VPWR VPWR _21350_/X sky130_fd_sc_hd__o22a_4
XFILLER_124_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17719__B _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20301_ _20772_/A VGND VGND VPWR VPWR _20533_/A sky130_fd_sc_hd__buf_2
X_21281_ _21269_/A VGND VGND VPWR VPWR _21281_/X sky130_fd_sc_hd__buf_2
XANTENNA__14424__A _13687_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13192__A1 _11857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23020_ _22949_/A _23020_/B VGND VGND VPWR VPWR _23020_/X sky130_fd_sc_hd__or2_4
X_20232_ _24276_/Q _20231_/X VGND VGND VPWR VPWR _20232_/X sky130_fd_sc_hd__or2_4
XFILLER_144_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22451__B2 _22445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22641__A _22648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20163_ _24448_/Q VGND VGND VPWR VPWR _20163_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21257__A _21269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22203__B2 _22198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20094_ _20093_/X VGND VGND VPWR VPWR _20099_/B sky130_fd_sc_hd__inv_2
XANTENNA__17454__B _17481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12879__A _12906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11783__A _13092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23922_ _23922_/CLK _23922_/D VGND VGND VPWR VPWR _23922_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15255__A _14003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23853_ _24045_/CLK _21436_/X VGND VGND VPWR VPWR _16140_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24342__CLK _24342_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22506__A2 _22501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22804_ _22803_/X VGND VGND VPWR VPWR _22804_/X sky130_fd_sc_hd__buf_2
X_23784_ _23561_/CLK _23784_/D VGND VGND VPWR VPWR _23784_/Q sky130_fd_sc_hd__dfxtp_4
X_20996_ _20259_/A _20996_/B VGND VGND VPWR VPWR _20996_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15702__B _15702_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24349__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22735_ _21024_/A _22708_/A _23093_/Q _22698_/A VGND VGND VPWR VPWR _22735_/X sky130_fd_sc_hd__o22a_4
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16086__A _16016_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13503__A _12941_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22666_ _22449_/X _22665_/X _15759_/B _22662_/X VGND VGND VPWR VPWR _23140_/D sky130_fd_sc_hd__o22a_4
XFILLER_139_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21720__A _21727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24405_ _23409_/CLK _18885_/X HRESETn VGND VGND VPWR VPWR _24405_/Q sky130_fd_sc_hd__dfrtp_4
X_21617_ _21617_/A VGND VGND VPWR VPWR _21617_/X sky130_fd_sc_hd__buf_2
X_22597_ _22418_/X _22594_/X _16774_/B _22591_/X VGND VGND VPWR VPWR _23185_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16814__A _16611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21493__A2 _21492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12350_ _12370_/A _12223_/B VGND VGND VPWR VPWR _12350_/X sky130_fd_sc_hd__or2_4
XFILLER_127_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24336_ _24277_/CLK _19170_/X HRESETn VGND VGND VPWR VPWR _24336_/Q sky130_fd_sc_hd__dfrtp_4
X_21548_ _20509_/A VGND VGND VPWR VPWR _21548_/X sky130_fd_sc_hd__buf_2
XFILLER_138_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20336__A _20336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12281_ _13300_/A _12392_/B VGND VGND VPWR VPWR _12281_/X sky130_fd_sc_hd__or2_4
XANTENNA__11958__A _16148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21479_ _21243_/X _21478_/X _23827_/Q _21475_/X VGND VGND VPWR VPWR _23827_/D sky130_fd_sc_hd__o22a_4
X_24267_ _24495_/CLK _19348_/X HRESETn VGND VGND VPWR VPWR _24267_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14020_ _13696_/A _14018_/X _14019_/X VGND VGND VPWR VPWR _14020_/X sky130_fd_sc_hd__and3_4
XFILLER_84_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23218_ _23537_/CLK _22546_/X VGND VGND VPWR VPWR _16621_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_101_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22551__A _22558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24198_ _23511_/CLK _19782_/X HRESETn VGND VGND VPWR VPWR _11663_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_106_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23149_ _24045_/CLK _22653_/X VGND VGND VPWR VPWR _16139_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_161_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14988__B _23349_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15971_ _15971_/A _15971_/B _15970_/X VGND VGND VPWR VPWR _15971_/X sky130_fd_sc_hd__or3_4
XFILLER_1_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17364__B _17445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12789__A _12800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17710_ _17710_/A _17710_/B VGND VGND VPWR VPWR _17768_/B sky130_fd_sc_hd__or2_4
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15165__A _14574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14922_ _14922_/A _23190_/Q VGND VGND VPWR VPWR _14922_/X sky130_fd_sc_hd__or2_4
X_18690_ _18288_/A _17950_/X VGND VGND VPWR VPWR _18690_/Y sky130_fd_sc_hd__nor2_4
XFILLER_152_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17641_ _17641_/A _18035_/B _17641_/C _17640_/X VGND VGND VPWR VPWR _17642_/C sky130_fd_sc_hd__or4_4
X_14853_ _12218_/A _23734_/Q VGND VGND VPWR VPWR _14854_/C sky130_fd_sc_hd__or2_4
XFILLER_64_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ _12485_/A _23741_/Q VGND VGND VPWR VPWR _13805_/C sky130_fd_sc_hd__or2_4
X_17572_ _17569_/X _17572_/B VGND VGND VPWR VPWR _17572_/X sky130_fd_sc_hd__or2_4
XFILLER_112_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14784_ _14783_/X VGND VGND VPWR VPWR _15091_/A sky130_fd_sc_hd__buf_2
X_11996_ _12102_/A _11827_/B VGND VGND VPWR VPWR _11996_/X sky130_fd_sc_hd__or2_4
X_19311_ _19230_/X VGND VGND VPWR VPWR _19311_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16523_ _16452_/Y _16523_/B VGND VGND VPWR VPWR _16526_/A sky130_fd_sc_hd__and2_4
X_13735_ _15457_/A VGND VGND VPWR VPWR _13744_/A sky130_fd_sc_hd__buf_2
XFILLER_45_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21181__B2 _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13413__A _13413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19242_ _19242_/A _19289_/A VGND VGND VPWR VPWR _19243_/B sky130_fd_sc_hd__and2_4
X_16454_ _16454_/A _16388_/B VGND VGND VPWR VPWR _16455_/C sky130_fd_sc_hd__or2_4
X_13666_ _13666_/A VGND VGND VPWR VPWR _15406_/A sky130_fd_sc_hd__buf_2
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22726__A _22705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15405_ _15405_/A _15401_/X _15405_/C VGND VGND VPWR VPWR _15405_/X sky130_fd_sc_hd__or3_4
X_12617_ _13063_/A VGND VGND VPWR VPWR _12976_/A sky130_fd_sc_hd__buf_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19173_ _19156_/B VGND VGND VPWR VPWR _19173_/Y sky130_fd_sc_hd__inv_2
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16385_ _16384_/X VGND VGND VPWR VPWR _16385_/Y sky130_fd_sc_hd__inv_2
X_13597_ _14311_/A _13702_/B VGND VGND VPWR VPWR _13597_/X sky130_fd_sc_hd__or2_4
XFILLER_12_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12029__A _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18124_ _17988_/X _17923_/X _17933_/X _17927_/X VGND VGND VPWR VPWR _18125_/B sky130_fd_sc_hd__a22oi_4
X_15336_ _13704_/A _23448_/Q VGND VGND VPWR VPWR _15337_/C sky130_fd_sc_hd__or2_4
X_12548_ _12894_/A _12548_/B VGND VGND VPWR VPWR _12548_/X sky130_fd_sc_hd__or2_4
XANTENNA__21484__A2 _21478_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18885__B1 _24405_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22681__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18055_ _18320_/A _18054_/Y VGND VGND VPWR VPWR _18055_/X sky130_fd_sc_hd__and2_4
XANTENNA__11868__A _11867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15267_ _15267_/A _23672_/Q VGND VGND VPWR VPWR _15267_/X sky130_fd_sc_hd__or2_4
X_12479_ _12878_/A VGND VGND VPWR VPWR _12867_/A sky130_fd_sc_hd__buf_2
XFILLER_145_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24215__CLK _24248_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17006_ _17006_/A _16976_/X _17005_/X _16973_/X VGND VGND VPWR VPWR _17906_/C sky130_fd_sc_hd__or4_4
X_14218_ _14254_/A _14117_/B VGND VGND VPWR VPWR _14218_/X sky130_fd_sc_hd__or2_4
XANTENNA__15059__B _15059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15198_ _14226_/A VGND VGND VPWR VPWR _15198_/X sky130_fd_sc_hd__buf_2
XANTENNA__22461__A _22461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14149_ _14149_/A _14149_/B _14148_/X VGND VGND VPWR VPWR _14149_/X sky130_fd_sc_hd__and3_4
XFILLER_112_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18957_ _19009_/A VGND VGND VPWR VPWR _18957_/X sky130_fd_sc_hd__buf_2
XANTENNA__12699__A _11935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17908_ _17908_/A _17908_/B VGND VGND VPWR VPWR _17909_/A sky130_fd_sc_hd__and2_4
XANTENNA__20747__A1 _20635_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20747__B2 _20746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18888_ _11609_/X _18888_/B _17113_/X _18887_/X VGND VGND VPWR VPWR _18888_/X sky130_fd_sc_hd__or4_4
XFILLER_67_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17839_ _17837_/X _17166_/X _17838_/X _17171_/X VGND VGND VPWR VPWR _17839_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17290__A _14700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15803__A _12863_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20850_ _20644_/X _20849_/X _24284_/Q _20758_/X VGND VGND VPWR VPWR _20850_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19509_ _19680_/A _19546_/A _19675_/A VGND VGND VPWR VPWR _19509_/X sky130_fd_sc_hd__o21a_4
XFILLER_35_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20781_ _20287_/A VGND VGND VPWR VPWR _20781_/X sky130_fd_sc_hd__buf_2
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21172__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13323__A _12866_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22520_ _22456_/X _22515_/X _15569_/B _22519_/X VGND VGND VPWR VPWR _23233_/D sky130_fd_sc_hd__o22a_4
XFILLER_168_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14138__B _23967_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18833__B _12097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22451_ _22449_/X _22450_/X _15657_/B _22445_/X VGND VGND VPWR VPWR _23268_/D sky130_fd_sc_hd__o22a_4
XFILLER_10_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21402_ _21388_/A VGND VGND VPWR VPWR _21402_/X sky130_fd_sc_hd__buf_2
X_22382_ _22132_/X _22376_/X _23301_/Q _22380_/X VGND VGND VPWR VPWR _22382_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13977__B _23168_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21333_ _21254_/X _21327_/X _16279_/B _21331_/X VGND VGND VPWR VPWR _23919_/D sky130_fd_sc_hd__o22a_4
X_24121_ _23544_/CLK _22783_/X HRESETn VGND VGND VPWR VPWR _24121_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21264_ _21264_/A VGND VGND VPWR VPWR _21264_/X sky130_fd_sc_hd__buf_2
X_24052_ _23668_/CLK _21088_/X VGND VGND VPWR VPWR _21080_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21227__A2 _21226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22424__B2 _22421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23003_ _18350_/X _23003_/B VGND VGND VPWR VPWR _23004_/C sky130_fd_sc_hd__or2_4
X_20215_ _20214_/X VGND VGND VPWR VPWR _20218_/B sky130_fd_sc_hd__inv_2
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21195_ _21195_/A VGND VGND VPWR VPWR _21195_/X sky130_fd_sc_hd__buf_2
XFILLER_131_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20146_ _20146_/A _20145_/Y VGND VGND VPWR VPWR _20147_/B sky130_fd_sc_hd__or2_4
XANTENNA__22727__A2 _22722_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20077_ _20064_/X _18500_/A _20070_/X _20076_/X VGND VGND VPWR VPWR _20077_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12402__A _12950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20738__A1 _18494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24472__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23905_ _23744_/CLK _23905_/D VGND VGND VPWR VPWR _15552_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15713__A _12851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ _16684_/A _11831_/X _11850_/C VGND VGND VPWR VPWR _11850_/X sky130_fd_sc_hd__or3_4
X_23836_ _23515_/CLK _23836_/D VGND VGND VPWR VPWR _14388_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _11781_/A VGND VGND VPWR VPWR _12354_/A sky130_fd_sc_hd__buf_2
XANTENNA__17367__B1 _17358_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23767_ _23770_/CLK _21597_/X VGND VGND VPWR VPWR _15130_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21163__B2 _21159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14329__A _14329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20979_ _22480_/A VGND VGND VPWR VPWR _21311_/A sky130_fd_sc_hd__buf_2
XFILLER_53_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _13520_/A _13514_/X _13520_/C VGND VGND VPWR VPWR _13529_/B sky130_fd_sc_hd__or3_4
X_22718_ _21570_/A _22715_/X _15501_/B _22712_/X VGND VGND VPWR VPWR _23106_/D sky130_fd_sc_hd__o22a_4
XFILLER_25_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23698_ _23852_/CLK _23698_/D VGND VGND VPWR VPWR _23698_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13451_ _12869_/A _13451_/B _13451_/C VGND VGND VPWR VPWR _13452_/C sky130_fd_sc_hd__and3_4
X_22649_ _22420_/X _22644_/X _16428_/B _22648_/X VGND VGND VPWR VPWR _23152_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16544__A _12106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12402_ _12950_/A VGND VGND VPWR VPWR _12402_/X sky130_fd_sc_hd__buf_2
XFILLER_142_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16170_ _13408_/A VGND VGND VPWR VPWR _16215_/A sky130_fd_sc_hd__buf_2
XANTENNA__21466__A2 _21462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13382_ _13400_/A _13373_/X _13382_/C VGND VGND VPWR VPWR _13383_/C sky130_fd_sc_hd__and3_4
XANTENNA__22663__B2 _22662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20066__A _19950_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11688__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15121_ _14911_/X _17339_/A _15120_/Y VGND VGND VPWR VPWR _15121_/X sky130_fd_sc_hd__o21a_4
X_12333_ _11701_/A _12333_/B _12332_/X VGND VGND VPWR VPWR _12343_/B sky130_fd_sc_hd__and3_4
X_24319_ _24287_/CLK _24319_/D HRESETn VGND VGND VPWR VPWR _24319_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14064__A _11736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21218__A2 _21212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15052_ _15078_/A _15050_/X _15052_/C VGND VGND VPWR VPWR _15058_/B sky130_fd_sc_hd__and3_4
X_12264_ _11606_/A VGND VGND VPWR VPWR _12264_/X sky130_fd_sc_hd__buf_2
XANTENNA__20216__D _20216_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22415__B2 _22409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24388__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14999__A _15022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14003_ _14003_/A _14003_/B _14003_/C VGND VGND VPWR VPWR _14004_/C sky130_fd_sc_hd__and3_4
X_19860_ _19678_/B _19744_/X _19675_/A VGND VGND VPWR VPWR _19895_/C sky130_fd_sc_hd__o21a_4
X_12195_ _12501_/A VGND VGND VPWR VPWR _13630_/A sky130_fd_sc_hd__buf_2
X_18811_ _18789_/A VGND VGND VPWR VPWR _18811_/X sky130_fd_sc_hd__buf_2
X_19791_ HRDATA[0] VGND VGND VPWR VPWR _19791_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22718__A2 _22715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13408__A _13408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15954_ _16006_/A VGND VGND VPWR VPWR _15961_/A sky130_fd_sc_hd__buf_2
X_18742_ _18499_/X _18740_/X _18527_/X _18741_/X VGND VGND VPWR VPWR _18742_/X sky130_fd_sc_hd__o22a_4
XFILLER_48_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14905_ _14905_/A _23702_/Q VGND VGND VPWR VPWR _14907_/B sky130_fd_sc_hd__or2_4
X_18673_ _17101_/A _18673_/B VGND VGND VPWR VPWR _18674_/C sky130_fd_sc_hd__or2_4
X_15885_ _13496_/A _15823_/B VGND VGND VPWR VPWR _15885_/X sky130_fd_sc_hd__or2_4
XANTENNA__24142__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17624_ _17341_/A VGND VGND VPWR VPWR _17624_/Y sky130_fd_sc_hd__inv_2
X_14836_ _14693_/A _14836_/B _14835_/X VGND VGND VPWR VPWR _14840_/B sky130_fd_sc_hd__and3_4
XFILLER_56_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17555_ _17641_/A VGND VGND VPWR VPWR _17583_/A sky130_fd_sc_hd__inv_2
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14767_ _14766_/X VGND VGND VPWR VPWR _14767_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22642__A2_N _22641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11979_ _12012_/A _11795_/B VGND VGND VPWR VPWR _11979_/X sky130_fd_sc_hd__or2_4
XANTENNA__21154__B2 _21152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16506_ _16481_/X _16443_/B VGND VGND VPWR VPWR _16507_/C sky130_fd_sc_hd__or2_4
X_13718_ _15372_/A VGND VGND VPWR VPWR _13719_/A sky130_fd_sc_hd__buf_2
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17486_ _17485_/X VGND VGND VPWR VPWR _17486_/Y sky130_fd_sc_hd__inv_2
X_14698_ _13894_/A _14698_/B _14697_/X VGND VGND VPWR VPWR _14699_/C sky130_fd_sc_hd__and3_4
XFILLER_60_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22456__A _20744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16437_ _16094_/A _16435_/X _16436_/X VGND VGND VPWR VPWR _16441_/B sky130_fd_sc_hd__and3_4
X_19225_ _22945_/A _24309_/Q _19224_/Y VGND VGND VPWR VPWR _24309_/D sky130_fd_sc_hd__o21a_4
XANTENNA__24395__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13649_ _12288_/A _13649_/B _13648_/X VGND VGND VPWR VPWR _13649_/X sky130_fd_sc_hd__or3_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19156_ _19156_/A _19156_/B VGND VGND VPWR VPWR _19157_/B sky130_fd_sc_hd__and2_4
X_16368_ _16465_/A _16366_/X _16367_/X VGND VGND VPWR VPWR _16369_/C sky130_fd_sc_hd__and3_4
XANTENNA__21457__A2 _21455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22654__B2 _22648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_51_0_HCLK clkbuf_6_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18107_ _18107_/A VGND VGND VPWR VPWR _18111_/C sky130_fd_sc_hd__inv_2
X_15319_ _15319_/A _23736_/Q VGND VGND VPWR VPWR _15320_/C sky130_fd_sc_hd__or2_4
X_19087_ _11523_/A VGND VGND VPWR VPWR _19087_/Y sky130_fd_sc_hd__inv_2
X_16299_ _16003_/A _16295_/X _16298_/X VGND VGND VPWR VPWR _16299_/X sky130_fd_sc_hd__or3_4
XANTENNA__22903__B _22902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18038_ _18037_/X _17561_/B VGND VGND VPWR VPWR _18038_/Y sky130_fd_sc_hd__nor2_4
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22191__A _22176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17285__A _11611_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14702__A _14613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20000_ _18017_/X _19983_/X _19999_/Y _19994_/X VGND VGND VPWR VPWR _20000_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20968__B2 _20282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19989_ _17897_/X _19983_/X _19988_/Y _19979_/X VGND VGND VPWR VPWR _19989_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22709__A2 _22708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13318__A _13318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21951_ _21821_/X _21946_/X _16409_/B _21950_/X VGND VGND VPWR VPWR _23568_/D sky130_fd_sc_hd__o22a_4
XFILLER_28_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21393__B2 _21388_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16629__A _16682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20902_ _20899_/X _20901_/X _20262_/X VGND VGND VPWR VPWR _20902_/Y sky130_fd_sc_hd__o21ai_4
X_21882_ _21881_/X _21875_/X _15222_/B _21809_/X VGND VGND VPWR VPWR _23607_/D sky130_fd_sc_hd__o22a_4
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _23557_/CLK _23621_/D VGND VGND VPWR VPWR _23621_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833_ _20930_/A _20832_/X VGND VGND VPWR VPWR _20833_/Y sky130_fd_sc_hd__nor2_4
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21696__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22893__A1 _17261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23552_ _24096_/CLK _21973_/X VGND VGND VPWR VPWR _23552_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20764_ _18525_/X _20702_/X _20753_/X _20763_/Y VGND VGND VPWR VPWR _20764_/X sky130_fd_sc_hd__a211o_4
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22366__A _22366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22503_ _22428_/X _22501_/X _16149_/B _22498_/X VGND VGND VPWR VPWR _22503_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12892__A _12864_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23483_ _23323_/CLK _22080_/X VGND VGND VPWR VPWR _23483_/Q sky130_fd_sc_hd__dfxtp_4
X_20695_ _20231_/A VGND VGND VPWR VPWR _20695_/X sky130_fd_sc_hd__buf_2
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22434_ _22432_/X _22426_/X _12579_/B _22433_/X VGND VGND VPWR VPWR _22434_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22645__B2 _22641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23285__CLK _23392_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22365_ _22103_/X _22362_/X _16766_/B _22359_/X VGND VGND VPWR VPWR _22365_/X sky130_fd_sc_hd__o22a_4
XFILLER_163_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24104_ _23337_/CLK _24104_/D VGND VGND VPWR VPWR _24104_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_163_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21316_ _21315_/X _21269_/A _23925_/Q _21239_/X VGND VGND VPWR VPWR _23925_/D sky130_fd_sc_hd__o22a_4
XFILLER_151_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22296_ _22125_/X _22294_/X _12991_/B _22291_/X VGND VGND VPWR VPWR _23368_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20614__A _20510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24035_ _23939_/CLK _21113_/X VGND VGND VPWR VPWR _15799_/B sky130_fd_sc_hd__dfxtp_4
X_21247_ _21532_/A VGND VGND VPWR VPWR _21247_/X sky130_fd_sc_hd__buf_2
XFILLER_117_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21178_ _20938_/X _21176_/X _14721_/B _21173_/X VGND VGND VPWR VPWR _23993_/D sky130_fd_sc_hd__o22a_4
XFILLER_77_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13228__A _12354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20129_ _11640_/B _20128_/X _11639_/A _18685_/Y VGND VGND VPWR VPWR _20129_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19577__A1 _20364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21445__A _21438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12951_ _12951_/A _23625_/Q VGND VGND VPWR VPWR _12953_/B sky130_fd_sc_hd__or2_4
XFILLER_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20187__A2 IRQ[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16539__A _12015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11971__A _13453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11902_ _11902_/A VGND VGND VPWR VPWR _13427_/A sky130_fd_sc_hd__buf_2
XANTENNA__15443__A _12190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15670_ _12726_/A _15666_/X _15669_/X VGND VGND VPWR VPWR _15670_/X sky130_fd_sc_hd__or3_4
XFILLER_93_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12882_ _12882_/A _12882_/B VGND VGND VPWR VPWR _12882_/X sky130_fd_sc_hd__and2_4
XFILLER_34_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19329__A1 _17037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14621_ _14676_/A _14621_/B _14621_/C VGND VGND VPWR VPWR _14621_/X sky130_fd_sc_hd__and3_4
X_23819_ _24074_/CLK _21490_/X VGND VGND VPWR VPWR _12565_/B sky130_fd_sc_hd__dfxtp_4
X_11833_ _11833_/A _23828_/Q VGND VGND VPWR VPWR _11833_/X sky130_fd_sc_hd__or2_4
XANTENNA__15162__B _15162_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14059__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24060__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17340_ _15118_/X _17340_/B VGND VGND VPWR VPWR _17341_/B sky130_fd_sc_hd__or2_4
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14552_ _14552_/A VGND VGND VPWR VPWR _14552_/Y sky130_fd_sc_hd__inv_2
XPHY_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21687__A2 _21684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11764_ _12156_/A _23796_/Q VGND VGND VPWR VPWR _11765_/C sky130_fd_sc_hd__or2_4
XPHY_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22276__A _22291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _12941_/A VGND VGND VPWR VPWR _13503_/X sky130_fd_sc_hd__buf_2
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17271_ _17911_/B VGND VGND VPWR VPWR _17271_/Y sky130_fd_sc_hd__inv_2
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _14482_/X VGND VGND VPWR VPWR _14483_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16274__A _16099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11695_ _11653_/A VGND VGND VPWR VPWR _13694_/A sky130_fd_sc_hd__buf_2
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19010_ _19024_/A VGND VGND VPWR VPWR _19010_/X sky130_fd_sc_hd__buf_2
X_16222_ _16222_/A _16222_/B _16222_/C VGND VGND VPWR VPWR _16238_/B sky130_fd_sc_hd__and3_4
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21439__A2 _21434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13434_ _13475_/A _13428_/X _13434_/C VGND VGND VPWR VPWR _13434_/X sky130_fd_sc_hd__or3_4
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16153_ _16156_/A _23117_/Q VGND VGND VPWR VPWR _16153_/X sky130_fd_sc_hd__or2_4
XFILLER_166_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13365_ _13375_/A _13365_/B VGND VGND VPWR VPWR _13366_/C sky130_fd_sc_hd__or2_4
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12307__A _12741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15104_ _15080_/A _15104_/B VGND VGND VPWR VPWR _15105_/C sky130_fd_sc_hd__or2_4
XFILLER_155_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12316_ _13045_/A _12312_/X _12316_/C VGND VGND VPWR VPWR _12316_/X sky130_fd_sc_hd__or3_4
X_16084_ _11815_/X _16068_/X _16083_/X VGND VGND VPWR VPWR _16085_/C sky130_fd_sc_hd__or3_4
XFILLER_142_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13296_ _13319_/A _13296_/B VGND VGND VPWR VPWR _13296_/X sky130_fd_sc_hd__or2_4
XFILLER_138_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19912_ _20241_/A VGND VGND VPWR VPWR _19913_/A sky130_fd_sc_hd__inv_2
X_15035_ _11877_/A _15033_/X _15035_/C VGND VGND VPWR VPWR _15036_/C sky130_fd_sc_hd__and3_4
X_12247_ _12708_/A _12247_/B _12247_/C VGND VGND VPWR VPWR _12247_/X sky130_fd_sc_hd__or3_4
XANTENNA__15618__A _11675_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19843_ _19849_/A _19839_/X _19842_/Y VGND VGND VPWR VPWR _19843_/X sky130_fd_sc_hd__o21a_4
X_12178_ _16684_/A _12178_/B _12178_/C VGND VGND VPWR VPWR _12178_/X sky130_fd_sc_hd__or3_4
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13138__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24323__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19774_ _19474_/X HRDATA[2] VGND VGND VPWR VPWR _19774_/X sky130_fd_sc_hd__and2_4
XFILLER_96_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16986_ _16986_/A _16985_/X VGND VGND VPWR VPWR _16986_/X sky130_fd_sc_hd__or2_4
XANTENNA__19568__A1 _20339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19568__B2 HRDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18725_ _16933_/Y _18720_/Y _16932_/X _18724_/X VGND VGND VPWR VPWR _20155_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21355__A _21322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15937_ _11889_/X VGND VGND VPWR VPWR _15944_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12977__A _12977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16449__A _11865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21375__B2 _21374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11881__A _11881_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15353__A _13695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15868_ _13543_/X _15868_/B VGND VGND VPWR VPWR _15868_/X sky130_fd_sc_hd__or2_4
X_18656_ _18565_/A _18651_/B _18652_/X _18655_/Y VGND VGND VPWR VPWR _18656_/X sky130_fd_sc_hd__a211o_4
XFILLER_149_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24403__CLK _23409_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17607_ _17391_/X _17606_/X _17385_/X _17393_/X VGND VGND VPWR VPWR _17607_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15072__B _23445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14819_ _14819_/A _14743_/B VGND VGND VPWR VPWR _14821_/B sky130_fd_sc_hd__or2_4
X_15799_ _12847_/A _15799_/B VGND VGND VPWR VPWR _15799_/X sky130_fd_sc_hd__or2_4
X_18587_ _18545_/A _18587_/B VGND VGND VPWR VPWR _18587_/X sky130_fd_sc_hd__and2_4
XANTENNA__21127__B2 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21678__A2 _21677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17538_ _12980_/X _17460_/B VGND VGND VPWR VPWR _17538_/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21090__A _21104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17469_ _17469_/A _17468_/Y VGND VGND VPWR VPWR _18165_/B sky130_fd_sc_hd__or2_4
XFILLER_149_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19208_ _24317_/Q _19138_/B _19207_/Y VGND VGND VPWR VPWR _24317_/D sky130_fd_sc_hd__o21a_4
XANTENNA__13601__A _13601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20480_ _24268_/Q VGND VGND VPWR VPWR _20480_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22627__B2 _22626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19139_ _24318_/Q _19138_/X VGND VGND VPWR VPWR _19205_/A sky130_fd_sc_hd__and2_4
XANTENNA__16912__A _16911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22150_ _22149_/X _22147_/X _13738_/B _22142_/X VGND VGND VPWR VPWR _23454_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17727__B _17399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21101_ _21101_/A VGND VGND VPWR VPWR _21101_/X sky130_fd_sc_hd__buf_2
XANTENNA__15528__A _12186_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22081_ _22041_/A VGND VGND VPWR VPWR _22081_/X sky130_fd_sc_hd__buf_2
XANTENNA__14432__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21032_ _21031_/X VGND VGND VPWR VPWR _21033_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_58_0_HCLK clkbuf_7_59_0_HCLK/A VGND VGND VPWR VPWR _24045_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__13990__B _23136_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12887__A _12867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22983_ _22982_/X VGND VGND VPWR VPWR HADDR[13] sky130_fd_sc_hd__inv_2
XFILLER_41_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21366__B2 _21331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21934_ _21881_/X _21930_/X _15147_/B _21899_/A VGND VGND VPWR VPWR _21934_/X sky130_fd_sc_hd__o22a_4
XFILLER_167_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21865_ _20819_/A VGND VGND VPWR VPWR _21865_/X sky130_fd_sc_hd__buf_2
XANTENNA__18574__A _18399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _23668_/CLK _23604_/D VGND VGND VPWR VPWR _23604_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21669__A2 _21663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ _20857_/A _20815_/X VGND VGND VPWR VPWR _20816_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22866__A1 _17284_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21796_ _21584_/X _21791_/X _23644_/Q _21795_/X VGND VGND VPWR VPWR _21796_/X sky130_fd_sc_hd__o22a_4
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23535_ _23246_/CLK _22002_/X VGND VGND VPWR VPWR _16248_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20747_ _20635_/X _20745_/X _24097_/Q _20746_/X VGND VGND VPWR VPWR _20747_/X sky130_fd_sc_hd__o22a_4
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14607__A _13652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13511__A _12950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23466_ _23404_/CLK _23466_/D VGND VGND VPWR VPWR _12797_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22618__B2 _22612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20678_ _24451_/Q VGND VGND VPWR VPWR _20679_/A sky130_fd_sc_hd__inv_2
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22417_ _22416_/X _22414_/X _16609_/B _22409_/X VGND VGND VPWR VPWR _23282_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19495__B1 HRDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17918__A _17109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23397_ _23397_/CLK _23397_/D VGND VGND VPWR VPWR _23397_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13150_ _12738_/A _13148_/X _13150_/C VGND VGND VPWR VPWR _13150_/X sky130_fd_sc_hd__and3_4
X_22348_ _14570_/B VGND VGND VPWR VPWR _23322_/D sky130_fd_sc_hd__buf_2
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12101_ _12078_/X _12101_/B _12100_/X VGND VGND VPWR VPWR _12101_/X sky130_fd_sc_hd__or3_4
XANTENNA__11966__A _13981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13081_ _13089_/A _13013_/B VGND VGND VPWR VPWR _13082_/C sky130_fd_sc_hd__or2_4
X_22279_ _22275_/A VGND VGND VPWR VPWR _22294_/A sky130_fd_sc_hd__buf_2
XANTENNA__14342__A _13916_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24018_ _23404_/CLK _24018_/D VGND VGND VPWR VPWR _24018_/Q sky130_fd_sc_hd__dfxtp_4
X_12032_ _16700_/A _12114_/B VGND VGND VPWR VPWR _12036_/B sky130_fd_sc_hd__or2_4
XFILLER_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16840_ _13271_/X _16839_/X _13264_/X VGND VGND VPWR VPWR _16841_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__14996__B _24021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16771_ _16757_/X _23601_/Q VGND VGND VPWR VPWR _16772_/C sky130_fd_sc_hd__or2_4
XFILLER_24_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13983_ _13983_/A _14052_/B VGND VGND VPWR VPWR _13983_/X sky130_fd_sc_hd__or2_4
XANTENNA__16269__A _15971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12797__A _12834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21357__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15722_ _12780_/X _15660_/B VGND VGND VPWR VPWR _15722_/X sky130_fd_sc_hd__or2_4
XANTENNA__15173__A _12484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18510_ _17436_/B _18509_/X _17439_/X VGND VGND VPWR VPWR _18510_/X sky130_fd_sc_hd__o21a_4
X_12934_ _12972_/A _12932_/X _12933_/X VGND VGND VPWR VPWR _12938_/B sky130_fd_sc_hd__and3_4
XFILLER_20_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19490_ _19525_/A _19545_/A VGND VGND VPWR VPWR _19494_/A sky130_fd_sc_hd__or2_4
XANTENNA__17091__C _17077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18441_ _18314_/A _18438_/Y _18439_/Y _18440_/X VGND VGND VPWR VPWR _18441_/X sky130_fd_sc_hd__or4_4
X_15653_ _15652_/Y VGND VGND VPWR VPWR _15653_/X sky130_fd_sc_hd__buf_2
XANTENNA__13405__B _13405_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12865_ _12889_/A _12865_/B _12865_/C VGND VGND VPWR VPWR _12866_/C sky130_fd_sc_hd__and3_4
XANTENNA__21109__B2 _21108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14604_ _13596_/A _14604_/B VGND VGND VPWR VPWR _14604_/X sky130_fd_sc_hd__or2_4
XANTENNA__15901__A _13547_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18372_ _17906_/A _18370_/X _24147_/Q _18371_/Y VGND VGND VPWR VPWR _18372_/X sky130_fd_sc_hd__o22a_4
X_11816_ _11815_/X VGND VGND VPWR VPWR _16684_/A sky130_fd_sc_hd__buf_2
XFILLER_159_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22857__A1 _17327_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15584_ _15620_/A _15523_/B VGND VGND VPWR VPWR _15585_/C sky130_fd_sc_hd__or2_4
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _15778_/A VGND VGND VPWR VPWR _12834_/A sky130_fd_sc_hd__buf_2
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17324_/B VGND VGND VPWR VPWR _17323_/Y sky130_fd_sc_hd__inv_2
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _13751_/A _14477_/B VGND VGND VPWR VPWR _14535_/X sky130_fd_sc_hd__or2_4
XFILLER_57_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11746_/X _23764_/Q VGND VGND VPWR VPWR _11748_/C sky130_fd_sc_hd__or2_4
XANTENNA__20332__A2 _20309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13421__A _13330_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20238__B _20844_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22609__A1 _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17254_ _17253_/X VGND VGND VPWR VPWR _17256_/B sky130_fd_sc_hd__inv_2
XFILLER_159_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22609__B2 _22605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14466_ _12498_/A _23483_/Q VGND VGND VPWR VPWR _14466_/X sky130_fd_sc_hd__or2_4
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _13383_/A VGND VGND VPWR VPWR _16053_/A sky130_fd_sc_hd__buf_2
X_16205_ _16205_/A _16205_/B _16205_/C VGND VGND VPWR VPWR _16206_/C sky130_fd_sc_hd__or3_4
XFILLER_146_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13417_ _13417_/A _13417_/B _13417_/C VGND VGND VPWR VPWR _13417_/X sky130_fd_sc_hd__and3_4
XFILLER_174_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22085__A2 _22081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17185_ _17130_/X _17183_/X _17124_/X _17184_/X VGND VGND VPWR VPWR _17185_/X sky130_fd_sc_hd__o22a_4
X_14397_ _14367_/A _14397_/B VGND VGND VPWR VPWR _14398_/C sky130_fd_sc_hd__or2_4
XANTENNA__12037__A _16713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16136_ _16109_/A _24077_/Q VGND VGND VPWR VPWR _16136_/X sky130_fd_sc_hd__or2_4
XFILLER_6_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13348_ _13376_/A _13345_/X _13347_/X VGND VGND VPWR VPWR _13348_/X sky130_fd_sc_hd__and3_4
XFILLER_115_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21832__A2 _21827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11876__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16067_ _11693_/X _16063_/X _16067_/C VGND VGND VPWR VPWR _16068_/C sky130_fd_sc_hd__or3_4
X_13279_ _13279_/A VGND VGND VPWR VPWR _13313_/A sky130_fd_sc_hd__buf_2
XFILLER_170_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15018_ _15018_/A _15016_/X _15017_/X VGND VGND VPWR VPWR _15018_/X sky130_fd_sc_hd__and3_4
XANTENNA__15067__B _23925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20399__A2 _20776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19826_ _19809_/A _19824_/X _19826_/C VGND VGND VPWR VPWR _19826_/X sky130_fd_sc_hd__and3_4
XANTENNA__17563__A _16383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21085__A _21118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19757_ HRDATA[20] VGND VGND VPWR VPWR _20917_/B sky130_fd_sc_hd__buf_2
X_16969_ _24136_/Q VGND VGND VPWR VPWR _17740_/A sky130_fd_sc_hd__inv_2
XANTENNA__15083__A _14682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18708_ _17974_/X _17627_/X _17919_/X _17347_/X VGND VGND VPWR VPWR _18709_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__12500__A _12871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19688_ _19797_/A _19679_/X _19685_/Y _19687_/X VGND VGND VPWR VPWR _19689_/B sky130_fd_sc_hd__a211o_4
XANTENNA__21813__A _21528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18639_ _18518_/A _17632_/A _17797_/A VGND VGND VPWR VPWR _18639_/X sky130_fd_sc_hd__a21o_4
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20571__A2 _20562_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15811__A _12854_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21650_ _21592_/X _21648_/X _14780_/B _21645_/X VGND VGND VPWR VPWR _23737_/D sky130_fd_sc_hd__o22a_4
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20601_ _24422_/Q _20427_/X _20157_/A _20471_/X VGND VGND VPWR VPWR _20601_/X sky130_fd_sc_hd__o22a_4
X_21581_ _21580_/X _21578_/X _13722_/B _21573_/X VGND VGND VPWR VPWR _21581_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14427__A _14431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20148__B _20147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13331__A _13475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23320_ _23416_/CLK _23320_/D VGND VGND VPWR VPWR _22350_/A sky130_fd_sc_hd__dfxtp_4
X_20532_ _20418_/X _20531_/X _24106_/Q _20510_/X VGND VGND VPWR VPWR _24106_/D sky130_fd_sc_hd__o22a_4
XFILLER_162_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22644__A _22658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20463_ _22113_/A VGND VGND VPWR VPWR _20464_/A sky130_fd_sc_hd__buf_2
XANTENNA__22076__A2 _22074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23251_ _23347_/CLK _23251_/D VGND VGND VPWR VPWR _12173_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19477__B1 _20246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16642__A _16682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22202_ _22134_/X _22201_/X _15698_/B _22198_/X VGND VGND VPWR VPWR _23428_/D sky130_fd_sc_hd__o22a_4
XFILLER_146_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_21_0_HCLK clkbuf_4_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23182_ _23246_/CLK _23182_/D VGND VGND VPWR VPWR _16041_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21823__A2 _21815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20394_ _22420_/A VGND VGND VPWR VPWR _21821_/A sky130_fd_sc_hd__buf_2
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20164__A IRQ[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11786__A _16222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22133_ _22132_/X _22123_/X _13518_/B _22130_/X VGND VGND VPWR VPWR _23461_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19953__A _19953_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14162__A _12453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22064_ _22057_/A VGND VGND VPWR VPWR _22064_/X sky130_fd_sc_hd__buf_2
XFILLER_47_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21015_ _20344_/A _21014_/X _19126_/A _20269_/A VGND VGND VPWR VPWR _21015_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17473__A _17473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23473__CLK _23409_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21339__B2 _21338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12410__A _12410_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22966_ _22961_/A _22966_/B VGND VGND VPWR VPWR _22966_/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21917_ _21850_/X _21916_/X _15735_/B _21913_/X VGND VGND VPWR VPWR _21917_/X sky130_fd_sc_hd__o22a_4
XFILLER_70_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22897_ _22897_/A _22896_/X VGND VGND VPWR VPWR HWDATA[29] sky130_fd_sc_hd__nor2_4
XANTENNA__16817__A _16683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22411__A2_N _22409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15721__A _13099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12650_ _12650_/A VGND VGND VPWR VPWR _12941_/A sky130_fd_sc_hd__buf_2
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21848_ _21848_/A VGND VGND VPWR VPWR _21848_/X sky130_fd_sc_hd__buf_2
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20339__A _18780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19704__A1 _20844_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _17251_/A _17398_/A _17048_/A _18782_/B VGND VGND VPWR VPWR _17078_/C sky130_fd_sc_hd__or4_4
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _12581_/A VGND VGND VPWR VPWR _12600_/A sky130_fd_sc_hd__buf_2
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21779_ _21556_/X _21777_/X _23656_/Q _21774_/X VGND VGND VPWR VPWR _23656_/D sky130_fd_sc_hd__o22a_4
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21511__B2 _21510_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14320_ _11914_/A _14320_/B _14320_/C VGND VGND VPWR VPWR _14324_/B sky130_fd_sc_hd__and3_4
XFILLER_15_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ _24358_/Q _11532_/B VGND VGND VPWR VPWR _19030_/A sky130_fd_sc_hd__or2_4
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23518_ _23518_/CLK _23518_/D VGND VGND VPWR VPWR _13707_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24498_ _24472_/CLK _24498_/D HRESETn VGND VGND VPWR VPWR _19988_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17191__A1 _17140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14056__B _24064_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _14623_/A _23487_/Q VGND VGND VPWR VPWR _14251_/X sky130_fd_sc_hd__or2_4
XFILLER_156_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23449_ _24057_/CLK _22162_/X VGND VGND VPWR VPWR _14731_/B sky130_fd_sc_hd__dfxtp_4
X_13202_ _13232_/A _13199_/X _13202_/C VGND VGND VPWR VPWR _13202_/X sky130_fd_sc_hd__and3_4
X_14182_ _11720_/A VGND VGND VPWR VPWR _14226_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13133_ _12708_/A _13129_/X _13133_/C VGND VGND VPWR VPWR _13133_/X sky130_fd_sc_hd__or3_4
XFILLER_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15168__A _13589_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18990_ _19021_/A VGND VGND VPWR VPWR _18990_/X sky130_fd_sc_hd__buf_2
XANTENNA__14072__A _12329_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13064_ _13094_/A _12995_/B VGND VGND VPWR VPWR _13066_/B sky130_fd_sc_hd__or2_4
XFILLER_140_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17941_ _17833_/X _17936_/X _17811_/X _17940_/Y VGND VGND VPWR VPWR _17941_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19582__B _19788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23816__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12015_ _12015_/A _23892_/Q VGND VGND VPWR VPWR _12016_/C sky130_fd_sc_hd__or2_4
XFILLER_79_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19640__B1 HRDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17872_ _18413_/A VGND VGND VPWR VPWR _18562_/A sky130_fd_sc_hd__buf_2
XFILLER_120_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14800__A _14647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_41_0_HCLK clkbuf_6_20_0_HCLK/X VGND VGND VPWR VPWR _23246_/CLK sky130_fd_sc_hd__clkbuf_1
X_19611_ _20380_/B _19573_/X _19610_/X _19576_/X VGND VGND VPWR VPWR _19611_/X sky130_fd_sc_hd__a211o_4
XFILLER_94_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16823_ _16821_/A _16821_/B _16822_/Y VGND VGND VPWR VPWR _16823_/X sky130_fd_sc_hd__a21o_4
XFILLER_65_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13416__A _13416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19542_ _24170_/Q _19481_/X HRDATA[22] _19482_/X VGND VGND VPWR VPWR _19542_/X sky130_fd_sc_hd__o22a_4
X_16754_ _11742_/X VGND VGND VPWR VPWR _16759_/A sky130_fd_sc_hd__buf_2
X_13966_ _11931_/A _13966_/B _13965_/X VGND VGND VPWR VPWR _13966_/X sky130_fd_sc_hd__or3_4
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22729__A _22722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12917_ _12957_/A _12915_/X _12916_/X VGND VGND VPWR VPWR _12917_/X sky130_fd_sc_hd__and3_4
X_15705_ _11902_/A _15705_/B VGND VGND VPWR VPWR _15706_/C sky130_fd_sc_hd__or2_4
XANTENNA__13135__B _23783_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19943__B2 _19773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16685_ _11671_/X _16685_/B _16685_/C VGND VGND VPWR VPWR _16685_/X sky130_fd_sc_hd__and3_4
X_19473_ HRDATA[31] VGND VGND VPWR VPWR _20246_/B sky130_fd_sc_hd__buf_2
XFILLER_111_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13897_ _14507_/A _13897_/B VGND VGND VPWR VPWR _13898_/C sky130_fd_sc_hd__or2_4
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21750__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18424_ _17387_/Y _18424_/B VGND VGND VPWR VPWR _18424_/X sky130_fd_sc_hd__or2_4
XANTENNA__15631__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12848_ _12848_/A _12916_/B VGND VGND VPWR VPWR _12848_/X sky130_fd_sc_hd__or2_4
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15636_ _15612_/A _15634_/X _15635_/X VGND VGND VPWR VPWR _15636_/X sky130_fd_sc_hd__and3_4
XFILLER_61_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15567_ _14430_/A _24097_/Q VGND VGND VPWR VPWR _15568_/C sky130_fd_sc_hd__or2_4
X_18355_ _18307_/X _18354_/X _20047_/A _18307_/X VGND VGND VPWR VPWR _24486_/D sky130_fd_sc_hd__a2bb2o_4
X_12779_ _12778_/X VGND VGND VPWR VPWR _13343_/A sky130_fd_sc_hd__buf_2
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21502__B2 _21496_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13151__A _13338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14518_ _12401_/A _14516_/X _14518_/C VGND VGND VPWR VPWR _14518_/X sky130_fd_sc_hd__and3_4
X_17306_ _17306_/A VGND VGND VPWR VPWR _17308_/B sky130_fd_sc_hd__inv_2
XFILLER_148_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15498_ _12635_/A _15496_/X _15497_/X VGND VGND VPWR VPWR _15498_/X sky130_fd_sc_hd__and3_4
X_18286_ _17977_/X _17991_/Y _17985_/X _17996_/Y VGND VGND VPWR VPWR _18286_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22464__A _20818_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22058__A2 _22053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14449_ _14310_/A _14445_/X _14448_/X VGND VGND VPWR VPWR _14449_/X sky130_fd_sc_hd__or3_4
X_17237_ _17230_/X _17234_/X _17236_/X VGND VGND VPWR VPWR _17237_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16462__A _16362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23346__CLK _23204_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17168_ _17128_/X _17158_/X _17836_/A _17167_/X VGND VGND VPWR VPWR _17168_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16119_ _16144_/A _16117_/X _16119_/C VGND VGND VPWR VPWR _16120_/C sky130_fd_sc_hd__and3_4
XANTENNA__19773__A HRDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17099_ _17057_/B _18674_/A VGND VGND VPWR VPWR _17099_/Y sky130_fd_sc_hd__nor2_4
XFILLER_66_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21018__B1 _20662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21808__A _21808_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21569__B2 _21561_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15806__A _12867_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14710__A _12484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19809_ _19809_/A VGND VGND VPWR VPWR _19809_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22518__B1 _15511_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22820_ _22819_/X _15048_/X VGND VGND VPWR VPWR _22820_/X sky130_fd_sc_hd__or2_4
XFILLER_84_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22639__A _22672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19934__B2 _20422_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22751_ _22750_/Y _24125_/Q _22750_/Y _24125_/Q VGND VGND VPWR VPWR _22769_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15541__A _14431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21702_ _21596_/X _21698_/X _15179_/B _21667_/A VGND VGND VPWR VPWR _21702_/X sky130_fd_sc_hd__o22a_4
XFILLER_77_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22682_ _22478_/X _22679_/X _23128_/Q _22676_/X VGND VGND VPWR VPWR _23128_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24121__CLK _23544_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24421_ _23475_/CLK _18865_/X HRESETn VGND VGND VPWR VPWR _24421_/Q sky130_fd_sc_hd__dfrtp_4
X_21633_ _21563_/X _21627_/X _23749_/Q _21631_/X VGND VGND VPWR VPWR _23749_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15260__B _15260_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22297__A2 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19948__A _17816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14157__A _14269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24497__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24352_ _24382_/CLK _24352_/D HRESETn VGND VGND VPWR VPWR _24352_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__13982__A1 _13853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21564_ _21563_/X _21554_/X _23781_/Q _21561_/X VGND VGND VPWR VPWR _23781_/D sky130_fd_sc_hd__o22a_4
XFILLER_139_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23303_ _23303_/CLK _22379_/X VGND VGND VPWR VPWR _13208_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22049__A2 _22046_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20515_ _20343_/A VGND VGND VPWR VPWR _20515_/X sky130_fd_sc_hd__buf_2
X_24283_ _24287_/CLK _19308_/X HRESETn VGND VGND VPWR VPWR _24283_/Q sky130_fd_sc_hd__dfrtp_4
X_21495_ _21273_/X _21492_/X _23815_/Q _21489_/X VGND VGND VPWR VPWR _23815_/D sky130_fd_sc_hd__o22a_4
XFILLER_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24271__CLK _24271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23234_ _23303_/CLK _22518_/X VGND VGND VPWR VPWR _15511_/B sky130_fd_sc_hd__dfxtp_4
X_20446_ _20259_/A VGND VGND VPWR VPWR _20446_/X sky130_fd_sc_hd__buf_2
XFILLER_162_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23165_ _23229_/CLK _23165_/D VGND VGND VPWR VPWR _13900_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12405__A _12402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20377_ _20377_/A VGND VGND VPWR VPWR _21534_/A sky130_fd_sc_hd__buf_2
XFILLER_106_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22116_ _22115_/X _22111_/X _12259_/B _22106_/X VGND VGND VPWR VPWR _22116_/X sky130_fd_sc_hd__o22a_4
X_23096_ _23098_/CLK _23096_/D VGND VGND VPWR VPWR _15304_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22047_ _21813_/X _22046_/X _23507_/Q _22043_/X VGND VGND VPWR VPWR _23507_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22221__A2 _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23989__CLK _23203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_28_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21980__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13820_ _15411_/A _13818_/X _13819_/X VGND VGND VPWR VPWR _13820_/X sky130_fd_sc_hd__and3_4
X_23998_ _23496_/CLK _21171_/X VGND VGND VPWR VPWR _23998_/Q sky130_fd_sc_hd__dfxtp_4
X_13751_ _13751_/A _23966_/Q VGND VGND VPWR VPWR _13752_/C sky130_fd_sc_hd__or2_4
X_22949_ _22949_/A _18575_/X VGND VGND VPWR VPWR _22949_/X sky130_fd_sc_hd__or2_4
XANTENNA__21732__B2 _21731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12702_ _12702_/A VGND VGND VPWR VPWR _13279_/A sky130_fd_sc_hd__buf_2
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16470_ _16370_/X _16470_/B _16470_/C VGND VGND VPWR VPWR _16470_/X sky130_fd_sc_hd__or3_4
X_13682_ _12190_/A _13765_/B VGND VGND VPWR VPWR _13684_/B sky130_fd_sc_hd__or2_4
XFILLER_70_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15421_ _14480_/A _15398_/X _15405_/X _15412_/X _15420_/X VGND VGND VPWR VPWR _15421_/X
+ sky130_fd_sc_hd__a32o_4
X_12633_ _12953_/A _12631_/X _12633_/C VGND VGND VPWR VPWR _12633_/X sky130_fd_sc_hd__and3_4
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15170__B _15170_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22288__A2 _22287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23369__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15352_ _15328_/A _24056_/Q VGND VGND VPWR VPWR _15352_/X sky130_fd_sc_hd__or2_4
XFILLER_54_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18140_ _18113_/X _18120_/Y _18136_/X _18138_/Y _18139_/X VGND VGND VPWR VPWR _18140_/X
+ sky130_fd_sc_hd__a32o_4
X_12564_ _12499_/A _12564_/B VGND VGND VPWR VPWR _12566_/B sky130_fd_sc_hd__or2_4
XFILLER_19_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22284__A _22284_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ _13689_/A _14276_/X _14284_/X _14292_/X _14302_/X VGND VGND VPWR VPWR _14303_/X
+ sky130_fd_sc_hd__a32o_4
X_18071_ _18070_/A _16994_/B _18028_/Y VGND VGND VPWR VPWR _23049_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__24167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11515_ _24342_/Q _19126_/A VGND VGND VPWR VPWR _11515_/Y sky130_fd_sc_hd__nor2_4
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17378__A _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15283_ _12433_/A _23896_/Q VGND VGND VPWR VPWR _15285_/B sky130_fd_sc_hd__or2_4
XFILLER_106_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12495_ _12495_/A VGND VGND VPWR VPWR _13666_/A sky130_fd_sc_hd__buf_2
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17022_ _17021_/X VGND VGND VPWR VPWR _17022_/X sky130_fd_sc_hd__buf_2
XFILLER_172_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14234_ _14229_/A VGND VGND VPWR VPWR _14235_/A sky130_fd_sc_hd__buf_2
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21799__A1 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21799__B2 _21795_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14165_ _14165_/A _23103_/Q VGND VGND VPWR VPWR _14167_/B sky130_fd_sc_hd__or2_4
XFILLER_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13116_ _13088_/A _23496_/Q VGND VGND VPWR VPWR _13118_/B sky130_fd_sc_hd__or2_4
XFILLER_125_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18973_ _18963_/X _18971_/X _18972_/Y _18968_/X VGND VGND VPWR VPWR _18973_/X sky130_fd_sc_hd__o22a_4
X_14096_ _14096_/A VGND VGND VPWR VPWR _14137_/A sky130_fd_sc_hd__buf_2
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22748__B1 _23086_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13047_ _12882_/A _13024_/X _13031_/X _13038_/X _13046_/X VGND VGND VPWR VPWR _13047_/X
+ sky130_fd_sc_hd__a32o_4
X_17924_ _17923_/X VGND VGND VPWR VPWR _17924_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14530__A _11781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17419__A1_N _14086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17855_ _17850_/X _17237_/Y _17812_/X _17854_/Y VGND VGND VPWR VPWR _17855_/X sky130_fd_sc_hd__o22a_4
XFILLER_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16806_ _16621_/A _23729_/Q VGND VGND VPWR VPWR _16806_/X sky130_fd_sc_hd__or2_4
XFILLER_19_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17786_ _16935_/X _17651_/X _17653_/X _17785_/X VGND VGND VPWR VPWR _17786_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14998_ _13954_/A _14998_/B _14997_/X VGND VGND VPWR VPWR _14999_/C sky130_fd_sc_hd__and3_4
XFILLER_81_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22459__A _22459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19525_ _19525_/A VGND VGND VPWR VPWR _19682_/A sky130_fd_sc_hd__buf_2
XANTENNA__24144__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16737_ _12058_/A _16813_/B VGND VGND VPWR VPWR _16737_/X sky130_fd_sc_hd__or2_4
XFILLER_46_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13949_ _13949_/A VGND VGND VPWR VPWR _13949_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16457__A _11714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21723__B2 _21717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15361__A _15321_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19456_ _19455_/Y VGND VGND VPWR VPWR _19457_/A sky130_fd_sc_hd__buf_2
X_16668_ _16786_/A _16668_/B _16667_/X VGND VGND VPWR VPWR _16668_/X sky130_fd_sc_hd__and3_4
XANTENNA__20931__C1 _20930_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18407_ _18407_/A _17385_/X VGND VGND VPWR VPWR _18409_/C sky130_fd_sc_hd__nor2_4
XANTENNA__15080__B _23541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15619_ _11710_/A _15552_/B VGND VGND VPWR VPWR _15619_/X sky130_fd_sc_hd__or2_4
X_19387_ _19381_/X _19386_/X _19381_/X _24244_/Q VGND VGND VPWR VPWR _19387_/X sky130_fd_sc_hd__a2bb2o_4
X_16599_ _11876_/X _16599_/B _16599_/C VGND VGND VPWR VPWR _16600_/B sky130_fd_sc_hd__or3_4
XANTENNA__24294__CLK _24294_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18338_ _18338_/A VGND VGND VPWR VPWR _18338_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22194__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18269_ _18206_/X _18170_/X _18206_/X _18164_/X VGND VGND VPWR VPWR _18269_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20300_ _20210_/Y _20225_/X _20225_/X _20299_/X VGND VGND VPWR VPWR _24116_/D sky130_fd_sc_hd__a2bb2o_4
X_21280_ _21280_/A VGND VGND VPWR VPWR _21280_/X sky130_fd_sc_hd__buf_2
X_20231_ _20231_/A VGND VGND VPWR VPWR _20231_/X sky130_fd_sc_hd__buf_2
XFILLER_143_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12225__A _11935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20162_ IRQ[13] VGND VGND VPWR VPWR _20162_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22739__B1 _22736_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22203__A2 _22201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20093_ _11585_/X _11558_/X VGND VGND VPWR VPWR _20093_/X sky130_fd_sc_hd__or2_4
XANTENNA__14440__A _13010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23921_ _23761_/CLK _23921_/D VGND VGND VPWR VPWR _23921_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21527__A2_N _21525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21962__A1 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21962__B2 _21957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23852_ _23852_/CLK _23852_/D VGND VGND VPWR VPWR _12390_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_57_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22369__A _22376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22803_ _22802_/X VGND VGND VPWR VPWR _22803_/X sky130_fd_sc_hd__buf_2
XFILLER_77_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23783_ _23750_/CLK _23783_/D VGND VGND VPWR VPWR _23783_/Q sky130_fd_sc_hd__dfxtp_4
X_20995_ _20781_/X _20994_/X _24310_/Q _20791_/X VGND VGND VPWR VPWR _20996_/B sky130_fd_sc_hd__o22a_4
XANTENNA__21714__B2 _21710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15271__A _12453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22734_ _21313_/A _22729_/X _14902_/B _22698_/A VGND VGND VPWR VPWR _23094_/D sky130_fd_sc_hd__o22a_4
XFILLER_129_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16086__B _16085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22665_ _22658_/A VGND VGND VPWR VPWR _22665_/X sky130_fd_sc_hd__buf_2
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24404_ _23409_/CLK _24404_/D HRESETn VGND VGND VPWR VPWR _24404_/Q sky130_fd_sc_hd__dfstp_4
X_21616_ _21534_/X _21613_/X _23761_/Q _21610_/X VGND VGND VPWR VPWR _23761_/D sky130_fd_sc_hd__o22a_4
XFILLER_138_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22596_ _22416_/X _22594_/X _16638_/B _22591_/X VGND VGND VPWR VPWR _22596_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24335_ _24277_/CLK _24335_/D HRESETn VGND VGND VPWR VPWR _19156_/A sky130_fd_sc_hd__dfrtp_4
X_21547_ _21546_/X _21542_/X _23788_/Q _21537_/X VGND VGND VPWR VPWR _21547_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14615__A _14615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12280_ _12240_/A VGND VGND VPWR VPWR _13300_/A sky130_fd_sc_hd__buf_2
X_24266_ _24495_/CLK _19349_/X HRESETn VGND VGND VPWR VPWR _20526_/A sky130_fd_sc_hd__dfrtp_4
X_21478_ _21492_/A VGND VGND VPWR VPWR _21478_/X sky130_fd_sc_hd__buf_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23217_ _23537_/CLK _23217_/D VGND VGND VPWR VPWR _16761_/B sky130_fd_sc_hd__dfxtp_4
X_20429_ _18891_/X VGND VGND VPWR VPWR _20429_/X sky130_fd_sc_hd__buf_2
XANTENNA__24017__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24197_ _23991_/CLK _19790_/X HRESETn VGND VGND VPWR VPWR _11750_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21448__A _21441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23148_ _23500_/CLK _22654_/X VGND VGND VPWR VPWR _12389_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11974__A _16138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15446__A _15446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15970_ _15993_/A _15967_/X _15970_/C VGND VGND VPWR VPWR _15970_/X sky130_fd_sc_hd__and3_4
X_23079_ _19975_/X _23079_/B VGND VGND VPWR VPWR _23080_/C sky130_fd_sc_hd__or2_4
XFILLER_0_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24167__CLK _23991_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14921_ _15369_/A _14921_/B _14920_/X VGND VGND VPWR VPWR _14921_/X sky130_fd_sc_hd__or3_4
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17640_ _17640_/A _17599_/X _17640_/C _17640_/D VGND VGND VPWR VPWR _17640_/X sky130_fd_sc_hd__and4_4
X_14852_ _14096_/A _14852_/B VGND VGND VPWR VPWR _14852_/X sky130_fd_sc_hd__or2_4
XFILLER_91_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22279__A _22275_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13803_ _14307_/A _13876_/B VGND VGND VPWR VPWR _13803_/X sky130_fd_sc_hd__or2_4
X_14783_ _15330_/A VGND VGND VPWR VPWR _14783_/X sky130_fd_sc_hd__buf_2
X_17571_ _17571_/A VGND VGND VPWR VPWR _17572_/B sky130_fd_sc_hd__inv_2
XFILLER_17_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11995_ _11943_/X _11993_/X _11995_/C VGND VGND VPWR VPWR _11999_/B sky130_fd_sc_hd__and3_4
XANTENNA__16277__A _11971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19310_ _19231_/A _19230_/X _19309_/Y VGND VGND VPWR VPWR _24282_/D sky130_fd_sc_hd__o21a_4
XFILLER_1_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15181__A _15018_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13734_ _13774_/A _13732_/X _13734_/C VGND VGND VPWR VPWR _13734_/X sky130_fd_sc_hd__and3_4
XFILLER_21_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16522_ _16521_/X VGND VGND VPWR VPWR _16523_/B sky130_fd_sc_hd__buf_2
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21181__A2 _21176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19241_ _24292_/Q _19240_/X VGND VGND VPWR VPWR _19289_/A sky130_fd_sc_hd__and2_4
X_16453_ _11715_/A _16387_/B VGND VGND VPWR VPWR _16455_/B sky130_fd_sc_hd__or2_4
XANTENNA__19588__A _19539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13665_ _13622_/A VGND VGND VPWR VPWR _15408_/A sky130_fd_sc_hd__buf_2
XFILLER_108_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12616_ _12616_/A VGND VGND VPWR VPWR _12962_/A sky130_fd_sc_hd__buf_2
X_15404_ _15404_/A _15404_/B _15403_/X VGND VGND VPWR VPWR _15405_/C sky130_fd_sc_hd__and3_4
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19172_ _19156_/A _19156_/B _19171_/Y VGND VGND VPWR VPWR _24335_/D sky130_fd_sc_hd__o21a_4
X_16384_ _16309_/X _16383_/A VGND VGND VPWR VPWR _16384_/X sky130_fd_sc_hd__or2_4
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ _13596_/A VGND VGND VPWR VPWR _14311_/A sky130_fd_sc_hd__buf_2
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15335_ _13699_/A _23160_/Q VGND VGND VPWR VPWR _15337_/B sky130_fd_sc_hd__or2_4
X_18123_ _17849_/X _18122_/Y VGND VGND VPWR VPWR _18123_/X sky130_fd_sc_hd__or2_4
X_12547_ _12911_/A VGND VGND VPWR VPWR _12874_/A sky130_fd_sc_hd__buf_2
XFILLER_129_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18885__A1 _16866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22681__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14525__A _12410_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20246__B _20246_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15266_ _12287_/A _15262_/X _15266_/C VGND VGND VPWR VPWR _15266_/X sky130_fd_sc_hd__or3_4
X_18054_ _17874_/X _18052_/X _18053_/X VGND VGND VPWR VPWR _18054_/Y sky130_fd_sc_hd__o21ai_4
X_12478_ _12537_/A VGND VGND VPWR VPWR _12878_/A sky130_fd_sc_hd__buf_2
XANTENNA__14244__B _23103_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17005_ _17005_/A VGND VGND VPWR VPWR _17005_/X sky130_fd_sc_hd__buf_2
X_14217_ _14201_/A _14217_/B _14217_/C VGND VGND VPWR VPWR _14221_/B sky130_fd_sc_hd__and3_4
X_15197_ _15196_/X _15134_/B VGND VGND VPWR VPWR _15200_/B sky130_fd_sc_hd__or2_4
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14148_ _14148_/A _23423_/Q VGND VGND VPWR VPWR _14148_/X sky130_fd_sc_hd__or2_4
XFILLER_99_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18956_ _18948_/D VGND VGND VPWR VPWR _19009_/A sky130_fd_sc_hd__inv_2
X_14079_ _12329_/A _23648_/Q VGND VGND VPWR VPWR _14080_/C sky130_fd_sc_hd__or2_4
XFILLER_140_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24355__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14260__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22197__B2 _22191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17907_ _17904_/X _17964_/B _17903_/A VGND VGND VPWR VPWR _17908_/B sky130_fd_sc_hd__o21ai_4
XFILLER_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18887_ _12028_/X _16710_/A VGND VGND VPWR VPWR _18887_/X sky130_fd_sc_hd__or2_4
XANTENNA__18667__A _18399_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21944__B2 _21943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23534__CLK _23246_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_11_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_82_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17838_ _17838_/A VGND VGND VPWR VPWR _17838_/X sky130_fd_sc_hd__buf_2
XFILLER_54_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17769_ _17675_/X _17702_/X VGND VGND VPWR VPWR _17769_/X sky130_fd_sc_hd__or2_4
XANTENNA__16187__A _16187_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ _19508_/A VGND VGND VPWR VPWR _19675_/A sky130_fd_sc_hd__inv_2
XANTENNA__15091__A _15091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13604__A _15415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20780_ _20233_/Y VGND VGND VPWR VPWR _20780_/X sky130_fd_sc_hd__buf_2
XANTENNA__21172__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22917__A _22916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19439_ _19439_/A VGND VGND VPWR VPWR _19512_/A sky130_fd_sc_hd__inv_2
XFILLER_23_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22450_ _22438_/A VGND VGND VPWR VPWR _22450_/X sky130_fd_sc_hd__buf_2
XFILLER_148_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22121__B2 _22118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21401_ _21285_/X _21398_/X _15505_/B _21395_/X VGND VGND VPWR VPWR _23874_/D sky130_fd_sc_hd__o22a_4
X_22381_ _22129_/X _22376_/X _23302_/Q _22380_/X VGND VGND VPWR VPWR _22381_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18876__A1 _17272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14435__A _12461_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24120_ _23544_/CLK _22780_/X HRESETn VGND VGND VPWR VPWR _22753_/A sky130_fd_sc_hd__dfrtp_4
X_21332_ _21251_/X _21327_/X _16421_/B _21331_/X VGND VGND VPWR VPWR _21332_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14154__B _23487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24051_ _23889_/CLK _21091_/X VGND VGND VPWR VPWR _24051_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_163_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21263_ _20509_/A VGND VGND VPWR VPWR _21263_/X sky130_fd_sc_hd__buf_2
XANTENNA__22424__A2 _22414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16650__A _16678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20435__A1 _18101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23002_ _22910_/X VGND VGND VPWR VPWR _23003_/B sky130_fd_sc_hd__buf_2
X_20214_ _21603_/A _21028_/A _21133_/A _21234_/A VGND VGND VPWR VPWR _20214_/X sky130_fd_sc_hd__or4_4
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21194_ _20378_/X _21191_/X _23985_/Q _21188_/X VGND VGND VPWR VPWR _21194_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11794__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15266__A _12287_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20145_ _20145_/A VGND VGND VPWR VPWR _20145_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14170__A _14170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22188__B2 _22184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20076_ _18530_/X _20055_/X _20075_/Y _20066_/X VGND VGND VPWR VPWR _20076_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20900__A HRDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21935__B2 _21899_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17064__B1 _20216_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17481__A _11876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18800__A1 _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23904_ _23904_/CLK _23904_/D VGND VGND VPWR VPWR _14052_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22099__A _22123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23835_ _23515_/CLK _21461_/X VGND VGND VPWR VPWR _14460_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11780_/A VGND VGND VPWR VPWR _11781_/A sky130_fd_sc_hd__buf_2
X_23766_ _23770_/CLK _23766_/D VGND VGND VPWR VPWR _23766_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20978_ _24215_/Q _20895_/X _20977_/Y VGND VGND VPWR VPWR _22480_/A sky130_fd_sc_hd__o21a_4
XANTENNA__21163__A2 _21162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22360__B2 _22359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21731__A _21724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22717_ _21283_/A _22715_/X _15840_/B _22712_/X VGND VGND VPWR VPWR _22717_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23697_ _23761_/CLK _23697_/D VGND VGND VPWR VPWR _23697_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ _12868_/A _13518_/B VGND VGND VPWR VPWR _13451_/C sky130_fd_sc_hd__or2_4
XFILLER_55_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22648_ _22648_/A VGND VGND VPWR VPWR _22648_/X sky130_fd_sc_hd__buf_2
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20347__A _20270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22112__B2 _22106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12401_ _12401_/A VGND VGND VPWR VPWR _12950_/A sky130_fd_sc_hd__buf_2
XANTENNA__11969__A _11969_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13381_ _13399_/A _13381_/B _13381_/C VGND VGND VPWR VPWR _13382_/C sky130_fd_sc_hd__or3_4
XANTENNA__18867__A1 _15916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22663__A2 _22658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22579_ _22539_/A VGND VGND VPWR VPWR _22579_/X sky130_fd_sc_hd__buf_2
X_15120_ _15048_/X _15116_/X _15119_/X VGND VGND VPWR VPWR _15120_/Y sky130_fd_sc_hd__o21ai_4
X_12332_ _12829_/A _23532_/Q VGND VGND VPWR VPWR _12332_/X sky130_fd_sc_hd__or2_4
X_24318_ _24292_/CLK _19206_/X HRESETn VGND VGND VPWR VPWR _24318_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17078__D _18888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15051_ _12329_/A _23509_/Q VGND VGND VPWR VPWR _15052_/C sky130_fd_sc_hd__or2_4
XFILLER_147_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12263_ _12912_/A _12208_/X _12225_/X _12247_/X _12262_/X VGND VGND VPWR VPWR _12263_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18619__A1 _16927_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24249_ _24248_/CLK _24249_/D HRESETn VGND VGND VPWR VPWR _24249_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22415__A2 _22414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14002_ _13637_/A _23648_/Q VGND VGND VPWR VPWR _14003_/C sky130_fd_sc_hd__or2_4
X_12194_ _12194_/A VGND VGND VPWR VPWR _12501_/A sky130_fd_sc_hd__buf_2
XANTENNA__15176__A _14988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18810_ _18786_/A VGND VGND VPWR VPWR _18810_/X sky130_fd_sc_hd__buf_2
XFILLER_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19790_ _19732_/X _19785_/X _19789_/X _16675_/A _19719_/X VGND VGND VPWR VPWR _19790_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14080__A _11698_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21906__A _21906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18741_ _17752_/X _17753_/X _17752_/X _17753_/X VGND VGND VPWR VPWR _18741_/X sky130_fd_sc_hd__a2bb2o_4
X_15953_ _13330_/A VGND VGND VPWR VPWR _16006_/A sky130_fd_sc_hd__buf_2
XFILLER_27_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21926__B2 _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14904_ _13591_/A _14902_/X _14903_/X VGND VGND VPWR VPWR _14904_/X sky130_fd_sc_hd__and3_4
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18672_ _18517_/A _17315_/Y VGND VGND VPWR VPWR _18674_/B sky130_fd_sc_hd__or2_4
X_15884_ _15903_/A _15822_/B VGND VGND VPWR VPWR _15884_/X sky130_fd_sc_hd__or2_4
XFILLER_110_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17623_ _17623_/A VGND VGND VPWR VPWR _18714_/B sky130_fd_sc_hd__inv_2
X_14835_ _14823_/A _14751_/B VGND VGND VPWR VPWR _14835_/X sky130_fd_sc_hd__or2_4
XFILLER_64_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13424__A _13327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17554_ _17971_/B _17554_/B VGND VGND VPWR VPWR _17641_/A sky130_fd_sc_hd__or2_4
X_14766_ _13951_/X _11627_/A _14735_/X _11604_/A _14765_/X VGND VGND VPWR VPWR _14766_/X
+ sky130_fd_sc_hd__a32o_4
X_11978_ _11975_/A _11793_/B VGND VGND VPWR VPWR _11978_/X sky130_fd_sc_hd__or2_4
XANTENNA__21154__A2 _21148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22737__A _22737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16505_ _16479_/X _16442_/B VGND VGND VPWR VPWR _16505_/X sky130_fd_sc_hd__or2_4
XANTENNA__24182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21641__A _21608_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13717_ _13717_/A VGND VGND VPWR VPWR _15372_/A sky130_fd_sc_hd__buf_2
X_17485_ _12680_/X _17487_/B VGND VGND VPWR VPWR _17485_/X sky130_fd_sc_hd__or2_4
X_14697_ _15625_/A _14697_/B _14696_/X VGND VGND VPWR VPWR _14697_/X sky130_fd_sc_hd__or3_4
XFILLER_71_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19224_ _19131_/B VGND VGND VPWR VPWR _19224_/Y sky130_fd_sc_hd__inv_2
X_16436_ _16101_/A _16436_/B VGND VGND VPWR VPWR _16436_/X sky130_fd_sc_hd__or2_4
X_13648_ _11878_/A _13646_/X _13648_/C VGND VGND VPWR VPWR _13648_/X sky130_fd_sc_hd__and3_4
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19155_ _19155_/A _19155_/B VGND VGND VPWR VPWR _19156_/B sky130_fd_sc_hd__and2_4
XANTENNA__18858__A1 _17156_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16367_ _16454_/A _16304_/B VGND VGND VPWR VPWR _16367_/X sky130_fd_sc_hd__or2_4
XANTENNA__22654__A2 _22651_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13579_ _12422_/A _12682_/Y _12423_/A _13578_/Y VGND VGND VPWR VPWR _13580_/A sky130_fd_sc_hd__a211o_4
XANTENNA__14255__A _15606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_2_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18106_ _18068_/X _18105_/X _20008_/A _18068_/X VGND VGND VPWR VPWR _24494_/D sky130_fd_sc_hd__a2bb2o_4
X_15318_ _15318_/A _23352_/Q VGND VGND VPWR VPWR _15318_/X sky130_fd_sc_hd__or2_4
X_16298_ _15961_/A _16296_/X _16297_/X VGND VGND VPWR VPWR _16298_/X sky130_fd_sc_hd__and3_4
X_19086_ _19082_/X _19085_/X _19082_/X _11524_/A VGND VGND VPWR VPWR _19086_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17566__A _11611_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18037_ _18376_/A VGND VGND VPWR VPWR _18037_/X sky130_fd_sc_hd__buf_2
X_15249_ _11812_/A _15233_/X _15248_/X VGND VGND VPWR VPWR _15250_/C sky130_fd_sc_hd__or3_4
XANTENNA__16470__A _16370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20417__A1 _20302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20417__B2 _20396_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14702__B _14701_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12503__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19988_ _19988_/A VGND VGND VPWR VPWR _19988_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24482__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18939_ _15380_/A _18934_/X _24376_/Q _18935_/X VGND VGND VPWR VPWR _18939_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21917__B2 _21913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15814__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21950_ _21950_/A VGND VGND VPWR VPWR _21950_/X sky130_fd_sc_hd__buf_2
XFILLER_39_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21393__A2 _21391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18794__B1 _24465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20901_ _20900_/Y _20873_/X _20512_/B _20697_/X VGND VGND VPWR VPWR _20901_/X sky130_fd_sc_hd__a2bb2o_4
X_21881_ _21311_/A VGND VGND VPWR VPWR _21881_/X sky130_fd_sc_hd__buf_2
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23620_ _23303_/CLK _23620_/D VGND VGND VPWR VPWR _15755_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_82_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20832_ _20781_/X _20831_/X _24317_/Q _20791_/X VGND VGND VPWR VPWR _20832_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17349__A1 _15382_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18546__B1 _17792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21551__A _20531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23551_ _23582_/CLK _23551_/D VGND VGND VPWR VPWR _23551_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20763_ _20652_/A _20762_/X VGND VGND VPWR VPWR _20763_/Y sky130_fd_sc_hd__nor2_4
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22502_ _22425_/X _22501_/X _16000_/B _22498_/X VGND VGND VPWR VPWR _23246_/D sky130_fd_sc_hd__o22a_4
XFILLER_22_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_18_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR _24158_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23482_ _23515_/CLK _22082_/X VGND VGND VPWR VPWR _14597_/B sky130_fd_sc_hd__dfxtp_4
X_20694_ _20635_/X _20693_/X _15834_/B _20614_/X VGND VGND VPWR VPWR _20694_/X sky130_fd_sc_hd__o22a_4
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22433_ _22433_/A VGND VGND VPWR VPWR _22433_/X sky130_fd_sc_hd__buf_2
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19956__A _19956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14165__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22645__A2 _22644_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22364_ _22101_/X _22362_/X _16627_/B _22359_/X VGND VGND VPWR VPWR _22364_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17521__A1 _17518_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17521__B2 _17520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24103_ _24039_/CLK _20597_/X VGND VGND VPWR VPWR _24103_/Q sky130_fd_sc_hd__dfxtp_4
X_21315_ _21024_/A VGND VGND VPWR VPWR _21315_/X sky130_fd_sc_hd__buf_2
X_22295_ _22122_/X _22294_/X _23369_/Q _22291_/X VGND VGND VPWR VPWR _22295_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16380__A _13417_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24034_ _23587_/CLK _21114_/X VGND VGND VPWR VPWR _15465_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_137_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21246_ _21243_/X _21245_/X _23955_/Q _21240_/X VGND VGND VPWR VPWR _21246_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12413__A _15851_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21177_ _20915_/X _21176_/X _14568_/B _21173_/X VGND VGND VPWR VPWR _23994_/D sky130_fd_sc_hd__o22a_4
XFILLER_77_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20128_ _20194_/A _20127_/X _11636_/A VGND VGND VPWR VPWR _20128_/X sky130_fd_sc_hd__o21a_4
XFILLER_104_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20630__A _20535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21908__B2 _21906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12950_ _12950_/A _12948_/X _12950_/C VGND VGND VPWR VPWR _12950_/X sky130_fd_sc_hd__and3_4
XANTENNA__15724__A _12766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22030__B1 _14485_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20059_ _20058_/X VGND VGND VPWR VPWR _24146_/D sky130_fd_sc_hd__inv_2
X_11901_ _12854_/A VGND VGND VPWR VPWR _11902_/A sky130_fd_sc_hd__buf_2
XANTENNA__22581__B2 _22576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12881_ _12881_/A _12877_/X _12881_/C VGND VGND VPWR VPWR _12882_/B sky130_fd_sc_hd__or3_4
XANTENNA__15443__B _15501_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13244__A _12354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ _11832_/A _23124_/Q VGND VGND VPWR VPWR _11834_/B sky130_fd_sc_hd__or2_4
XANTENNA__24205__CLK _23126_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14620_ _14820_/A _23514_/Q VGND VGND VPWR VPWR _14621_/C sky130_fd_sc_hd__or2_4
X_23818_ _23852_/CLK _23818_/D VGND VGND VPWR VPWR _12825_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18754__B _11633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14059__B _23136_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14483_/Y _14548_/X _15389_/B VGND VGND VPWR VPWR _14552_/A sky130_fd_sc_hd__o21a_4
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23749_ _23493_/CLK _23749_/D VGND VGND VPWR VPWR _23749_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11763_ _11717_/X _11763_/B VGND VGND VPWR VPWR _11763_/X sky130_fd_sc_hd__or2_4
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _12402_/X _13500_/X _13501_/X VGND VGND VPWR VPWR _13502_/X sky130_fd_sc_hd__and3_4
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _11855_/A _11629_/A _14451_/X _11606_/A _14481_/X VGND VGND VPWR VPWR _14482_/X
+ sky130_fd_sc_hd__a32o_4
X_17270_ _17915_/B _17269_/Y VGND VGND VPWR VPWR _17911_/B sky130_fd_sc_hd__or2_4
X_11694_ _11693_/X VGND VGND VPWR VPWR _11694_/X sky130_fd_sc_hd__buf_2
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16221_ _16205_/A _16221_/B _16221_/C VGND VGND VPWR VPWR _16222_/C sky130_fd_sc_hd__or3_4
X_13433_ _13330_/A _13433_/B _13433_/C VGND VGND VPWR VPWR _13434_/C sky130_fd_sc_hd__and3_4
XANTENNA__11699__A _12604_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24355__CLK _24388_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16152_ _16138_/A _16152_/B _16151_/X VGND VGND VPWR VPWR _16152_/X sky130_fd_sc_hd__or3_4
XFILLER_139_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13364_ _13374_/A _13364_/B VGND VGND VPWR VPWR _13366_/B sky130_fd_sc_hd__or2_4
XFILLER_10_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17512__A1 _13049_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17512__B2 _17511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12315_ _12748_/A _12315_/B _12315_/C VGND VGND VPWR VPWR _12316_/C sky130_fd_sc_hd__and3_4
X_15103_ _15103_/A _23701_/Q VGND VGND VPWR VPWR _15105_/B sky130_fd_sc_hd__or2_4
X_16083_ _16187_/A _16083_/B _16082_/X VGND VGND VPWR VPWR _16083_/X sky130_fd_sc_hd__and3_4
X_13295_ _13330_/A _13292_/X _13294_/X VGND VGND VPWR VPWR _13295_/X sky130_fd_sc_hd__and3_4
XFILLER_127_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14803__A _14669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19911_ _19906_/X _20871_/A _19910_/X VGND VGND VPWR VPWR _19911_/Y sky130_fd_sc_hd__o21ai_4
X_15034_ _13630_/A _23637_/Q VGND VGND VPWR VPWR _15035_/C sky130_fd_sc_hd__or2_4
XFILLER_154_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12246_ _12298_/A _12241_/X _12246_/C VGND VGND VPWR VPWR _12247_/C sky130_fd_sc_hd__and3_4
XANTENNA__13419__A _13455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21072__B2 _21070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19842_ _19842_/A VGND VGND VPWR VPWR _19842_/Y sky130_fd_sc_hd__inv_2
X_12177_ _11686_/X _12177_/B _12176_/X VGND VGND VPWR VPWR _12178_/C sky130_fd_sc_hd__and3_4
XANTENNA__12323__A _13052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19773_ HRDATA[18] VGND VGND VPWR VPWR _19773_/X sky130_fd_sc_hd__buf_2
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16985_ _17905_/A _17906_/B VGND VGND VPWR VPWR _16985_/X sky130_fd_sc_hd__or2_4
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18724_ _18721_/Y _18723_/X _18721_/Y _18723_/X VGND VGND VPWR VPWR _18724_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15936_ _11882_/X VGND VGND VPWR VPWR _15936_/X sky130_fd_sc_hd__buf_2
XFILLER_7_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18655_ _18654_/X VGND VGND VPWR VPWR _18655_/Y sky130_fd_sc_hd__inv_2
X_15867_ _13514_/A _15865_/X _15866_/X VGND VGND VPWR VPWR _15867_/X sky130_fd_sc_hd__and3_4
XFILLER_58_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17606_ _17362_/X _17371_/A _17375_/B VGND VGND VPWR VPWR _17606_/X sky130_fd_sc_hd__a21o_4
X_14818_ _14840_/A _14814_/X _14818_/C VGND VGND VPWR VPWR _14826_/B sky130_fd_sc_hd__or3_4
XFILLER_91_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18586_ _18518_/A _17401_/X _17797_/A VGND VGND VPWR VPWR _18586_/X sky130_fd_sc_hd__a21o_4
X_15798_ _13324_/A _15796_/X _15797_/X VGND VGND VPWR VPWR _15798_/X sky130_fd_sc_hd__and3_4
XANTENNA__21127__A2 _21125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17537_ _17475_/B VGND VGND VPWR VPWR _17537_/Y sky130_fd_sc_hd__inv_2
X_14749_ _14331_/A _14745_/X _14749_/C VGND VGND VPWR VPWR _14749_/X sky130_fd_sc_hd__or3_4
XANTENNA__12993__A _12877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17468_ _17467_/X VGND VGND VPWR VPWR _17468_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14014__B1 _11603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19207_ _19138_/X VGND VGND VPWR VPWR _19207_/Y sky130_fd_sc_hd__inv_2
X_16419_ _11971_/X _16419_/B VGND VGND VPWR VPWR _16419_/X sky130_fd_sc_hd__and2_4
XFILLER_73_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19776__A _19705_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17399_ _17398_/Y _17280_/B VGND VGND VPWR VPWR _17399_/X sky130_fd_sc_hd__or2_4
XFILLER_146_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21835__B1 _12646_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19138_ _24317_/Q _19138_/B VGND VGND VPWR VPWR _19138_/X sky130_fd_sc_hd__and2_4
XFILLER_173_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17296__A _17296_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15809__A _12874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19069_ _19052_/X _19067_/X _19068_/X _19063_/A VGND VGND VPWR VPWR _24353_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14713__A _13596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21100_ _20486_/X _21097_/X _24044_/Q _21094_/X VGND VGND VPWR VPWR _24044_/D sky130_fd_sc_hd__o22a_4
XFILLER_172_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22080_ _21872_/X _22074_/X _23483_/Q _22078_/X VGND VGND VPWR VPWR _22080_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22930__A _22930_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21031_ _21184_/A _21134_/B _21184_/C _21134_/D VGND VGND VPWR VPWR _21031_/X sky130_fd_sc_hd__or4_4
XANTENNA__22260__B1 _13760_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21546__A _20486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15544__A _14421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24228__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22982_ _22977_/X _18367_/A _22959_/X _22981_/X VGND VGND VPWR VPWR _22982_/X sky130_fd_sc_hd__a211o_4
XFILLER_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21366__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22563__B2 _22562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21933_ _21879_/X _21930_/X _15333_/B _21927_/X VGND VGND VPWR VPWR _23576_/D sky130_fd_sc_hd__o22a_4
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13064__A _13094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21864_ _21862_/X _21863_/X _23615_/Q _21858_/X VGND VGND VPWR VPWR _21864_/X sky130_fd_sc_hd__o22a_4
XFILLER_167_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21281__A _21269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23603_ _23764_/CLK _21896_/X VGND VGND VPWR VPWR _23603_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23252__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20815_ _20695_/X _20806_/Y _20813_/X _20814_/Y _20714_/X VGND VGND VPWR VPWR _20815_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21795_ _21774_/A VGND VGND VPWR VPWR _21795_/X sky130_fd_sc_hd__buf_2
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23534_ _23246_/CLK _22004_/X VGND VGND VPWR VPWR _15940_/B sky130_fd_sc_hd__dfxtp_4
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20746_ _20510_/A VGND VGND VPWR VPWR _20746_/X sky130_fd_sc_hd__buf_2
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23465_ _23337_/CLK _22124_/X VGND VGND VPWR VPWR _23465_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20677_ _20677_/A _20617_/B VGND VGND VPWR VPWR _20677_/Y sky130_fd_sc_hd__nand2_4
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22416_ _20360_/A VGND VGND VPWR VPWR _22416_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23396_ _23588_/CLK _23396_/D VGND VGND VPWR VPWR _15762_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_104_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23001__A _23043_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22347_ _23323_/Q VGND VGND VPWR VPWR _23323_/D sky130_fd_sc_hd__buf_2
XANTENNA__15719__A _12758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12319__B1 _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12100_ _12061_/A _12098_/X _12100_/C VGND VGND VPWR VPWR _12100_/X sky130_fd_sc_hd__and3_4
X_13080_ _13055_/A VGND VGND VPWR VPWR _13089_/A sky130_fd_sc_hd__buf_2
X_22278_ _22272_/Y _22277_/X _22095_/X _22277_/X VGND VGND VPWR VPWR _23380_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24017_ _23761_/CLK _24017_/D VGND VGND VPWR VPWR _24017_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12031_ _16711_/A VGND VGND VPWR VPWR _16700_/A sky130_fd_sc_hd__buf_2
XANTENNA__21054__B2 _21049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21229_ _20959_/X _21226_/X _23960_/Q _21223_/X VGND VGND VPWR VPWR _21229_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20360__A _20360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11982__A _11973_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16770_ _16755_/X _23953_/Q VGND VGND VPWR VPWR _16772_/B sky130_fd_sc_hd__or2_4
X_13982_ _13853_/A _13959_/X _13966_/X _13973_/X _13981_/X VGND VGND VPWR VPWR _13982_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21357__A2 _21355_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22554__B2 _22548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15721_ _13099_/A _15719_/X _15720_/X VGND VGND VPWR VPWR _15721_/X sky130_fd_sc_hd__and3_4
X_12933_ _12940_/A _23593_/Q VGND VGND VPWR VPWR _12933_/X sky130_fd_sc_hd__or2_4
XFILLER_160_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18765__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18440_ _18440_/A _17394_/A VGND VGND VPWR VPWR _18440_/X sky130_fd_sc_hd__and2_4
XANTENNA__13047__A1 _12882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15652_ _15651_/X VGND VGND VPWR VPWR _15652_/Y sky130_fd_sc_hd__inv_2
X_12864_ _12864_/A _23305_/Q VGND VGND VPWR VPWR _12865_/C sky130_fd_sc_hd__or2_4
XANTENNA__21109__A2 _21104_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22287__A _22294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18484__B _17445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22306__B2 _22305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21191__A _21198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14603_ _11933_/A _14599_/X _14602_/X VGND VGND VPWR VPWR _14603_/X sky130_fd_sc_hd__or3_4
X_11815_ _13416_/A VGND VGND VPWR VPWR _11815_/X sky130_fd_sc_hd__buf_2
X_18371_ _18370_/X VGND VGND VPWR VPWR _18371_/Y sky130_fd_sc_hd__inv_2
X_12795_ _13205_/A VGND VGND VPWR VPWR _15778_/A sky130_fd_sc_hd__buf_2
X_15583_ _11710_/A _15522_/B VGND VGND VPWR VPWR _15585_/B sky130_fd_sc_hd__or2_4
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17322_ _17319_/Y _17018_/X _17026_/X _17321_/X VGND VGND VPWR VPWR _17324_/B sky130_fd_sc_hd__o22a_4
X_14534_ _14510_/A _14534_/B VGND VGND VPWR VPWR _14536_/B sky130_fd_sc_hd__or2_4
X_11746_ _16080_/A VGND VGND VPWR VPWR _11746_/X sky130_fd_sc_hd__buf_2
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _16687_/A _17024_/X _17031_/X _17252_/Y VGND VGND VPWR VPWR _17253_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22609__A2 _22608_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11677_ _13530_/A VGND VGND VPWR VPWR _13383_/A sky130_fd_sc_hd__buf_2
X_14465_ _12546_/A _14461_/X _14464_/X VGND VGND VPWR VPWR _14465_/X sky130_fd_sc_hd__or3_4
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16204_ _16220_/A _16202_/X _16204_/C VGND VGND VPWR VPWR _16205_/C sky130_fd_sc_hd__and3_4
X_13416_ _13416_/A _13416_/B _13415_/X VGND VGND VPWR VPWR _13417_/C sky130_fd_sc_hd__or3_4
Xclkbuf_7_64_0_HCLK clkbuf_7_65_0_HCLK/A VGND VGND VPWR VPWR _24137_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17184_ _17015_/X _17131_/X _17339_/A _17133_/X VGND VGND VPWR VPWR _17184_/X sky130_fd_sc_hd__o22a_4
X_14396_ _14366_/A _14396_/B VGND VGND VPWR VPWR _14396_/X sky130_fd_sc_hd__or2_4
X_16135_ _16108_/A _23629_/Q VGND VGND VPWR VPWR _16135_/X sky130_fd_sc_hd__or2_4
X_13347_ _13385_/A _13274_/B VGND VGND VPWR VPWR _13347_/X sky130_fd_sc_hd__or2_4
XFILLER_128_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16066_ _16066_/A _16064_/X _16066_/C VGND VGND VPWR VPWR _16067_/C sky130_fd_sc_hd__and3_4
X_13278_ _13309_/A _23366_/Q VGND VGND VPWR VPWR _13281_/B sky130_fd_sc_hd__or2_4
XANTENNA__22750__A SYSTICKCLKDIV[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14252__B _24095_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22242__B1 _12655_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12229_ _12727_/A _23692_/Q VGND VGND VPWR VPWR _12229_/X sky130_fd_sc_hd__or2_4
XFILLER_130_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15017_ _15017_/A _23957_/Q VGND VGND VPWR VPWR _15017_/X sky130_fd_sc_hd__or2_4
XFILLER_170_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23125__CLK _23456_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19825_ _19898_/B _19808_/A VGND VGND VPWR VPWR _19826_/C sky130_fd_sc_hd__or2_4
XFILLER_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20270__A _18889_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11892__A _11891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19756_ HRDATA[4] VGND VGND VPWR VPWR _19756_/Y sky130_fd_sc_hd__inv_2
X_16968_ _24138_/Q VGND VGND VPWR VPWR _17732_/A sky130_fd_sc_hd__inv_2
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18707_ _18624_/X _18705_/X _18706_/Y _11642_/X VGND VGND VPWR VPWR _18707_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__22545__B2 _22541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15919_ _15521_/X _15656_/X _16855_/A _15919_/D VGND VGND VPWR VPWR _15919_/X sky130_fd_sc_hd__or4_4
X_19687_ _19687_/A _19815_/B _19687_/C _19687_/D VGND VGND VPWR VPWR _19687_/X sky130_fd_sc_hd__and4_4
XANTENNA__12500__B _12500_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16899_ _16899_/A _16898_/X VGND VGND VPWR VPWR _16899_/Y sky130_fd_sc_hd__nand2_4
XFILLER_92_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18638_ _17111_/X _18091_/Y _17224_/X _18637_/X VGND VGND VPWR VPWR _18638_/X sky130_fd_sc_hd__a211o_4
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18569_ _18477_/X _18556_/Y _18504_/X _18568_/X VGND VGND VPWR VPWR _18569_/X sky130_fd_sc_hd__o22a_4
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14708__A _13791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20600_ _20847_/A VGND VGND VPWR VPWR _20652_/A sky130_fd_sc_hd__buf_2
XANTENNA__13612__A _11932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21580_ _20819_/A VGND VGND VPWR VPWR _21580_/X sky130_fd_sc_hd__buf_2
XFILLER_33_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22925__A _18681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20531_ _20531_/A VGND VGND VPWR VPWR _20531_/X sky130_fd_sc_hd__buf_2
XFILLER_137_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23250_ _23537_/CLK _22496_/X VGND VGND VPWR VPWR _16679_/B sky130_fd_sc_hd__dfxtp_4
X_20462_ _24237_/Q _20420_/X _20461_/X VGND VGND VPWR VPWR _22113_/A sky130_fd_sc_hd__o21a_4
X_22201_ _22194_/A VGND VGND VPWR VPWR _22201_/X sky130_fd_sc_hd__buf_2
X_23181_ _23533_/CLK _23181_/D VGND VGND VPWR VPWR _16193_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21284__B2 _21276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22481__B1 _15122_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20393_ _24240_/Q _20304_/X _20392_/Y VGND VGND VPWR VPWR _22420_/A sky130_fd_sc_hd__o21a_4
XANTENNA__14443__A _14304_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22132_ _20632_/A VGND VGND VPWR VPWR _22132_/X sky130_fd_sc_hd__buf_2
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14162__B _23647_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13059__A _13094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22063_ _21843_/X _22060_/X _23495_/Q _22057_/X VGND VGND VPWR VPWR _22063_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21036__B2 _21035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21014_ _20425_/A _21013_/X _19226_/B _20349_/A VGND VGND VPWR VPWR _21014_/X sky130_fd_sc_hd__o22a_4
XFILLER_47_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21276__A _21264_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12898__A _12871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15274__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21339__A2 _21334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22965_ _22964_/X VGND VGND VPWR VPWR HADDR[10] sky130_fd_sc_hd__inv_2
XFILLER_90_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21916_ _21909_/A VGND VGND VPWR VPWR _21916_/X sky130_fd_sc_hd__buf_2
XFILLER_16_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22896_ _16687_/A _22885_/X _19909_/X _22895_/X VGND VGND VPWR VPWR _22896_/X sky130_fd_sc_hd__o22a_4
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21847_ _21845_/X _21839_/X _13388_/B _21846_/X VGND VGND VPWR VPWR _23622_/D sky130_fd_sc_hd__o22a_4
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20339__B _20339_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _24210_/Q VGND VGND VPWR VPWR _18782_/B sky130_fd_sc_hd__buf_2
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12580_/A VGND VGND VPWR VPWR _12581_/A sky130_fd_sc_hd__buf_2
X_21778_ _21553_/X _21777_/X _12902_/B _21774_/X VGND VGND VPWR VPWR _23657_/D sky130_fd_sc_hd__o22a_4
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22835__A _22884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17715__B2 _17368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21511__A2 _21506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14337__B _14337_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _24357_/Q _11530_/X VGND VGND VPWR VPWR _11532_/B sky130_fd_sc_hd__or2_4
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20729_ _20493_/A VGND VGND VPWR VPWR _20730_/B sky130_fd_sc_hd__buf_2
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23517_ _23518_/CLK _23517_/D VGND VGND VPWR VPWR _13800_/B sky130_fd_sc_hd__dfxtp_4
X_24497_ _24158_/CLK _24497_/D HRESETn VGND VGND VPWR VPWR _19993_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _13865_/A _14246_/X _14249_/X VGND VGND VPWR VPWR _14250_/X sky130_fd_sc_hd__or3_4
X_23448_ _23290_/CLK _23448_/D VGND VGND VPWR VPWR _23448_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _13200_/X _23751_/Q VGND VGND VPWR VPWR _13202_/C sky130_fd_sc_hd__or2_4
XANTENNA__11977__A _16148_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15449__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14181_ _14225_/A _23263_/Q VGND VGND VPWR VPWR _14185_/B sky130_fd_sc_hd__or2_4
X_23379_ _23379_/CLK _22281_/X VGND VGND VPWR VPWR _12119_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_152_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14353__A _14390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13132_ _13276_/A _13130_/X _13131_/X VGND VGND VPWR VPWR _13133_/C sky130_fd_sc_hd__and3_4
XFILLER_152_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13063_ _13063_/A VGND VGND VPWR VPWR _13100_/A sky130_fd_sc_hd__buf_2
X_17940_ _17940_/A VGND VGND VPWR VPWR _17940_/Y sky130_fd_sc_hd__inv_2
X_12014_ _11960_/A _21655_/A VGND VGND VPWR VPWR _12016_/B sky130_fd_sc_hd__or2_4
XANTENNA__21186__A _21219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17871_ _17249_/X VGND VGND VPWR VPWR _18413_/A sky130_fd_sc_hd__buf_2
Xclkbuf_4_6_0_HCLK clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19610_ _19703_/A HRDATA[11] VGND VGND VPWR VPWR _19610_/X sky130_fd_sc_hd__and2_4
XFILLER_120_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17651__B1 _17014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16822_ _16822_/A VGND VGND VPWR VPWR _16822_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12601__A _12927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22527__B2 _22526_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19541_ _19480_/X _19540_/X HRDATA[5] _19484_/X VGND VGND VPWR VPWR _19888_/B sky130_fd_sc_hd__o22a_4
X_16753_ _16635_/A _16753_/B _16753_/C VGND VGND VPWR VPWR _16760_/B sky130_fd_sc_hd__and3_4
XFILLER_4_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13965_ _13965_/A _13965_/B _13965_/C VGND VGND VPWR VPWR _13965_/X sky130_fd_sc_hd__and3_4
XFILLER_98_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15704_ _13332_/A _15704_/B VGND VGND VPWR VPWR _15706_/B sky130_fd_sc_hd__or2_4
XANTENNA__15912__A _13566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12916_ _12923_/A _12916_/B VGND VGND VPWR VPWR _12916_/X sky130_fd_sc_hd__or2_4
X_19472_ _19465_/A VGND VGND VPWR VPWR _19806_/A sky130_fd_sc_hd__buf_2
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16684_ _16684_/A _16668_/X _16684_/C VGND VGND VPWR VPWR _16685_/C sky130_fd_sc_hd__or3_4
XFILLER_74_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17954__A1 _18411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13896_ _14386_/A _13896_/B VGND VGND VPWR VPWR _13896_/X sky130_fd_sc_hd__or2_4
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21750__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18423_ _18413_/X _17391_/X _18417_/X _18168_/X _18422_/Y VGND VGND VPWR VPWR _18424_/B
+ sky130_fd_sc_hd__a32o_4
X_15635_ _15642_/A _15574_/B VGND VGND VPWR VPWR _15635_/X sky130_fd_sc_hd__or2_4
X_12847_ _12847_/A _12915_/B VGND VGND VPWR VPWR _12847_/X sky130_fd_sc_hd__or2_4
XFILLER_61_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13432__A _13431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18354_ _18215_/X _18351_/X _18240_/X _18353_/X VGND VGND VPWR VPWR _18354_/X sky130_fd_sc_hd__o22a_4
X_15566_ _14420_/A _15566_/B VGND VGND VPWR VPWR _15566_/X sky130_fd_sc_hd__or2_4
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _13051_/A VGND VGND VPWR VPWR _12778_/X sky130_fd_sc_hd__buf_2
XFILLER_159_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21502__A2 _21499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22745__A _22745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14247__B _23711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17305_ _17289_/X _17301_/Y _17304_/X VGND VGND VPWR VPWR _17305_/X sky130_fd_sc_hd__a21o_4
X_14517_ _14517_/A _23963_/Q VGND VGND VPWR VPWR _14518_/C sky130_fd_sc_hd__or2_4
X_11729_ _16033_/A VGND VGND VPWR VPWR _16080_/A sky130_fd_sc_hd__buf_2
XANTENNA__15717__B1 _12264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18285_ _17976_/X _17941_/X _17882_/X VGND VGND VPWR VPWR _18285_/Y sky130_fd_sc_hd__o21ai_4
X_15497_ _15502_/A _15497_/B VGND VGND VPWR VPWR _15497_/X sky130_fd_sc_hd__or2_4
XANTENNA__16743__A _11943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17236_ _17825_/A _17236_/B VGND VGND VPWR VPWR _17236_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14448_ _14448_/A _14446_/X _14447_/X VGND VGND VPWR VPWR _14448_/X sky130_fd_sc_hd__and3_4
XANTENNA__20265__A _20264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11887__A _11887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15359__A _13704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17167_ _17160_/X _17163_/X _17838_/A _17166_/X VGND VGND VPWR VPWR _17167_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22463__B1 _23263_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14379_ _14540_/A _14376_/X _14378_/X VGND VGND VPWR VPWR _14379_/X sky130_fd_sc_hd__and3_4
XANTENNA__14263__A _14263_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16118_ _16147_/A _16203_/B VGND VGND VPWR VPWR _16119_/C sky130_fd_sc_hd__or2_4
XFILLER_142_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17098_ _18485_/A VGND VGND VPWR VPWR _18674_/A sky130_fd_sc_hd__buf_2
XFILLER_89_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21018__A1 _18774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17574__A _16162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16049_ _16049_/A _23566_/Q VGND VGND VPWR VPWR _16050_/C sky130_fd_sc_hd__or2_4
XANTENNA__21569__A2 _21566_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19808_ _19808_/A VGND VGND VPWR VPWR _19808_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13607__A _13607_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21189__A2_N _21188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22518__B2 _22512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19739_ _19732_/X _19735_/X _19738_/X _17820_/X _19719_/X VGND VGND VPWR VPWR _19739_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15822__A _12884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22750_ SYSTICKCLKDIV[7] VGND VGND VPWR VPWR _22750_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21701_ _21594_/X _21698_/X _15307_/B _21695_/X VGND VGND VPWR VPWR _23704_/D sky130_fd_sc_hd__o22a_4
XFILLER_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22681_ _22476_/X _22679_/X _14743_/B _22676_/X VGND VGND VPWR VPWR _22681_/X sky130_fd_sc_hd__o22a_4
XFILLER_164_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14438__A _12492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24420_ _23475_/CLK _24420_/D HRESETn VGND VGND VPWR VPWR _24420_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13342__A _13341_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21632_ _21560_/X _21627_/X _13280_/B _21631_/X VGND VGND VPWR VPWR _21632_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19698__A1 _17005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19698__B2 HRDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14157__B _24095_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24351_ _24382_/CLK _24351_/D HRESETn VGND VGND VPWR VPWR _19075_/A sky130_fd_sc_hd__dfstp_4
XFILLER_166_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21563_ _21848_/A VGND VGND VPWR VPWR _21563_/X sky130_fd_sc_hd__buf_2
XANTENNA__16653__A _16053_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23302_ _24102_/CLK _22381_/X VGND VGND VPWR VPWR _23302_/Q sky130_fd_sc_hd__dfxtp_4
X_20514_ _20261_/X VGND VGND VPWR VPWR _20514_/X sky130_fd_sc_hd__buf_2
XANTENNA__24416__CLK _23476_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24282_ _24292_/CLK _24282_/D HRESETn VGND VGND VPWR VPWR _19231_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15184__A1 _14302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21494_ _21271_/X _21492_/X _13110_/B _21489_/X VGND VGND VPWR VPWR _21494_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23233_ _23617_/CLK _23233_/D VGND VGND VPWR VPWR _15569_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_153_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20445_ _20444_/X _21007_/B _20308_/X VGND VGND VPWR VPWR _20445_/X sky130_fd_sc_hd__a21o_4
XANTENNA__19964__A _18407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14173__A _14012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23164_ _24096_/CLK _23164_/D VGND VGND VPWR VPWR _14362_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20376_ _24241_/Q _20304_/X _20375_/Y VGND VGND VPWR VPWR _20377_/A sky130_fd_sc_hd__o21a_4
XANTENNA__22390__A _22357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22115_ _20485_/A VGND VGND VPWR VPWR _22115_/X sky130_fd_sc_hd__buf_2
XFILLER_161_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23095_ _23095_/CLK _22733_/X VGND VGND VPWR VPWR _15176_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22757__A1 SYSTICKCLKDIV[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22046_ _22060_/A VGND VGND VPWR VPWR _22046_/X sky130_fd_sc_hd__buf_2
XFILLER_47_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13517__A _12971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12421__A _12320_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22509__A1 _22437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22509__B2 _22505_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21980__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21734__A _21727_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23997_ _23997_/CLK _23997_/D VGND VGND VPWR VPWR _23997_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15732__A _13100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13750_ _14541_/A _13750_/B VGND VGND VPWR VPWR _13750_/X sky130_fd_sc_hd__or2_4
X_22948_ _22922_/A VGND VGND VPWR VPWR _22949_/A sky130_fd_sc_hd__buf_2
XANTENNA__21732__A2 _21727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12701_ _13277_/A _23690_/Q VGND VGND VPWR VPWR _12704_/B sky130_fd_sc_hd__or2_4
XFILLER_43_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13681_ _15442_/A _13681_/B _13680_/X VGND VGND VPWR VPWR _13681_/X sky130_fd_sc_hd__or3_4
Xclkbuf_4_14_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22879_ _17574_/Y _22836_/X _22875_/X _22878_/X VGND VGND VPWR VPWR _22880_/B sky130_fd_sc_hd__o22a_4
XANTENNA__14348__A _14348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15420_ _15420_/A _15419_/X VGND VGND VPWR VPWR _15420_/X sky130_fd_sc_hd__and2_4
X_12632_ _12632_/A _12632_/B VGND VGND VPWR VPWR _12633_/C sky130_fd_sc_hd__or2_4
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22565__A _22558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12563_ _12904_/A _12563_/B _12562_/X VGND VGND VPWR VPWR _12563_/X sky130_fd_sc_hd__or3_4
X_15351_ _15326_/A _15351_/B VGND VGND VPWR VPWR _15351_/X sky130_fd_sc_hd__or2_4
XFILLER_157_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16563__A _12015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ _11514_/A VGND VGND VPWR VPWR _11516_/A sky130_fd_sc_hd__inv_2
X_14302_ _14302_/A _14301_/X VGND VGND VPWR VPWR _14302_/X sky130_fd_sc_hd__and2_4
X_18070_ _18070_/A _17009_/B VGND VGND VPWR VPWR _18070_/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15282_ _13586_/A _15259_/X _15266_/X _15273_/X _15281_/X VGND VGND VPWR VPWR _15282_/X
+ sky130_fd_sc_hd__a32o_4
X_12494_ _12188_/A VGND VGND VPWR VPWR _12495_/A sky130_fd_sc_hd__buf_2
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17021_ _17020_/X VGND VGND VPWR VPWR _17021_/X sky130_fd_sc_hd__buf_2
XANTENNA__21248__B2 _21240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15179__A _15000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14233_ _14630_/A _14228_/X _14232_/X VGND VGND VPWR VPWR _14243_/B sky130_fd_sc_hd__or3_4
XFILLER_172_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14083__A _15649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14164_ _14277_/A _14164_/B _14164_/C VGND VGND VPWR VPWR _14164_/X sky130_fd_sc_hd__or3_4
XANTENNA__21909__A _21909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13115_ _13091_/A _13115_/B _13114_/X VGND VGND VPWR VPWR _13123_/B sky130_fd_sc_hd__or3_4
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24136__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18972_ _24401_/Q VGND VGND VPWR VPWR _18972_/Y sky130_fd_sc_hd__inv_2
X_14095_ _12473_/A VGND VGND VPWR VPWR _14096_/A sky130_fd_sc_hd__buf_2
XANTENNA__14811__A _11674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22748__A1 _19920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13046_ _13046_/A _13045_/X VGND VGND VPWR VPWR _13046_/X sky130_fd_sc_hd__and2_4
X_17923_ _17922_/X _17148_/X _17815_/X _17158_/X VGND VGND VPWR VPWR _17923_/X sky130_fd_sc_hd__o22a_4
XFILLER_61_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13427__A _13427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17854_ _17854_/A VGND VGND VPWR VPWR _17854_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12331__A _13205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16805_ _16767_/A _16803_/X _16804_/X VGND VGND VPWR VPWR _16805_/X sky130_fd_sc_hd__and3_4
X_17785_ _17654_/X _17784_/X _17654_/X _17784_/X VGND VGND VPWR VPWR _17785_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14997_ _13953_/A _23285_/Q VGND VGND VPWR VPWR _14997_/X sky130_fd_sc_hd__or2_4
XFILLER_94_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16738__A _12064_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19524_ _19524_/A VGND VGND VPWR VPWR _19624_/B sky130_fd_sc_hd__buf_2
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16736_ _16732_/A _16736_/B _16736_/C VGND VGND VPWR VPWR _16740_/B sky130_fd_sc_hd__and3_4
X_13948_ _13863_/X _13946_/Y VGND VGND VPWR VPWR _13949_/A sky130_fd_sc_hd__or2_4
Xclkbuf_1_1_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_1_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21723__A2 _21720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19455_ _19452_/X VGND VGND VPWR VPWR _19455_/Y sky130_fd_sc_hd__inv_2
X_16667_ _16675_/A _16667_/B _16666_/X VGND VGND VPWR VPWR _16667_/X sky130_fd_sc_hd__or3_4
XANTENNA__14258__A _11680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13879_ _14375_/A _13876_/X _13879_/C VGND VGND VPWR VPWR _13879_/X sky130_fd_sc_hd__and3_4
XANTENNA__13162__A _13279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18406_ _18406_/A _18406_/B VGND VGND VPWR VPWR _18409_/B sky130_fd_sc_hd__and2_4
XANTENNA__23313__CLK _23761_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15618_ _11675_/A _15600_/X _15618_/C VGND VGND VPWR VPWR _15618_/X sky130_fd_sc_hd__or3_4
X_19386_ _19383_/X _23078_/B _19328_/Y _19385_/Y VGND VGND VPWR VPWR _19386_/X sky130_fd_sc_hd__o22a_4
X_16598_ _12001_/A _16598_/B _16597_/X VGND VGND VPWR VPWR _16599_/C sky130_fd_sc_hd__and3_4
XFILLER_148_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18337_ _18283_/A _18337_/B _18337_/C _18337_/D VGND VGND VPWR VPWR _18338_/A sky130_fd_sc_hd__or4_4
XANTENNA__21487__B2 _21482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17569__A _17139_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15549_ _12288_/A _15545_/X _15548_/X VGND VGND VPWR VPWR _15549_/X sky130_fd_sc_hd__or3_4
XFILLER_124_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24378__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18268_ _18198_/X _18264_/Y _18265_/X _18267_/Y VGND VGND VPWR VPWR _18268_/X sky130_fd_sc_hd__a211o_4
X_17219_ _17218_/X VGND VGND VPWR VPWR _17219_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_34_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_34_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18199_ _17833_/X _17180_/X _17877_/X _17218_/X VGND VGND VPWR VPWR _18199_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__12506__A _12506_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20230_ _20229_/X VGND VGND VPWR VPWR _20231_/A sky130_fd_sc_hd__buf_2
XFILLER_144_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15817__A _11970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20161_ _20161_/A VGND VGND VPWR VPWR _20161_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14721__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22739__B2 _23086_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20092_ _11586_/X VGND VGND VPWR VPWR _20124_/B sky130_fd_sc_hd__inv_2
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23920_ _24080_/CLK _21332_/X VGND VGND VPWR VPWR _16421_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21411__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12241__A _13164_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21962__A2 _21960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21554__A _21542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23851_ _24074_/CLK _21439_/X VGND VGND VPWR VPWR _12549_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16648__A _16672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22802_ _22799_/X _22801_/X VGND VGND VPWR VPWR _22802_/X sky130_fd_sc_hd__or2_4
X_23782_ _23397_/CLK _21562_/X VGND VGND VPWR VPWR _23782_/Q sky130_fd_sc_hd__dfxtp_4
X_20994_ _20782_/X _20993_/X _24342_/Q _20789_/X VGND VGND VPWR VPWR _20994_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21714__A2 _21713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22733_ _21311_/A _22729_/X _15176_/B _22698_/A VGND VGND VPWR VPWR _22733_/X sky130_fd_sc_hd__o22a_4
XFILLER_38_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13072__A _13100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18591__B2 _18590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22664_ _22447_/X _22658_/X _13462_/B _22662_/X VGND VGND VPWR VPWR _23141_/D sky130_fd_sc_hd__o22a_4
XFILLER_129_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21615_ _21532_/X _21613_/X _23762_/Q _21610_/X VGND VGND VPWR VPWR _21615_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_116_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR _23678_/CLK sky130_fd_sc_hd__clkbuf_1
X_24403_ _23409_/CLK _24403_/D HRESETn VGND VGND VPWR VPWR _24403_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22675__B1 _13838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23806__CLK _23101_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22595_ _22412_/X _22594_/X _12135_/B _22591_/X VGND VGND VPWR VPWR _23187_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19540__B1 HRDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20686__C1 _20685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13800__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21546_ _20486_/A VGND VGND VPWR VPWR _21546_/X sky130_fd_sc_hd__buf_2
X_24334_ _24294_/CLK _19174_/X HRESETn VGND VGND VPWR VPWR _19155_/A sky130_fd_sc_hd__dfrtp_4
X_24265_ _24495_/CLK _19351_/X HRESETn VGND VGND VPWR VPWR _24265_/Q sky130_fd_sc_hd__dfrtp_4
X_21477_ _21506_/A VGND VGND VPWR VPWR _21492_/A sky130_fd_sc_hd__buf_2
XANTENNA__12416__A _13564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22832__B _14767_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23216_ _23760_/CLK _23216_/D VGND VGND VPWR VPWR _16394_/B sky130_fd_sc_hd__dfxtp_4
X_20428_ _24430_/Q _20427_/X _24462_/Q _20282_/X VGND VGND VPWR VPWR _20428_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24196_ _24184_/CLK _19805_/X HRESETn VGND VGND VPWR VPWR _11653_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23147_ _24012_/CLK _22656_/X VGND VGND VPWR VPWR _12548_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15727__A _12762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20359_ _24242_/Q _20304_/X _20358_/Y VGND VGND VPWR VPWR _20360_/A sky130_fd_sc_hd__o21a_4
XANTENNA__21650__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23078_ _23078_/A _23078_/B VGND VGND VPWR VPWR _23078_/X sky130_fd_sc_hd__or2_4
XFILLER_0_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13247__A _13235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14920_ _14916_/X _14918_/X _14920_/C VGND VGND VPWR VPWR _14920_/X sky130_fd_sc_hd__and3_4
XFILLER_96_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22029_ _21869_/X _22024_/X _14339_/B _22028_/X VGND VGND VPWR VPWR _23516_/D sky130_fd_sc_hd__o22a_4
XFILLER_130_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14851_ _11618_/A _14849_/X _14850_/X VGND VGND VPWR VPWR _14851_/X sky130_fd_sc_hd__and3_4
XFILLER_21_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11990__A _11990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19359__B1 _19358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23336__CLK _23592_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13802_ _13617_/A VGND VGND VPWR VPWR _14307_/A sky130_fd_sc_hd__buf_2
X_17570_ _16085_/X _18076_/B VGND VGND VPWR VPWR _17571_/A sky130_fd_sc_hd__or2_4
X_14782_ _15106_/A _14778_/X _14782_/C VGND VGND VPWR VPWR _14782_/X sky130_fd_sc_hd__or3_4
X_11994_ _11990_/A _23860_/Q VGND VGND VPWR VPWR _11995_/C sky130_fd_sc_hd__or2_4
XANTENNA__22902__A1 _12021_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16521_ _13417_/A _16489_/X _16520_/X VGND VGND VPWR VPWR _16521_/X sky130_fd_sc_hd__and3_4
X_13733_ _13742_/A _13733_/B VGND VGND VPWR VPWR _13734_/C sky130_fd_sc_hd__or2_4
XANTENNA__14078__A _12322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19240_ _19240_/A _19240_/B VGND VGND VPWR VPWR _19240_/X sky130_fd_sc_hd__and2_4
XFILLER_56_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16452_ _16451_/X VGND VGND VPWR VPWR _16452_/Y sky130_fd_sc_hd__inv_2
X_13664_ _14331_/A VGND VGND VPWR VPWR _15412_/A sky130_fd_sc_hd__buf_2
XFILLER_32_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15403_ _13656_/A _15466_/B VGND VGND VPWR VPWR _15403_/X sky130_fd_sc_hd__or2_4
X_12615_ _11781_/A VGND VGND VPWR VPWR _12616_/A sky130_fd_sc_hd__buf_2
X_19171_ _19157_/B VGND VGND VPWR VPWR _19171_/Y sky130_fd_sc_hd__inv_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17389__A _17360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16383_ _16383_/A VGND VGND VPWR VPWR _16383_/X sky130_fd_sc_hd__buf_2
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ _13983_/A VGND VGND VPWR VPWR _13596_/A sky130_fd_sc_hd__buf_2
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19531__B1 HRDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18122_ _18122_/A VGND VGND VPWR VPWR _18122_/Y sky130_fd_sc_hd__inv_2
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15334_ _15372_/A _15334_/B _15333_/X VGND VGND VPWR VPWR _15338_/B sky130_fd_sc_hd__and3_4
X_12546_ _12546_/A VGND VGND VPWR VPWR _12911_/A sky130_fd_sc_hd__buf_2
XFILLER_61_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18053_ _17245_/X VGND VGND VPWR VPWR _18053_/X sky130_fd_sc_hd__buf_2
XFILLER_145_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15265_ _12426_/A _15263_/X _15264_/X VGND VGND VPWR VPWR _15266_/C sky130_fd_sc_hd__and3_4
X_12477_ _12477_/A VGND VGND VPWR VPWR _12537_/A sky130_fd_sc_hd__buf_2
XFILLER_144_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17004_ _18576_/B VGND VGND VPWR VPWR _17005_/A sky130_fd_sc_hd__inv_2
XANTENNA__18098__B1 _17919_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14216_ _14240_/A _23999_/Q VGND VGND VPWR VPWR _14217_/C sky130_fd_sc_hd__or2_4
XFILLER_160_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15196_ _14229_/A VGND VGND VPWR VPWR _15196_/X sky130_fd_sc_hd__buf_2
XFILLER_126_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14147_ _12433_/A _23391_/Q VGND VGND VPWR VPWR _14149_/B sky130_fd_sc_hd__or2_4
XANTENNA__15637__A _13884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18955_ _18955_/A VGND VGND VPWR VPWR _18955_/Y sky130_fd_sc_hd__inv_2
X_14078_ _12322_/A _23232_/Q VGND VGND VPWR VPWR _14080_/B sky130_fd_sc_hd__or2_4
XANTENNA__22197__A2 _22194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13029_ _12513_/A _13105_/B VGND VGND VPWR VPWR _13029_/X sky130_fd_sc_hd__or2_4
X_17906_ _17906_/A _17906_/B _17906_/C _16996_/B VGND VGND VPWR VPWR _17964_/B sky130_fd_sc_hd__or4_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18886_ _17251_/A _17398_/A _17037_/Y _17427_/A VGND VGND VPWR VPWR _18889_/B sky130_fd_sc_hd__or4_4
XANTENNA__12061__A _12061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21374__A _21381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17837_ _17160_/X VGND VGND VPWR VPWR _17837_/X sky130_fd_sc_hd__buf_2
XFILLER_67_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12996__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15372__A _15372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24261__CLK _24127_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17768_ _17711_/A _17768_/B _17768_/C VGND VGND VPWR VPWR _17768_/X sky130_fd_sc_hd__and3_4
XFILLER_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19507_ _19507_/A _19507_/B VGND VGND VPWR VPWR _19508_/A sky130_fd_sc_hd__or2_4
X_16719_ _12028_/X _16696_/X _16703_/X _16710_/X _16718_/X VGND VGND VPWR VPWR _16719_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23829__CLK _23456_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17699_ _17699_/A VGND VGND VPWR VPWR _17699_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19770__B1 _20561_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19438_ _19438_/A _19438_/B VGND VGND VPWR VPWR _19439_/A sky130_fd_sc_hd__or2_4
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20718__A _20718_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19369_ _19372_/A VGND VGND VPWR VPWR _19369_/X sky130_fd_sc_hd__buf_2
XANTENNA__14716__A _14325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21400_ _21283_/X _21398_/X _15844_/B _21395_/X VGND VGND VPWR VPWR _21400_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22121__A2 _22111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13620__A _15401_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22380_ _22358_/A VGND VGND VPWR VPWR _22380_/X sky130_fd_sc_hd__buf_2
XANTENNA__22933__A _22945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21331_ _21331_/A VGND VGND VPWR VPWR _21331_/X sky130_fd_sc_hd__buf_2
XFILLER_50_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12236__A _12236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21880__B2 _21870_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24050_ _23922_/CLK _24050_/D VGND VGND VPWR VPWR _24050_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21549__A _21549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21262_ _21261_/X _21257_/X _12357_/B _21252_/X VGND VGND VPWR VPWR _23948_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23209__CLK _23561_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23001_ _23043_/A _23001_/B VGND VGND VPWR VPWR _23001_/Y sky130_fd_sc_hd__nand2_4
XFILLER_116_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20213_ _22039_/A _22039_/B VGND VGND VPWR VPWR _21234_/A sky130_fd_sc_hd__or2_4
XANTENNA__15547__A _14421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21632__B2 _21631_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21193_ _20361_/X _21191_/X _23986_/Q _21188_/X VGND VGND VPWR VPWR _23986_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17465__A1_N _12753_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20144_ _20132_/Y _20143_/Y _20125_/X _20192_/A VGND VGND VPWR VPWR _20145_/A sky130_fd_sc_hd__a211o_4
XANTENNA__22188__A2 _22187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13067__A _13067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20075_ _24480_/Q VGND VGND VPWR VPWR _20075_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21396__B1 _13405_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21935__A2 _21930_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17064__B2 _17251_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23903_ _23518_/CLK _23903_/D VGND VGND VPWR VPWR _23903_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17481__B _17481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16378__A _11684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23834_ _23294_/CLK _23834_/D VGND VGND VPWR VPWR _14591_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21699__A1 _21589_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _20977_/A _20976_/X VGND VGND VPWR VPWR _20977_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21699__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23765_ _23904_/CLK _23765_/D VGND VGND VPWR VPWR _23765_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17367__A2 _17378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22716_ _21280_/A _22715_/X _23108_/Q _22712_/X VGND VGND VPWR VPWR _23108_/D sky130_fd_sc_hd__o22a_4
XFILLER_14_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23696_ _24080_/CLK _21718_/X VGND VGND VPWR VPWR _16403_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_80_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22647_ _22418_/X _22644_/X _16795_/B _22641_/X VGND VGND VPWR VPWR _23153_/D sky130_fd_sc_hd__o22a_4
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14626__A _14669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22112__A2 _22111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19513__B1 _17037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13530__A _13530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12400_ _12387_/A _12398_/X _12400_/C VGND VGND VPWR VPWR _12400_/X sky130_fd_sc_hd__and3_4
X_13380_ _13398_/A _13378_/X _13380_/C VGND VGND VPWR VPWR _13381_/C sky130_fd_sc_hd__and3_4
XFILLER_167_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17002__A _24212_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24481__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22578_ _22471_/X _22572_/X _14491_/B _22576_/X VGND VGND VPWR VPWR _22578_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24361__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12331_ _13205_/A VGND VGND VPWR VPWR _12829_/A sky130_fd_sc_hd__buf_2
XANTENNA__21871__A1 _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24317_ _24287_/CLK _24317_/D HRESETn VGND VGND VPWR VPWR _24317_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21871__B2 _21870_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21529_ _21523_/A VGND VGND VPWR VPWR _21542_/A sky130_fd_sc_hd__buf_2
XFILLER_166_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12262_ _13016_/A _12261_/X VGND VGND VPWR VPWR _12262_/X sky130_fd_sc_hd__and2_4
X_15050_ _12322_/A _23253_/Q VGND VGND VPWR VPWR _15050_/X sky130_fd_sc_hd__or2_4
XANTENNA__21459__A _21438_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24248_ _24248_/CLK _19375_/X HRESETn VGND VGND VPWR VPWR _24248_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20363__A _18779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24134__CLK _24134_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14001_ _11623_/A _23232_/Q VGND VGND VPWR VPWR _14003_/B sky130_fd_sc_hd__or2_4
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15457__A _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11985__A _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21623__B2 _21617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12193_ _12568_/A _12193_/B VGND VGND VPWR VPWR _12201_/B sky130_fd_sc_hd__or2_4
X_24179_ _23383_/CLK _24179_/D HRESETn VGND VGND VPWR VPWR _24179_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14361__A _14512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15176__B _15176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18740_ _16943_/A _18727_/X _18504_/X _22846_/B VGND VGND VPWR VPWR _18740_/X sky130_fd_sc_hd__o22a_4
X_15952_ _15952_/A _15952_/B _15952_/C VGND VGND VPWR VPWR _15952_/X sky130_fd_sc_hd__and3_4
XFILLER_110_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24284__CLK _24292_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21387__B1 _12314_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21926__A2 _21923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14903_ _14155_/A _14967_/B VGND VGND VPWR VPWR _14903_/X sky130_fd_sc_hd__or2_4
X_18671_ _17756_/X _17747_/X _17756_/X _17747_/X VGND VGND VPWR VPWR _18671_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17391__B _17448_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15883_ _12402_/X _15883_/B _15883_/C VGND VGND VPWR VPWR _15883_/X sky130_fd_sc_hd__and3_4
XFILLER_48_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17622_ _17324_/X VGND VGND VPWR VPWR _18693_/B sky130_fd_sc_hd__inv_2
XFILLER_56_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14834_ _14834_/A _14834_/B VGND VGND VPWR VPWR _14836_/B sky130_fd_sc_hd__or2_4
XANTENNA__13705__A _13705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17553_ _17120_/Y _17551_/B VGND VGND VPWR VPWR _17554_/B sky130_fd_sc_hd__and2_4
X_14765_ _15420_/A _14742_/X _14749_/X _14756_/X _14764_/X VGND VGND VPWR VPWR _14765_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11977_ _16148_/A _11977_/B _11977_/C VGND VGND VPWR VPWR _11977_/X sky130_fd_sc_hd__and3_4
XANTENNA__18555__A1 _18111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16504_ _11784_/X _16504_/B _16504_/C VGND VGND VPWR VPWR _16504_/X sky130_fd_sc_hd__and3_4
XANTENNA__22737__B _18576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13716_ _12596_/A VGND VGND VPWR VPWR _13756_/A sky130_fd_sc_hd__buf_2
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20362__A1 _20302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17484_ _17480_/Y _17022_/X _17029_/X _17483_/Y VGND VGND VPWR VPWR _17487_/B sky130_fd_sc_hd__o22a_4
XANTENNA__20362__B2 _20225_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14696_ _14647_/X _14696_/B _14696_/C VGND VGND VPWR VPWR _14696_/X sky130_fd_sc_hd__and3_4
XANTENNA__20538__A _20233_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19223_ _19223_/A VGND VGND VPWR VPWR _22945_/A sky130_fd_sc_hd__buf_2
X_16435_ _16112_/A _16435_/B VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__or2_4
X_13647_ _15444_/A _13738_/B VGND VGND VPWR VPWR _13648_/C sky130_fd_sc_hd__or2_4
XFILLER_158_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13440__A _12871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19154_ _19154_/A _19154_/B VGND VGND VPWR VPWR _19155_/B sky130_fd_sc_hd__and2_4
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16366_ _11715_/A _16303_/B VGND VGND VPWR VPWR _16366_/X sky130_fd_sc_hd__or2_4
XFILLER_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20114__A1 _20098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _12684_/X _13578_/B VGND VGND VPWR VPWR _13578_/Y sky130_fd_sc_hd__nor2_4
XFILLER_160_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14255__B _23647_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18105_ _18020_/X _18102_/X _18065_/X _18104_/X VGND VGND VPWR VPWR _18105_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15317_ _11654_/A _15317_/B _15317_/C VGND VGND VPWR VPWR _15317_/X sky130_fd_sc_hd__and3_4
X_19085_ _19074_/X _19083_/Y _19084_/Y _19079_/X VGND VGND VPWR VPWR _19085_/X sky130_fd_sc_hd__o22a_4
X_12529_ _14295_/A VGND VGND VPWR VPWR _12530_/A sky130_fd_sc_hd__buf_2
X_16297_ _15982_/A _16297_/B VGND VGND VPWR VPWR _16297_/X sky130_fd_sc_hd__or2_4
XANTENNA__12056__A _11943_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18036_ _17088_/A VGND VGND VPWR VPWR _18376_/A sky130_fd_sc_hd__buf_2
XANTENNA__23064__B1 _17957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15248_ _14614_/A _15240_/X _15248_/C VGND VGND VPWR VPWR _15248_/X sky130_fd_sc_hd__and3_4
XFILLER_132_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11895__A _12194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17818__B1 _17817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21614__B2 _21610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15367__A _12580_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15179_ _15000_/A _15179_/B VGND VGND VPWR VPWR _15181_/B sky130_fd_sc_hd__or2_4
XANTENNA__14271__A _12427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15086__B _23957_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19987_ _19987_/A VGND VGND VPWR VPWR _19987_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18938_ _14844_/X _18934_/X _24377_/Q _18935_/X VGND VGND VPWR VPWR _24377_/D sky130_fd_sc_hd__o22a_4
.ends

