* NGSPICE file created from NfiVe32_SYS.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

.subckt NfiVe32_SYS HADDR[0] HADDR[10] HADDR[11] HADDR[12] HADDR[13] HADDR[14] HADDR[15]
+ HADDR[16] HADDR[17] HADDR[18] HADDR[19] HADDR[1] HADDR[20] HADDR[21] HADDR[22] HADDR[23]
+ HADDR[24] HADDR[25] HADDR[26] HADDR[27] HADDR[28] HADDR[29] HADDR[2] HADDR[30] HADDR[31]
+ HADDR[3] HADDR[4] HADDR[5] HADDR[6] HADDR[7] HADDR[8] HADDR[9] HCLK HRDATA[0] HRDATA[10]
+ HRDATA[11] HRDATA[12] HRDATA[13] HRDATA[14] HRDATA[15] HRDATA[16] HRDATA[17] HRDATA[18]
+ HRDATA[19] HRDATA[1] HRDATA[20] HRDATA[21] HRDATA[22] HRDATA[23] HRDATA[24] HRDATA[25]
+ HRDATA[26] HRDATA[27] HRDATA[28] HRDATA[29] HRDATA[2] HRDATA[30] HRDATA[31] HRDATA[3]
+ HRDATA[4] HRDATA[5] HRDATA[6] HRDATA[7] HRDATA[8] HRDATA[9] HREADY HRESETn HSIZE[0]
+ HSIZE[1] HSIZE[2] HTRANS[0] HTRANS[1] HWDATA[0] HWDATA[10] HWDATA[11] HWDATA[12]
+ HWDATA[13] HWDATA[14] HWDATA[15] HWDATA[16] HWDATA[17] HWDATA[18] HWDATA[19] HWDATA[1]
+ HWDATA[20] HWDATA[21] HWDATA[22] HWDATA[23] HWDATA[24] HWDATA[25] HWDATA[26] HWDATA[27]
+ HWDATA[28] HWDATA[29] HWDATA[2] HWDATA[30] HWDATA[31] HWDATA[3] HWDATA[4] HWDATA[5]
+ HWDATA[6] HWDATA[7] HWDATA[8] HWDATA[9] HWRITE IRQ[0] IRQ[10] IRQ[11] IRQ[12] IRQ[13]
+ IRQ[14] IRQ[15] IRQ[16] IRQ[17] IRQ[18] IRQ[19] IRQ[1] IRQ[20] IRQ[21] IRQ[22] IRQ[23]
+ IRQ[24] IRQ[25] IRQ[26] IRQ[27] IRQ[28] IRQ[29] IRQ[2] IRQ[30] IRQ[31] IRQ[3] IRQ[4]
+ IRQ[5] IRQ[6] IRQ[7] IRQ[8] IRQ[9] NMI SYSTICKCLKDIV[0] SYSTICKCLKDIV[1] SYSTICKCLKDIV[2]
+ SYSTICKCLKDIV[3] SYSTICKCLKDIV[4] SYSTICKCLKDIV[5] SYSTICKCLKDIV[6] SYSTICKCLKDIV[7]
+ VPWR VGND
XANTENNA__21378__B1 _15839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15814__B _23885_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18869_ _20425_/A VGND VGND VPWR VPWR _20407_/A sky130_fd_sc_hd__buf_2
XFILLER_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18794__A1 _15646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16198__A _16198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20900_ _24387_/Q _20556_/A VGND VGND VPWR VPWR _20900_/Y sky130_fd_sc_hd__nand2_4
XFILLER_94_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13615__A _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21880_ _21887_/A VGND VGND VPWR VPWR _21880_/X sky130_fd_sc_hd__buf_2
XANTENNA__22928__A _18570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20831_ _20825_/X _20831_/B VGND VGND VPWR VPWR _20831_/Y sky130_fd_sc_hd__nor2_4
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15830__A _12522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20762_ _20762_/A VGND VGND VPWR VPWR _20762_/Y sky130_fd_sc_hd__inv_2
X_23550_ _23320_/CLK _23550_/D VGND VGND VPWR VPWR _23550_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19302__A _19317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20448__A _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22501_ _22439_/X _22500_/X _23209_/Q _22497_/X VGND VGND VPWR VPWR _22501_/X sky130_fd_sc_hd__o22a_4
XFILLER_74_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23481_ _23514_/CLK _23481_/D VGND VGND VPWR VPWR _23481_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20693_ _20673_/X _20679_/Y _20690_/X _20691_/Y _20692_/X VGND VGND VPWR VPWR _20693_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_5_13_0_HCLK_A clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22432_ _20696_/A VGND VGND VPWR VPWR _22432_/X sky130_fd_sc_hd__buf_2
XANTENNA__13350__A _13349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24157__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22363_ _22115_/X _22361_/X _15795_/B _22358_/X VGND VGND VPWR VPWR _23277_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16661__A _16624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21314_ _21237_/X _21312_/X _16124_/B _21309_/X VGND VGND VPWR VPWR _23895_/D sky130_fd_sc_hd__o22a_4
X_24102_ _24321_/CLK _24102_/D HRESETn VGND VGND VPWR VPWR _22741_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22294_ _22136_/X _22293_/X _14652_/B _22290_/X VGND VGND VPWR VPWR _23332_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16380__B _16380_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24033_ _23145_/CLK _21055_/X VGND VGND VPWR VPWR _15159_/B sky130_fd_sc_hd__dfxtp_4
X_21245_ _21244_/X _21235_/X _23924_/Q _21242_/X VGND VGND VPWR VPWR _23924_/D sky130_fd_sc_hd__o22a_4
XFILLER_2_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15277__A _15023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19972__A _19996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23181__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14181__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21176_ _21183_/A VGND VGND VPWR VPWR _21176_/X sky130_fd_sc_hd__buf_2
XFILLER_46_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20127_ _18603_/Y _18688_/X _20126_/X VGND VGND VPWR VPWR _20128_/B sky130_fd_sc_hd__o21a_4
XFILLER_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17492__A _17194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17037__A1 _18864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20058_ _20058_/A VGND VGND VPWR VPWR _20058_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22030__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15724__B _15724_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18785__A1 _13274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11900_ _15956_/A VGND VGND VPWR VPWR _15952_/A sky130_fd_sc_hd__buf_2
XANTENNA__13525__A _12981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22581__A2 _22579_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12880_ _12880_/A VGND VGND VPWR VPWR _13951_/A sky130_fd_sc_hd__buf_2
XFILLER_6_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11831_ _11821_/A _12014_/B VGND VGND VPWR VPWR _11831_/X sky130_fd_sc_hd__or2_4
X_23817_ _23910_/CLK _23817_/D VGND VGND VPWR VPWR _23817_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15740__A _12777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14550_ _13695_/X _14486_/B VGND VGND VPWR VPWR _14550_/X sky130_fd_sc_hd__or2_4
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11747_/X _11751_/X _11761_/X VGND VGND VPWR VPWR _11763_/C sky130_fd_sc_hd__or3_4
X_23748_ _23363_/CLK _23748_/D VGND VGND VPWR VPWR _14662_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_42_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20358__A _20342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _12965_/A VGND VGND VPWR VPWR _15879_/A sky130_fd_sc_hd__buf_2
XFILLER_14_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _12465_/A _14479_/X _14481_/C VGND VGND VPWR VPWR _14482_/C sky130_fd_sc_hd__and3_4
X_11693_ _11644_/A VGND VGND VPWR VPWR _14178_/A sky130_fd_sc_hd__buf_2
X_23679_ _23217_/CLK _23679_/D VGND VGND VPWR VPWR _23679_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16227_/A _16220_/B VGND VGND VPWR VPWR _16220_/X sky130_fd_sc_hd__or2_4
XANTENNA__13260__A _13260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _11913_/X _13430_/X _13431_/X VGND VGND VPWR VPWR _13433_/C sky130_fd_sc_hd__and3_4
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22097__B2 _22096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19866__B _19866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14075__B _14073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16151_ _16151_/A _16149_/X _16150_/X VGND VGND VPWR VPWR _16151_/X sky130_fd_sc_hd__and3_4
XANTENNA__19368__A2_N _17775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21844__A1 _21843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13363_ _11681_/X _13356_/X _13363_/C VGND VGND VPWR VPWR _13363_/X sky130_fd_sc_hd__or3_4
XFILLER_42_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17667__A _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22256__A2_N _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21844__B2 _21836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23524__CLK _23107_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15102_ _15069_/A _23071_/Q VGND VGND VPWR VPWR _15102_/X sky130_fd_sc_hd__or2_4
X_12314_ _15553_/A VGND VGND VPWR VPWR _12315_/A sky130_fd_sc_hd__buf_2
X_16082_ _13442_/X VGND VGND VPWR VPWR _16083_/A sky130_fd_sc_hd__buf_2
X_13294_ _13286_/X _24016_/Q VGND VGND VPWR VPWR _13294_/X sky130_fd_sc_hd__or2_4
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16290__B _16368_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15033_ _13925_/A _15033_/B VGND VGND VPWR VPWR _15035_/B sky130_fd_sc_hd__or2_4
X_19910_ _22723_/A VGND VGND VPWR VPWR _19910_/X sky130_fd_sc_hd__buf_2
X_12245_ _12235_/A VGND VGND VPWR VPWR _12725_/A sky130_fd_sc_hd__buf_2
XFILLER_29_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12176_ _11773_/X _12174_/X _12175_/X VGND VGND VPWR VPWR _12176_/X sky130_fd_sc_hd__and3_4
X_19841_ _19841_/A VGND VGND VPWR VPWR _21297_/A sky130_fd_sc_hd__buf_2
XFILLER_29_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13419__B _13336_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12323__B _12323_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20821__A HRDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18498__A _18498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16984_ _17661_/A _16983_/X VGND VGND VPWR VPWR _16984_/X sky130_fd_sc_hd__or2_4
X_19772_ _19873_/B _19592_/A _19640_/X VGND VGND VPWR VPWR _19772_/X sky130_fd_sc_hd__o21a_4
XFILLER_96_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13837__A1 _13594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15935_ _15934_/X _23512_/Q VGND VGND VPWR VPWR _15935_/X sky130_fd_sc_hd__or2_4
X_18723_ _17738_/X _17739_/X _17738_/X _17739_/X VGND VGND VPWR VPWR _18723_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_24_0_HCLK clkbuf_7_25_0_HCLK/A VGND VGND VPWR VPWR _24032_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18776__A1 _16374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13435__A _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18654_ _17742_/X _17743_/B _17742_/X _17743_/B VGND VGND VPWR VPWR _18654_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15866_ _13507_/X _15862_/X _15866_/C VGND VGND VPWR VPWR _15866_/X sky130_fd_sc_hd__or3_4
Xclkbuf_7_87_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR _23326_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21780__B1 _23617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14817_ _11766_/A _14817_/B _14817_/C VGND VGND VPWR VPWR _14818_/C sky130_fd_sc_hd__and3_4
X_17605_ _17605_/A VGND VGND VPWR VPWR _18621_/B sky130_fd_sc_hd__inv_2
XANTENNA__21652__A _21659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13154__B _23985_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18585_ _17618_/C _18585_/B VGND VGND VPWR VPWR _18585_/Y sky130_fd_sc_hd__nand2_4
X_15797_ _15820_/A _15793_/X _15797_/C VGND VGND VPWR VPWR _15797_/X sky130_fd_sc_hd__or3_4
XFILLER_17_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16746__A _11782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17536_ _16444_/Y _17016_/X _17023_/X _17535_/Y VGND VGND VPWR VPWR _17570_/A sky130_fd_sc_hd__o22a_4
XFILLER_83_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14748_ _14748_/A _14748_/B _14747_/X VGND VGND VPWR VPWR _14748_/X sky130_fd_sc_hd__and3_4
XANTENNA__16465__B _16405_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17467_ _11924_/A _17467_/B VGND VGND VPWR VPWR _17467_/X sky130_fd_sc_hd__and2_4
XFILLER_60_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14679_ _14679_/A _14679_/B VGND VGND VPWR VPWR _14679_/X sky130_fd_sc_hd__or2_4
XFILLER_60_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17751__A2 _17346_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16418_ _16083_/A _16416_/X _16418_/C VGND VGND VPWR VPWR _16418_/X sky130_fd_sc_hd__and3_4
X_19206_ _24257_/Q _19206_/B VGND VGND VPWR VPWR _19207_/B sky130_fd_sc_hd__and2_4
XFILLER_53_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17398_ _17395_/X _17397_/X VGND VGND VPWR VPWR _17603_/B sky130_fd_sc_hd__and2_4
XFILLER_14_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22483__A _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19137_ _19137_/A _19136_/X VGND VGND VPWR VPWR _19137_/X sky130_fd_sc_hd__and2_4
X_16349_ _16303_/X _16347_/X _16348_/X VGND VGND VPWR VPWR _16349_/X sky130_fd_sc_hd__and3_4
XFILLER_9_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16481__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19068_ _19068_/A VGND VGND VPWR VPWR _19068_/Y sky130_fd_sc_hd__inv_2
X_18019_ _18011_/X _17894_/X _18014_/Y _18016_/X _18018_/X VGND VGND VPWR VPWR _18019_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12514__A _13014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21030_ _21030_/A VGND VGND VPWR VPWR _21030_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22260__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21403__A2_N _21402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15825__A _12520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20810__A2 _20809_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17743__C _17742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22012__B2 _22006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15544__B _23563_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22981_ _18334_/X _23004_/B VGND VGND VPWR VPWR _22981_/X sky130_fd_sc_hd__or2_4
XFILLER_68_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22563__A2 _22536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13345__A _12859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21932_ _21804_/X _21931_/X _23544_/Q _21928_/X VGND VGND VPWR VPWR _21932_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21863_ _21293_/A VGND VGND VPWR VPWR _21863_/X sky130_fd_sc_hd__buf_2
XFILLER_83_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16656__A _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23602_ _23986_/CLK _21820_/X VGND VGND VPWR VPWR _23602_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15560__A _15533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20814_ _20616_/X _20802_/X _20757_/X _20813_/Y VGND VGND VPWR VPWR _20814_/X sky130_fd_sc_hd__a211o_4
XFILLER_58_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21794_ _21791_/X _21793_/X _23613_/Q _21788_/X VGND VGND VPWR VPWR _23613_/D sky130_fd_sc_hd__o22a_4
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20178__A _19313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23533_ _23922_/CLK _21947_/X VGND VGND VPWR VPWR _15802_/B sky130_fd_sc_hd__dfxtp_4
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20745_ _20634_/A _20744_/X VGND VGND VPWR VPWR _20745_/Y sky130_fd_sc_hd__nand2_4
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14176__A _11638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17742__A2 _17111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20676_ HRDATA[13] _20675_/X VGND VGND VPWR VPWR _20676_/X sky130_fd_sc_hd__or2_4
X_23464_ _23304_/CLK _23464_/D VGND VGND VPWR VPWR _23464_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22415_ _22100_/A VGND VGND VPWR VPWR _22415_/X sky130_fd_sc_hd__buf_2
XANTENNA__20629__A2 _20628_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23395_ _23270_/CLK _22195_/X VGND VGND VPWR VPWR _14766_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16391__A _16002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14904__A _14998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22346_ _22086_/X _22340_/X _16253_/B _22344_/X VGND VGND VPWR VPWR _22346_/X sky130_fd_sc_hd__o22a_4
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23697__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22277_ _22107_/X _22272_/X _13287_/B _22276_/X VGND VGND VPWR VPWR _23344_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12424__A _12386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12030_ _12029_/X VGND VGND VPWR VPWR _12031_/B sky130_fd_sc_hd__inv_2
XFILLER_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21228_ _21227_/X _21223_/X _23931_/Q _21218_/X VGND VGND VPWR VPWR _21228_/X sky130_fd_sc_hd__o22a_4
X_24016_ _23983_/CLK _21087_/X VGND VGND VPWR VPWR _24016_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21054__A2 _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21737__A _21752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13239__B _23953_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12143__B _23677_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11542__A2 IRQ[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15735__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21159_ _20982_/X _21154_/X _14873_/B _21115_/X VGND VGND VPWR VPWR _21159_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17739__A2_N _17122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22003__B2 _21999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15454__B _15454_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13981_ _12472_/A _23786_/Q VGND VGND VPWR VPWR _13982_/C sky130_fd_sc_hd__or2_4
XANTENNA__14492__A1 _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14492__B2 _14491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15720_ _13101_/A _15716_/X _15719_/X VGND VGND VPWR VPWR _15720_/X sky130_fd_sc_hd__or3_4
XANTENNA__13255__A _13243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12932_ _12958_/A _12857_/B VGND VGND VPWR VPWR _12932_/X sky130_fd_sc_hd__or2_4
XANTENNA__17950__A _18171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18222__A3 _18215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22568__A _22583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15651_ _15582_/X _15648_/X _15650_/Y VGND VGND VPWR VPWR _15914_/B sky130_fd_sc_hd__a21o_4
X_12863_ _12890_/A VGND VGND VPWR VPWR _12870_/A sky130_fd_sc_hd__buf_2
XFILLER_46_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16566__A _12011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19707__B1 _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14602_ _15030_/A _14676_/B VGND VGND VPWR VPWR _14602_/X sky130_fd_sc_hd__or2_4
X_11814_ _11819_/A _11814_/B VGND VGND VPWR VPWR _11814_/X sky130_fd_sc_hd__or2_4
X_18370_ _17874_/A _18392_/B VGND VGND VPWR VPWR _18370_/Y sky130_fd_sc_hd__nor2_4
X_15582_ _11842_/A _13595_/X _15551_/X _11596_/A _15581_/X VGND VGND VPWR VPWR _15582_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_76_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12794_ _12794_/A VGND VGND VPWR VPWR _12795_/A sky130_fd_sc_hd__buf_2
XANTENNA__20088__A _20071_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _18662_/A VGND VGND VPWR VPWR _17321_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14533_ _14533_/A _14533_/B VGND VGND VPWR VPWR _14534_/C sky130_fd_sc_hd__or2_4
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _16229_/A VGND VGND VPWR VPWR _11745_/X sky130_fd_sc_hd__buf_2
XANTENNA__19877__A _19877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17733__A2 _17106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18781__A _18781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17249_/A _17811_/A VGND VGND VPWR VPWR _17252_/X sky130_fd_sc_hd__or2_4
X_14464_ _14464_/A _14462_/X _14464_/C VGND VGND VPWR VPWR _14464_/X sky130_fd_sc_hd__and3_4
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _11737_/A VGND VGND VPWR VPWR _13992_/A sky130_fd_sc_hd__buf_2
XFILLER_41_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ _16203_/A _16201_/X _16203_/C VGND VGND VPWR VPWR _16203_/X sky130_fd_sc_hd__and3_4
XANTENNA__12558__A1 _11980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13415_ _13415_/A _13415_/B _13415_/C VGND VGND VPWR VPWR _13423_/B sky130_fd_sc_hd__or3_4
XANTENNA__17397__A _17178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17183_ _14263_/X _17137_/X _17182_/Y _17065_/X VGND VGND VPWR VPWR _17183_/X sky130_fd_sc_hd__o22a_4
X_14395_ _15618_/A _14305_/B VGND VGND VPWR VPWR _14396_/C sky130_fd_sc_hd__or2_4
XFILLER_70_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14814__A _14845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16134_ _16107_/A _16211_/B VGND VGND VPWR VPWR _16134_/X sky130_fd_sc_hd__or2_4
X_13346_ _15695_/A _13342_/X _13346_/C VGND VGND VPWR VPWR _13346_/X sky130_fd_sc_hd__or3_4
XANTENNA__15629__B _15573_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16065_ _16069_/A _23864_/Q VGND VGND VPWR VPWR _16065_/X sky130_fd_sc_hd__or2_4
X_13277_ _13277_/A _13276_/Y VGND VGND VPWR VPWR _13277_/X sky130_fd_sc_hd__or2_4
XANTENNA__12334__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15016_ _12301_/A _15016_/B _15015_/X VGND VGND VPWR VPWR _15017_/B sky130_fd_sc_hd__or3_4
XFILLER_64_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12228_ _12221_/X _12228_/B VGND VGND VPWR VPWR _12228_/X sky130_fd_sc_hd__or2_4
XFILLER_68_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21045__A2 _21044_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22242__B2 _22240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12053__B _23773_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19824_ _21581_/A VGND VGND VPWR VPWR _21112_/A sky130_fd_sc_hd__buf_2
XANTENNA__15645__A _13918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12159_ _11803_/A _12159_/B VGND VGND VPWR VPWR _12159_/X sky130_fd_sc_hd__or2_4
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19755_ _19720_/B VGND VGND VPWR VPWR _19755_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16967_ _17726_/A _18642_/A _17720_/A VGND VGND VPWR VPWR _18557_/A sky130_fd_sc_hd__or3_4
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18956__A _18971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13165__A _12745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22545__A2 _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18706_ _18681_/A _18705_/Y _17735_/X VGND VGND VPWR VPWR _18706_/X sky130_fd_sc_hd__a21o_4
X_15918_ _14075_/X _14265_/Y _14074_/X _15917_/Y VGND VGND VPWR VPWR _15919_/A sky130_fd_sc_hd__a211o_4
X_16898_ _16898_/A _16897_/X VGND VGND VPWR VPWR _16903_/C sky130_fd_sc_hd__nor2_4
X_19686_ _19686_/A _19861_/A VGND VGND VPWR VPWR _19867_/C sky130_fd_sc_hd__or2_4
X_15849_ _13548_/X _15849_/B VGND VGND VPWR VPWR _15849_/X sky130_fd_sc_hd__or2_4
X_18637_ _18082_/A _18042_/Y _17854_/X _18636_/X VGND VGND VPWR VPWR _18638_/A sky130_fd_sc_hd__a211o_4
XFILLER_77_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15380__A _15379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20308__A1 _17636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16907__C _16907_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18568_ _17390_/B _18566_/X _18063_/A _18567_/X VGND VGND VPWR VPWR _18568_/X sky130_fd_sc_hd__a211o_4
XFILLER_80_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17519_ _13270_/X _17510_/B VGND VGND VPWR VPWR _17519_/Y sky130_fd_sc_hd__nand2_4
XFILLER_75_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18499_ _18714_/A VGND VGND VPWR VPWR _18499_/X sky130_fd_sc_hd__buf_2
XFILLER_33_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12509__A _12509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20530_ _18256_/X _20424_/X _20516_/X _20529_/Y VGND VGND VPWR VPWR _20531_/A sky130_fd_sc_hd__a211o_4
XFILLER_32_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12228__B _12228_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20461_ _20588_/A _20461_/B VGND VGND VPWR VPWR _20461_/Y sky130_fd_sc_hd__nand2_4
XFILLER_53_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21808__B2 _21800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20445__B _20445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22200_ _11813_/B VGND VGND VPWR VPWR _22200_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17488__A1 _13350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23180_ _23404_/CLK _22546_/X VGND VGND VPWR VPWR _15462_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17488__B2 _17487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21284__A2 _21283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20392_ _24217_/Q _20282_/X _20391_/X VGND VGND VPWR VPWR _20393_/A sky130_fd_sc_hd__o21a_4
X_22131_ _22446_/A VGND VGND VPWR VPWR _22131_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12244__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22062_ _21857_/X _22059_/X _15296_/B _22056_/X VGND VGND VPWR VPWR _23458_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21036__A2 _21030_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21013_ _21012_/X VGND VGND VPWR VPWR _21013_/X sky130_fd_sc_hd__buf_2
XFILLER_99_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21972__A2_N _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19672__D _19672_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15555__A _15536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19027__A _19027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20795__A1 _24200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17660__A1 _16985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15274__B _15274_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18866__A _11599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22964_ _22982_/A _22962_/Y _22963_/X VGND VGND VPWR VPWR _22964_/X sky130_fd_sc_hd__and3_4
XFILLER_99_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20547__A1 _18283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22388__A _20276_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21915_ _23550_/Q VGND VGND VPWR VPWR _21915_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_70_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR _24305_/CLK sky130_fd_sc_hd__clkbuf_1
X_22895_ _22895_/A VGND VGND VPWR VPWR HADDR[2] sky130_fd_sc_hd__inv_2
XFILLER_56_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16386__A _15929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15290__A _14152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13803__A _13654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21846_ _21845_/X _21841_/X _23591_/Q _21836_/X VGND VGND VPWR VPWR _21846_/X sky130_fd_sc_hd__o22a_4
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14618__B _14698_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21777_ _21567_/X _21776_/X _14714_/B _21773_/X VGND VGND VPWR VPWR _23620_/D sky130_fd_sc_hd__o22a_4
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ _11530_/A _18959_/A VGND VGND VPWR VPWR _11530_/X sky130_fd_sc_hd__or2_4
X_23516_ _23515_/CLK _23516_/D VGND VGND VPWR VPWR _23516_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20728_ _20358_/B _20822_/B VGND VGND VPWR VPWR _20728_/X sky130_fd_sc_hd__or2_4
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20636__A _22112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23447_ _23383_/CLK _23447_/D VGND VGND VPWR VPWR _16189_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20659_ _20658_/X VGND VGND VPWR VPWR _20659_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14634__A _15036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13200_ _11850_/A _13200_/B VGND VGND VPWR VPWR _13200_/X sky130_fd_sc_hd__and2_4
X_14180_ _14225_/A _14078_/B VGND VGND VPWR VPWR _14183_/B sky130_fd_sc_hd__or2_4
X_23378_ _23314_/CLK _23378_/D VGND VGND VPWR VPWR _23378_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20483__B1 _20482_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13131_ _13109_/A _13129_/X _13131_/C VGND VGND VPWR VPWR _13131_/X sky130_fd_sc_hd__and3_4
X_22329_ _15212_/B VGND VGND VPWR VPWR _22329_/X sky130_fd_sc_hd__buf_2
XANTENNA__12154__A _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22224__A1 _22103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13062_ _13726_/A VGND VGND VPWR VPWR _15480_/A sky130_fd_sc_hd__buf_2
XANTENNA__22224__B2 _22219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21467__A _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17664__B _17664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12013_ _12020_/A VGND VGND VPWR VPWR _16541_/A sky130_fd_sc_hd__buf_2
XANTENNA__11993__A _11993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17870_ _17862_/X _17867_/X _17869_/X VGND VGND VPWR VPWR _17871_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__20786__A1 _20681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20786__B2 _20625_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16821_ _16897_/A _16820_/X _16897_/A _16820_/X VGND VGND VPWR VPWR _16821_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22527__A2 _22522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16752_ _16747_/X _16752_/B _16751_/X VGND VGND VPWR VPWR _16752_/X sky130_fd_sc_hd__and3_4
X_19540_ _19817_/C _19637_/A VGND VGND VPWR VPWR _19541_/B sky130_fd_sc_hd__or2_4
XANTENNA__17680__A _17680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13964_ _13968_/A _13964_/B _13964_/C VGND VGND VPWR VPWR _13965_/C sky130_fd_sc_hd__and3_4
XFILLER_19_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20538__A1 _20511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20538__B2 _20488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15703_ _12742_/A _15762_/B VGND VGND VPWR VPWR _15703_/X sky130_fd_sc_hd__or2_4
XFILLER_111_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12915_ _12915_/A _23091_/Q VGND VGND VPWR VPWR _12915_/X sky130_fd_sc_hd__or2_4
X_16683_ _16686_/A _16744_/B VGND VGND VPWR VPWR _16683_/X sky130_fd_sc_hd__or2_4
X_19471_ _19471_/A VGND VGND VPWR VPWR _19754_/A sky130_fd_sc_hd__buf_2
XFILLER_47_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15912__B _15911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18926__D _18934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13895_ _13895_/A _13815_/B VGND VGND VPWR VPWR _13895_/X sky130_fd_sc_hd__or2_4
XANTENNA__16296__A _11884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15634_ _14499_/A _15634_/B _15634_/C VGND VGND VPWR VPWR _15635_/C sky130_fd_sc_hd__and3_4
X_18422_ _18244_/A _18419_/Y _18420_/Y _18421_/X VGND VGND VPWR VPWR _18422_/X sky130_fd_sc_hd__or4_4
XFILLER_64_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13713__A _13697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12846_ _12435_/A VGND VGND VPWR VPWR _12849_/A sky130_fd_sc_hd__buf_2
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18353_ _18383_/A _18383_/B _18342_/A VGND VGND VPWR VPWR _18354_/B sky130_fd_sc_hd__o21ai_4
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15565_ _11859_/A _15561_/X _15565_/C VGND VGND VPWR VPWR _15565_/X sky130_fd_sc_hd__or3_4
X_12777_ _13087_/A VGND VGND VPWR VPWR _12777_/X sky130_fd_sc_hd__buf_2
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18903__A1 _17191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12329__A _12711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17304_ _17297_/X _17309_/B VGND VGND VPWR VPWR _17305_/A sky130_fd_sc_hd__or2_4
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14536_/A _14516_/B VGND VGND VPWR VPWR _14517_/C sky130_fd_sc_hd__or2_4
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _11727_/X VGND VGND VPWR VPWR _16048_/A sky130_fd_sc_hd__buf_2
X_18284_ _18171_/X _18262_/X _18202_/X _18283_/X VGND VGND VPWR VPWR _18284_/X sky130_fd_sc_hd__o22a_4
X_15496_ _13735_/A _15432_/B VGND VGND VPWR VPWR _15496_/X sky130_fd_sc_hd__or2_4
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__B _23741_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17235_ _17251_/A _17226_/Y _17824_/A _17234_/Y VGND VGND VPWR VPWR _17235_/X sky130_fd_sc_hd__o22a_4
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14447_ _12885_/A _14447_/B VGND VGND VPWR VPWR _14447_/X sky130_fd_sc_hd__or2_4
X_11659_ _11658_/X VGND VGND VPWR VPWR _16077_/A sky130_fd_sc_hd__buf_2
XFILLER_35_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14544__A _13711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17166_ _14565_/Y _17100_/X _17165_/Y _17065_/X VGND VGND VPWR VPWR _17166_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18667__B1 _18198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14378_ _15598_/A _14283_/B VGND VGND VPWR VPWR _14378_/X sky130_fd_sc_hd__or2_4
XANTENNA__22463__B2 _22386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16117_ _16090_/A VGND VGND VPWR VPWR _16145_/A sky130_fd_sc_hd__buf_2
XFILLER_7_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13329_ _13301_/A _13329_/B VGND VGND VPWR VPWR _13329_/X sky130_fd_sc_hd__or2_4
X_17097_ _17097_/A VGND VGND VPWR VPWR _17097_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16048_ _16048_/A _16046_/X _16047_/X VGND VGND VPWR VPWR _16052_/B sky130_fd_sc_hd__and3_4
XANTENNA__12999__A _12852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15375__A _12598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20777__A1 _24201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19807_ _19710_/X _19800_/X _19806_/X _18759_/A _19490_/X VGND VGND VPWR VPWR _24171_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24338__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17999_ _17569_/A _17995_/X _17998_/X VGND VGND VPWR VPWR _17999_/Y sky130_fd_sc_hd__a21oi_4
X_19738_ _19419_/X _19737_/X _12101_/X _19678_/X VGND VGND VPWR VPWR _19738_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23392__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19395__B2 _24204_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15822__B _23821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19669_ _19668_/X VGND VGND VPWR VPWR _19669_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14719__A _13918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_57_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17945__A2 _17898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21700_ _21522_/X _21698_/X _23671_/Q _21695_/X VGND VGND VPWR VPWR _21700_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13623__A _13623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22680_ _21804_/A _22679_/X _23096_/Q _22676_/X VGND VGND VPWR VPWR _22680_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21631_ _21576_/X _21626_/X _14860_/B _21595_/A VGND VGND VPWR VPWR _21631_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17158__B1 _17156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16934__A _18171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12239__A _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24350_ _24344_/CLK _18929_/X HRESETn VGND VGND VPWR VPWR _24350_/Q sky130_fd_sc_hd__dfstp_4
X_21562_ _20838_/A VGND VGND VPWR VPWR _21562_/X sky130_fd_sc_hd__buf_2
XANTENNA__16905__B1 _16897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23301_ _24008_/CLK _23301_/D VGND VGND VPWR VPWR _22325_/A sky130_fd_sc_hd__dfxtp_4
X_20513_ _18577_/Y VGND VGND VPWR VPWR _20534_/A sky130_fd_sc_hd__buf_2
X_21493_ _21285_/X _21491_/X _14777_/B _21488_/X VGND VGND VPWR VPWR _23779_/D sky130_fd_sc_hd__o22a_4
X_24281_ _24344_/CLK _24281_/D HRESETn VGND VGND VPWR VPWR _19230_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_21_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14454__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20444_ _20444_/A VGND VGND VPWR VPWR _20444_/X sky130_fd_sc_hd__buf_2
X_23232_ _23233_/CLK _22461_/X VGND VGND VPWR VPWR _14856_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21257__A2 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22671__A _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20465__B1 _12316_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20375_ _20280_/X _20373_/X _24090_/Q _20374_/X VGND VGND VPWR VPWR _20375_/X sky130_fd_sc_hd__o22a_4
X_23163_ _24059_/CLK _23163_/D VGND VGND VPWR VPWR _16767_/B sky130_fd_sc_hd__dfxtp_4
X_22114_ _22112_/X _22113_/X _15677_/B _22108_/X VGND VGND VPWR VPWR _23438_/D sky130_fd_sc_hd__o22a_4
X_23094_ _23473_/CLK _23094_/D VGND VGND VPWR VPWR _12328_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22206__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17881__B2 _17880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22045_ _22031_/A VGND VGND VPWR VPWR _22045_/X sky130_fd_sc_hd__buf_2
XFILLER_0_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15285__A _14149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12702__A _15664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22509__A2 _22507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23996_ _24092_/CLK _21121_/X VGND VGND VPWR VPWR _23996_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21717__B1 _23659_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23007__A _23006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22947_ _22924_/X _18349_/A _22937_/X _22946_/X VGND VGND VPWR VPWR _22948_/A sky130_fd_sc_hd__a211o_4
XFILLER_84_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21193__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12700_ _12711_/A VGND VGND VPWR VPWR _12722_/A sky130_fd_sc_hd__buf_2
X_13680_ _15448_/A _13678_/X _13680_/C VGND VGND VPWR VPWR _13681_/C sky130_fd_sc_hd__and3_4
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22878_ _22872_/A _22878_/B VGND VGND VPWR VPWR HWDATA[30] sky130_fd_sc_hd__nor2_4
XFILLER_16_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12631_ _13737_/A VGND VGND VPWR VPWR _12954_/A sky130_fd_sc_hd__buf_2
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21829_ _21817_/A VGND VGND VPWR VPWR _21829_/X sky130_fd_sc_hd__buf_2
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22142__B1 _15277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15350_ _15334_/A _15350_/B _15350_/C VGND VGND VPWR VPWR _15354_/B sky130_fd_sc_hd__and3_4
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_0_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR _24202_/CLK sky130_fd_sc_hd__clkbuf_1
X_12562_ _13908_/A VGND VGND VPWR VPWR _13738_/A sky130_fd_sc_hd__buf_2
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21496__A2 _21491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14301_ _12257_/A _14301_/B VGND VGND VPWR VPWR _14301_/X sky130_fd_sc_hd__or2_4
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11513_ _24328_/Q _11513_/B VGND VGND VPWR VPWR _11514_/B sky130_fd_sc_hd__or2_4
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11988__A _16143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15281_ _11847_/A _15258_/X _15265_/X _15272_/X _15280_/X VGND VGND VPWR VPWR _15281_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12493_/A _12489_/X _12493_/C VGND VGND VPWR VPWR _12503_/B sky130_fd_sc_hd__and3_4
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17020_ _17020_/A VGND VGND VPWR VPWR _17021_/A sky130_fd_sc_hd__buf_2
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _14246_/A _14232_/B _14231_/X VGND VGND VPWR VPWR _14232_/X sky130_fd_sc_hd__and3_4
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21248__A2 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23265__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22445__B2 _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19310__B2 _19303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14163_ _14146_/X _14153_/X _14163_/C VGND VGND VPWR VPWR _14163_/X sky130_fd_sc_hd__or3_4
X_13114_ _13098_/A _23378_/Q VGND VGND VPWR VPWR _13116_/B sky130_fd_sc_hd__or2_4
XFILLER_98_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21197__A _21168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14094_ _12880_/A VGND VGND VPWR VPWR _15011_/A sky130_fd_sc_hd__buf_2
X_18971_ _18971_/A VGND VGND VPWR VPWR _18971_/X sky130_fd_sc_hd__buf_2
XFILLER_98_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15195__A _14195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13045_ _12553_/A _13045_/B VGND VGND VPWR VPWR _13045_/X sky130_fd_sc_hd__or2_4
X_17922_ _17911_/X _17233_/X _17912_/X _17211_/X VGND VGND VPWR VPWR _17922_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__13708__A _13708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12612__A _12612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18002__C _17762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21420__A2 _21419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17853_ _17853_/A VGND VGND VPWR VPWR _17853_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16804_ _16768_/X _24091_/Q VGND VGND VPWR VPWR _16805_/C sky130_fd_sc_hd__or2_4
XFILLER_78_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24105__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14996_ _14121_/A _23167_/Q VGND VGND VPWR VPWR _14998_/B sky130_fd_sc_hd__or2_4
X_17784_ _18442_/A VGND VGND VPWR VPWR _18206_/A sky130_fd_sc_hd__buf_2
XFILLER_82_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16738__B _23867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19523_ _19523_/A _19523_/B VGND VGND VPWR VPWR _19524_/B sky130_fd_sc_hd__or2_4
X_13947_ _12217_/A _13947_/B _13947_/C VGND VGND VPWR VPWR _13948_/C sky130_fd_sc_hd__and3_4
X_16735_ _11921_/X _23803_/Q VGND VGND VPWR VPWR _16736_/C sky130_fd_sc_hd__or2_4
XANTENNA__21184__A1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21184__B2 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13443__A _13437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16666_ _16670_/A _23868_/Q VGND VGND VPWR VPWR _16666_/X sky130_fd_sc_hd__or2_4
X_19454_ _19454_/A _19453_/Y VGND VGND VPWR VPWR _19454_/X sky130_fd_sc_hd__or2_4
X_13878_ _13878_/A _13791_/B VGND VGND VPWR VPWR _13880_/B sky130_fd_sc_hd__or2_4
XFILLER_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20931__A1 _18679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15617_ _15617_/A _23595_/Q VGND VGND VPWR VPWR _15619_/B sky130_fd_sc_hd__or2_4
X_18405_ _18405_/A _18404_/X VGND VGND VPWR VPWR _18405_/X sky130_fd_sc_hd__or2_4
X_12829_ _12829_/A _23860_/Q VGND VGND VPWR VPWR _12830_/C sky130_fd_sc_hd__or2_4
XFILLER_90_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16597_ _11675_/X VGND VGND VPWR VPWR _16597_/X sky130_fd_sc_hd__buf_2
X_19385_ _19385_/A VGND VGND VPWR VPWR _19385_/X sky130_fd_sc_hd__buf_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15548_ _12861_/A _15546_/X _15547_/X VGND VGND VPWR VPWR _15548_/X sky130_fd_sc_hd__and3_4
X_18336_ _18285_/C _17759_/X _17680_/X VGND VGND VPWR VPWR _18336_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21487__A2 _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22684__B2 _22683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20276__A _20276_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23608__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11898__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18267_ _18267_/A _18267_/B _18265_/Y _18267_/D VGND VGND VPWR VPWR _18268_/A sky130_fd_sc_hd__or4_4
X_15479_ _12646_/A _15477_/X _15478_/X VGND VGND VPWR VPWR _15479_/X sky130_fd_sc_hd__and3_4
XANTENNA__14274__A _15412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17218_ _17007_/X _17155_/X _14988_/X _17186_/X VGND VGND VPWR VPWR _17218_/X sky130_fd_sc_hd__o22a_4
X_18198_ _18198_/A VGND VGND VPWR VPWR _18198_/X sky130_fd_sc_hd__buf_2
XFILLER_89_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22436__B2 _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19784__B _19784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24190__CLK _24187_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12924__A1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17149_ _17220_/A _17140_/Y _17160_/A _17148_/Y VGND VGND VPWR VPWR _17149_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12924__B2 _12923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23758__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20160_ _20160_/A _20159_/Y VGND VGND VPWR VPWR _20160_/X sky130_fd_sc_hd__or2_4
XFILLER_89_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14721__B _14723_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13618__A _13614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20091_ _20091_/A VGND VGND VPWR VPWR _20091_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18407__A3 _18393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12522__A _12522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21947__B1 _15802_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15833__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23850_ _23819_/CLK _23850_/D VGND VGND VPWR VPWR _23850_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22801_ _22807_/A _15120_/Y VGND VGND VPWR VPWR _22801_/X sky130_fd_sc_hd__or2_4
XFILLER_113_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15552__B _23883_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23781_ _23781_/CLK _23781_/D VGND VGND VPWR VPWR _14484_/B sky130_fd_sc_hd__dfxtp_4
X_20993_ _20494_/A _20992_/X _24319_/Q _20453_/A VGND VGND VPWR VPWR _20993_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14449__A _13019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23138__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21175__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22732_ SYSTICKCLKDIV[3] _22730_/Y SYSTICKCLKDIV[2] _22756_/A VGND VGND VPWR VPWR
+ _22732_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22663_ _22462_/X _22636_/A _23103_/Q _22626_/A VGND VGND VPWR VPWR _22663_/X sky130_fd_sc_hd__o22a_4
XFILLER_94_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16664__A _16652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24402_ _23326_/CLK _18838_/X HRESETn VGND VGND VPWR VPWR _24402_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21614_ _21546_/X _21612_/X _15849_/B _21609_/X VGND VGND VPWR VPWR _21614_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21478__A2 _21477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22594_ _22427_/X _22593_/X _15732_/B _22590_/X VGND VGND VPWR VPWR _23150_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22675__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16383__B _16383_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24333_ _24365_/CLK _24333_/D HRESETn VGND VGND VPWR VPWR _24333_/Q sky130_fd_sc_hd__dfstp_4
X_21545_ _21543_/X _21544_/X _15722_/B _21539_/X VGND VGND VPWR VPWR _23758_/D sky130_fd_sc_hd__o22a_4
X_24264_ _24305_/CLK _24264_/D HRESETn VGND VGND VPWR VPWR _19213_/A sky130_fd_sc_hd__dfrtp_4
X_21476_ _21256_/X _21470_/X _13485_/B _21474_/X VGND VGND VPWR VPWR _21476_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20438__B1 _20437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23215_ _24082_/CLK _23215_/D VGND VGND VPWR VPWR _13568_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20427_ _20427_/A VGND VGND VPWR VPWR _20427_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24195_ _24199_/CLK _24195_/D HRESETn VGND VGND VPWR VPWR _24195_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19843__A2 _19837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23146_ _23561_/CLK _23146_/D VGND VGND VPWR VPWR _14025_/B sky130_fd_sc_hd__dfxtp_4
X_20358_ _20342_/A _20358_/B VGND VGND VPWR VPWR _20358_/X sky130_fd_sc_hd__and2_4
XANTENNA__21650__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13528__A _13507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20289_ _20424_/A VGND VGND VPWR VPWR _20578_/A sky130_fd_sc_hd__buf_2
X_23077_ _23973_/CLK _22706_/X VGND VGND VPWR VPWR _14547_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_4_2_0_HCLK_A clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12432__A _12338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22028_ _22020_/X VGND VGND VPWR VPWR _22028_/X sky130_fd_sc_hd__buf_2
XANTENNA__21745__A _21737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14850_ _14073_/A _14818_/X _14850_/C VGND VGND VPWR VPWR _14851_/A sky130_fd_sc_hd__and3_4
XANTENNA__15743__A _15743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24321__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13801_ _13659_/A _13873_/B VGND VGND VPWR VPWR _13801_/X sky130_fd_sc_hd__or2_4
XFILLER_21_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14781_ _12217_/A _14781_/B _14781_/C VGND VGND VPWR VPWR _14782_/C sky130_fd_sc_hd__and3_4
XFILLER_40_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15462__B _15462_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11993_ _11993_/A _23902_/Q VGND VGND VPWR VPWR _11995_/B sky130_fd_sc_hd__or2_4
X_23979_ _23688_/CLK _23979_/D VGND VGND VPWR VPWR _23979_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16520_ _16239_/X _16520_/B VGND VGND VPWR VPWR _16520_/X sky130_fd_sc_hd__or2_4
XANTENNA__13263__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13732_ _15493_/A _13627_/B VGND VGND VPWR VPWR _13732_/X sky130_fd_sc_hd__or2_4
XFILLER_17_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22576__A _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_40_0_HCLK clkbuf_6_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_40_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16451_ _11713_/X VGND VGND VPWR VPWR _16465_/A sky130_fd_sc_hd__buf_2
X_13663_ _15431_/A _13660_/X _13662_/X VGND VGND VPWR VPWR _13663_/X sky130_fd_sc_hd__and3_4
XFILLER_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15402_ _13622_/A _15465_/B VGND VGND VPWR VPWR _15402_/X sky130_fd_sc_hd__or2_4
X_12614_ _12604_/A _12614_/B VGND VGND VPWR VPWR _12614_/X sky130_fd_sc_hd__or2_4
X_19170_ _24303_/Q _19124_/B _19169_/Y VGND VGND VPWR VPWR _24303_/D sky130_fd_sc_hd__o21a_4
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16382_ _15948_/A _16380_/X _16382_/C VGND VGND VPWR VPWR _16382_/X sky130_fd_sc_hd__and3_4
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21469__A2 _21463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13594_ _11841_/A VGND VGND VPWR VPWR _13594_/X sky130_fd_sc_hd__buf_2
XANTENNA__20096__A NMI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18121_ _18107_/A _18081_/B _17259_/A _17531_/X VGND VGND VPWR VPWR _18121_/X sky130_fd_sc_hd__o22a_4
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15333_ _15333_/A _15274_/B VGND VGND VPWR VPWR _15334_/C sky130_fd_sc_hd__or2_4
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12545_ _12553_/A VGND VGND VPWR VPWR _12546_/A sky130_fd_sc_hd__buf_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18052_ _16924_/X VGND VGND VPWR VPWR _18224_/A sky130_fd_sc_hd__buf_2
X_15264_ _12860_/A _15262_/X _15263_/X VGND VGND VPWR VPWR _15264_/X sky130_fd_sc_hd__and3_4
X_12476_ _13020_/A VGND VGND VPWR VPWR _13029_/A sky130_fd_sc_hd__buf_2
X_17003_ _17003_/A VGND VGND VPWR VPWR _17003_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12326__B _12317_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14215_ _14215_/A _14215_/B _14215_/C VGND VGND VPWR VPWR _14221_/B sky130_fd_sc_hd__and3_4
X_15195_ _14195_/A _15193_/X _15195_/C VGND VGND VPWR VPWR _15199_/B sky130_fd_sc_hd__and3_4
XANTENNA__14822__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14146_ _14119_/X VGND VGND VPWR VPWR _14146_/X sky130_fd_sc_hd__buf_2
XFILLER_119_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15637__B _24075_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13438__A _13437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14077_ _14074_/X _14076_/Y VGND VGND VPWR VPWR _14077_/X sky130_fd_sc_hd__or2_4
X_18954_ _18954_/A VGND VGND VPWR VPWR _18954_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12342__A _13726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13028_ _12518_/A _13104_/B VGND VGND VPWR VPWR _13028_/X sky130_fd_sc_hd__or2_4
X_17905_ _17905_/A VGND VGND VPWR VPWR _17905_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21655__A _21662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18885_ _18892_/A VGND VGND VPWR VPWR _18885_/X sky130_fd_sc_hd__buf_2
XFILLER_117_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15653__A _12691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17836_ _17836_/A VGND VGND VPWR VPWR _17836_/X sky130_fd_sc_hd__buf_2
XFILLER_39_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_122_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR _23859_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16468__B _16408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17767_ _17946_/B _17765_/X _17946_/A VGND VGND VPWR VPWR _17767_/X sky130_fd_sc_hd__a21bo_4
XFILLER_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14979_ _14925_/A _14979_/B _14978_/X VGND VGND VPWR VPWR _14983_/B sky130_fd_sc_hd__and3_4
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14269__A _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21157__B2 _21151_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18964__A _18994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19506_ _19744_/A _19541_/A VGND VGND VPWR VPWR _19718_/A sky130_fd_sc_hd__or2_4
XFILLER_35_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13173__A _12255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16718_ _16718_/A _16718_/B _16717_/X VGND VGND VPWR VPWR _16719_/C sky130_fd_sc_hd__and3_4
XFILLER_63_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17698_ _17698_/A _17696_/A VGND VGND VPWR VPWR _17698_/X sky130_fd_sc_hd__or2_4
XFILLER_50_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19437_ HRDATA[1] VGND VGND VPWR VPWR _19437_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16649_ _16616_/A _16649_/B _16649_/C VGND VGND VPWR VPWR _16653_/B sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_4_13_0_HCLK_A clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19368_ _19367_/X _17775_/X _19367_/X _24220_/Q VGND VGND VPWR VPWR _19368_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18319_ _18206_/A _17492_/X VGND VGND VPWR VPWR _18319_/X sky130_fd_sc_hd__and2_4
XANTENNA__13620__B _13713_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19299_ _19205_/B VGND VGND VPWR VPWR _19299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23580__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21330_ _21316_/A VGND VGND VPWR VPWR _21330_/X sky130_fd_sc_hd__buf_2
XANTENNA__12236__B _12236_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18089__A1 _17762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21261_ _21831_/A VGND VGND VPWR VPWR _21261_/X sky130_fd_sc_hd__buf_2
XANTENNA__15828__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14732__A _14158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19825__A2 _19672_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18204__A _18204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23000_ _22989_/A _23000_/B _23000_/C VGND VGND VPWR VPWR _23000_/X sky130_fd_sc_hd__and3_4
X_20212_ _16907_/C _18757_/X _20516_/A VGND VGND VPWR VPWR _20212_/X sky130_fd_sc_hd__o21a_4
XFILLER_11_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21192_ _20671_/X _21190_/X _15815_/B _21187_/X VGND VGND VPWR VPWR _21192_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21632__A2 _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15547__B _23435_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20143_ _24424_/Q VGND VGND VPWR VPWR _20143_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19589__A1 _20358_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20074_ _11622_/A _20073_/X VGND VGND VPWR VPWR _20074_/Y sky130_fd_sc_hd__nor2_4
XFILLER_83_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16659__A _16640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21396__B2 _21359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23902_ _23320_/CLK _21303_/X VGND VGND VPWR VPWR _23902_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15563__A _15556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18261__A1 _17672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23833_ _23770_/CLK _23833_/D VGND VGND VPWR VPWR _16280_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21148__B2 _21144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22345__B1 _16391_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18874__A _18898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13083__A _13083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23764_ _24021_/CLK _21530_/X VGND VGND VPWR VPWR _12774_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21699__A2 _21698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20976_ _20976_/A VGND VGND VPWR VPWR _20976_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22396__A _20355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_27_0_HCLK clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22715_ _19770_/X _16996_/A _20576_/B VGND VGND VPWR VPWR _22723_/B sky130_fd_sc_hd__and3_4
X_23695_ _23987_/CLK _21661_/X VGND VGND VPWR VPWR _13487_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16394__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14907__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13811__A _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22646_ _22432_/X _22643_/X _15493_/B _22640_/X VGND VGND VPWR VPWR _23116_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22648__B2 _22647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22577_ _22398_/X _22572_/X _16407_/B _22576_/X VGND VGND VPWR VPWR _23162_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12427__A _13572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21320__B2 _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12330_ _12744_/A _12328_/X _12330_/C VGND VGND VPWR VPWR _12334_/B sky130_fd_sc_hd__and3_4
X_24316_ _24290_/CLK _19144_/X HRESETn VGND VGND VPWR VPWR _19137_/A sky130_fd_sc_hd__dfrtp_4
X_21528_ _21526_/X _21520_/X _12463_/B _21527_/X VGND VGND VPWR VPWR _21528_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12261_ _12260_/X VGND VGND VPWR VPWR _12743_/A sky130_fd_sc_hd__buf_2
X_24247_ _24216_/CLK _24247_/D HRESETn VGND VGND VPWR VPWR _24247_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15738__A _12794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21459_ _21227_/X _21456_/X _23803_/Q _21453_/X VGND VGND VPWR VPWR _21459_/X sky130_fd_sc_hd__o22a_4
X_14000_ _14000_/A VGND VGND VPWR VPWR _14021_/A sky130_fd_sc_hd__buf_2
XANTENNA__21084__B1 _24018_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12192_ _15412_/A VGND VGND VPWR VPWR _13055_/A sky130_fd_sc_hd__buf_2
X_24178_ _23584_/CLK _19738_/X HRESETn VGND VGND VPWR VPWR _14101_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20082__C _20076_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23129_ _23130_/CLK _23129_/D VGND VGND VPWR VPWR _16279_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13258__A _12350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15951_ _15984_/A _24024_/Q VGND VGND VPWR VPWR _15953_/B sky130_fd_sc_hd__or2_4
XANTENNA__17672__B _17497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16569__A _16569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22584__B1 _12620_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14902_ _15146_/A _23456_/Q VGND VGND VPWR VPWR _14902_/X sky130_fd_sc_hd__or2_4
XFILLER_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15882_ _15882_/A _15878_/X _15882_/C VGND VGND VPWR VPWR _15882_/X sky130_fd_sc_hd__or3_4
X_18670_ _18142_/A _17615_/X _18398_/X _17333_/X VGND VGND VPWR VPWR _18670_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__15904__C _15904_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17621_ _17621_/A _17421_/A _17621_/C _17621_/D VGND VGND VPWR VPWR _17622_/B sky130_fd_sc_hd__or4_4
XFILLER_40_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14833_ _11766_/A _14833_/B _14832_/X VGND VGND VPWR VPWR _14833_/X sky130_fd_sc_hd__and3_4
XFILLER_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21139__B2 _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14764_ _13603_/A _14762_/X _14763_/X VGND VGND VPWR VPWR _14764_/X sky130_fd_sc_hd__and3_4
X_17552_ _17552_/A _17457_/B VGND VGND VPWR VPWR _17552_/X sky130_fd_sc_hd__and2_4
X_11976_ _11976_/A VGND VGND VPWR VPWR _15420_/A sky130_fd_sc_hd__buf_2
X_13715_ _12617_/A VGND VGND VPWR VPWR _15495_/A sky130_fd_sc_hd__buf_2
X_16503_ _16355_/X _16499_/X _16503_/C VGND VGND VPWR VPWR _16503_/X sky130_fd_sc_hd__or3_4
XANTENNA__20898__B1 _20895_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17483_ _13591_/X _17480_/X VGND VGND VPWR VPWR _17483_/X sky130_fd_sc_hd__and2_4
X_14695_ _14679_/A _14695_/B VGND VGND VPWR VPWR _14695_/X sky130_fd_sc_hd__or2_4
XANTENNA__14817__A _11766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19222_ _24273_/Q _19263_/A VGND VGND VPWR VPWR _19261_/A sky130_fd_sc_hd__and2_4
XANTENNA__13721__A _13747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13646_ _13677_/A _13644_/X _13646_/C VGND VGND VPWR VPWR _13646_/X sky130_fd_sc_hd__and3_4
X_16434_ _16394_/X _16434_/B VGND VGND VPWR VPWR _16434_/X sky130_fd_sc_hd__or2_4
XFILLER_60_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22639__B2 _22633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16365_ _16365_/A _16365_/B VGND VGND VPWR VPWR _16366_/C sky130_fd_sc_hd__or2_4
X_19153_ _19132_/X VGND VGND VPWR VPWR _19153_/Y sky130_fd_sc_hd__inv_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13577_ _13493_/X _13577_/B VGND VGND VPWR VPWR _13578_/A sky130_fd_sc_hd__or2_4
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21311__B2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15316_ _13708_/A VGND VGND VPWR VPWR _15334_/A sky130_fd_sc_hd__buf_2
X_18104_ _18297_/A _17565_/Y VGND VGND VPWR VPWR _18105_/D sky130_fd_sc_hd__and2_4
XFILLER_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12528_ _12528_/A _12528_/B _12528_/C VGND VGND VPWR VPWR _12528_/X sky130_fd_sc_hd__or3_4
X_16296_ _11884_/X _16296_/B VGND VGND VPWR VPWR _16296_/X sky130_fd_sc_hd__or2_4
X_19084_ _18999_/A VGND VGND VPWR VPWR _19084_/X sky130_fd_sc_hd__buf_2
XANTENNA__21862__A2 _21853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_47_0_HCLK clkbuf_7_46_0_HCLK/A VGND VGND VPWR VPWR _23336_/CLK sky130_fd_sc_hd__clkbuf_1
X_15247_ _14202_/A _15247_/B _15246_/X VGND VGND VPWR VPWR _15248_/C sky130_fd_sc_hd__and3_4
X_18035_ _17837_/A _18033_/X _17845_/X _18034_/X VGND VGND VPWR VPWR _18035_/X sky130_fd_sc_hd__o22a_4
X_12459_ _12459_/A VGND VGND VPWR VPWR _12460_/A sky130_fd_sc_hd__buf_2
XANTENNA__14552__A _13711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15178_ _11608_/A _15178_/B _15177_/X VGND VGND VPWR VPWR _15178_/X sky130_fd_sc_hd__and3_4
XANTENNA__22811__A1 _17339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21614__A2 _21612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14271__B _14271_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14129_ _11847_/A _14086_/X _14099_/X _14118_/X _14128_/X VGND VGND VPWR VPWR _14129_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13168__A _12713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24120__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19986_ _19986_/A VGND VGND VPWR VPWR _19986_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12072__A _12068_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18937_ _18971_/A VGND VGND VPWR VPWR _18937_/X sky130_fd_sc_hd__buf_2
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21378__B2 _21373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19440__B1 _19437_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18868_ _18867_/X VGND VGND VPWR VPWR _20425_/A sky130_fd_sc_hd__buf_2
X_17819_ _17802_/X _17166_/X _17804_/X _17153_/X VGND VGND VPWR VPWR _17819_/X sky130_fd_sc_hd__o22a_4
X_18799_ _17178_/X _18795_/X _24424_/Q _18796_/X VGND VGND VPWR VPWR _18799_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18694__A _18327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20830_ _20732_/X _20829_/X _24294_/Q _20739_/X VGND VGND VPWR VPWR _20831_/B sky130_fd_sc_hd__o22a_4
XFILLER_19_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20761_ _24393_/Q _20595_/B VGND VGND VPWR VPWR _20761_/Y sky130_fd_sc_hd__nand2_4
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22500_ _22471_/A VGND VGND VPWR VPWR _22500_/X sky130_fd_sc_hd__buf_2
XANTENNA__13631__A _13631_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17103__A _18713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23480_ _23539_/CLK _22032_/X VGND VGND VPWR VPWR _23480_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20692_ _20288_/X VGND VGND VPWR VPWR _20692_/X sky130_fd_sc_hd__buf_2
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22431_ _22430_/X _22428_/X _15845_/B _22423_/X VGND VGND VPWR VPWR _23245_/D sky130_fd_sc_hd__o22a_4
XFILLER_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12247__A _12240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22362_ _22112_/X _22361_/X _15725_/B _22358_/X VGND VGND VPWR VPWR _22362_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20464__A _20464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24101_ _24321_/CLK _24101_/D HRESETn VGND VGND VPWR VPWR _24101_/Q sky130_fd_sc_hd__dfrtp_4
X_21313_ _21234_/X _21312_/X _23896_/Q _21309_/X VGND VGND VPWR VPWR _21313_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22293_ _22286_/A VGND VGND VPWR VPWR _22293_/X sky130_fd_sc_hd__buf_2
XANTENNA__14462__A _12441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24032_ _24032_/CLK _21056_/X VGND VGND VPWR VPWR _14892_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_11_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21244_ _20509_/A VGND VGND VPWR VPWR _21244_/X sky130_fd_sc_hd__buf_2
XANTENNA__22802__A1 _13685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15277__B _15277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_4_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21175_ _20394_/X _21169_/X _16273_/B _21173_/X VGND VGND VPWR VPWR _21175_/X sky130_fd_sc_hd__o22a_4
XFILLER_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20126_ _20077_/D _20125_/X VGND VGND VPWR VPWR _20126_/X sky130_fd_sc_hd__or2_4
XFILLER_63_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23476__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16389__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15293__A _14161_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20057_ _20057_/A VGND VGND VPWR VPWR _20057_/X sky130_fd_sc_hd__buf_2
XANTENNA__12710__A _12710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11830_ _11730_/X _11830_/B _11830_/C VGND VGND VPWR VPWR _11834_/B sky130_fd_sc_hd__and3_4
X_23816_ _23816_/CLK _21435_/X VGND VGND VPWR VPWR _13662_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20639__A _20421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23015__A _23015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11820_/A _11761_/B _11760_/X VGND VGND VPWR VPWR _11761_/X sky130_fd_sc_hd__and3_4
X_23747_ _23363_/CLK _23747_/D VGND VGND VPWR VPWR _14733_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ _20872_/X _20958_/X _15241_/B _20202_/X VGND VGND VPWR VPWR _20959_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20344__A2 _18814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14637__A _14782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _12982_/A VGND VGND VPWR VPWR _13500_/X sky130_fd_sc_hd__buf_2
XFILLER_42_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20358__B _20358_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17013__A _17013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13541__A _12413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _12512_/A _14480_/B VGND VGND VPWR VPWR _14481_/C sky130_fd_sc_hd__or2_4
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11691_/X VGND VGND VPWR VPWR _11692_/X sky130_fd_sc_hd__buf_2
X_23678_ _23774_/CLK _23678_/D VGND VGND VPWR VPWR _21683_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14356__B _14276_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _13463_/A _13504_/B VGND VGND VPWR VPWR _13431_/X sky130_fd_sc_hd__or2_4
XANTENNA__20077__C _20076_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22629_ _22636_/A VGND VGND VPWR VPWR _22629_/X sky130_fd_sc_hd__buf_2
XFILLER_70_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22097__A2 _22089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12157__A _12169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19498__B1 _19497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16150_ _16150_/A _16220_/B VGND VGND VPWR VPWR _16150_/X sky130_fd_sc_hd__or2_4
XFILLER_10_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13362_ _13357_/X _13362_/B _13362_/C VGND VGND VPWR VPWR _13363_/C sky130_fd_sc_hd__and3_4
XFILLER_107_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17667__B _17667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21844__A2 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20374__A _20202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15101_ _14055_/A _15093_/X _15100_/X VGND VGND VPWR VPWR _15101_/X sky130_fd_sc_hd__and3_4
XFILLER_5_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12313_ _11955_/A VGND VGND VPWR VPWR _15553_/A sky130_fd_sc_hd__buf_2
X_16081_ _16081_/A _16080_/Y VGND VGND VPWR VPWR _16081_/X sky130_fd_sc_hd__or2_4
X_13293_ _12540_/A _13291_/X _13293_/C VGND VGND VPWR VPWR _13293_/X sky130_fd_sc_hd__and3_4
X_15032_ _15032_/A _15032_/B _15032_/C VGND VGND VPWR VPWR _15032_/X sky130_fd_sc_hd__or3_4
XANTENNA__12337__A2 _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21057__B1 _15023_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12244_ _13055_/A VGND VGND VPWR VPWR _12706_/A sky130_fd_sc_hd__buf_2
XANTENNA__15187__B _15126_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23819__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12604__B _24021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19840_ _19819_/X _19839_/X _19766_/A VGND VGND VPWR VPWR _19840_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_29_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12175_ _11734_/A _24093_/Q VGND VGND VPWR VPWR _12175_/X sky130_fd_sc_hd__or2_4
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19771_ _19674_/X _19769_/Y _19770_/X _19551_/A VGND VGND VPWR VPWR _19771_/X sky130_fd_sc_hd__a2bb2o_4
X_16983_ _16945_/Y _16982_/X VGND VGND VPWR VPWR _16983_/X sky130_fd_sc_hd__or2_4
XFILLER_104_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16299__A _15929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18722_ _16935_/A _18710_/X _18485_/X _22824_/B VGND VGND VPWR VPWR _18722_/X sky130_fd_sc_hd__o22a_4
X_15934_ _15956_/A VGND VGND VPWR VPWR _15934_/X sky130_fd_sc_hd__buf_2
XFILLER_110_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23969__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18653_ _19994_/A VGND VGND VPWR VPWR _18653_/X sky130_fd_sc_hd__buf_2
XFILLER_36_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15865_ _13511_/X _15865_/B _15865_/C VGND VGND VPWR VPWR _15866_/C sky130_fd_sc_hd__and3_4
XANTENNA__20583__A2 _20582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21780__B2 _21737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17604_ _18587_/B VGND VGND VPWR VPWR _17619_/A sky130_fd_sc_hd__inv_2
XANTENNA__15931__A _11872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14816_ _14816_/A _14812_/X _14815_/X VGND VGND VPWR VPWR _14817_/C sky130_fd_sc_hd__or3_4
X_18584_ _17858_/X _17295_/X _18579_/X _18582_/X _18583_/X VGND VGND VPWR VPWR _18585_/B
+ sky130_fd_sc_hd__a32o_4
X_15796_ _15823_/A _15796_/B _15796_/C VGND VGND VPWR VPWR _15797_/C sky130_fd_sc_hd__and3_4
XFILLER_75_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17535_ _17535_/A VGND VGND VPWR VPWR _17535_/Y sky130_fd_sc_hd__inv_2
X_11959_ _13428_/A VGND VGND VPWR VPWR _11959_/X sky130_fd_sc_hd__buf_2
X_14747_ _15037_/A _14803_/B VGND VGND VPWR VPWR _14747_/X sky130_fd_sc_hd__or2_4
XANTENNA__20268__B _20494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13451__A _13447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_10_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14678_ _14397_/A _14678_/B _14677_/X VGND VGND VPWR VPWR _14678_/X sky130_fd_sc_hd__or3_4
X_17466_ _12559_/X VGND VGND VPWR VPWR _17466_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19205_ _19205_/A _19205_/B VGND VGND VPWR VPWR _19206_/B sky130_fd_sc_hd__and2_4
XFILLER_60_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13629_ _13645_/A VGND VGND VPWR VPWR _13630_/A sky130_fd_sc_hd__buf_2
X_16417_ _16397_/X _16417_/B VGND VGND VPWR VPWR _16418_/C sky130_fd_sc_hd__or2_4
XFILLER_20_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17858__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17397_ _17178_/X _17396_/Y VGND VGND VPWR VPWR _17397_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_5_5_0_HCLK_A clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16762__A _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19136_ _24315_/Q _19135_/X VGND VGND VPWR VPWR _19136_/X sky130_fd_sc_hd__and2_4
XFILLER_9_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16348_ _16188_/A _16280_/B VGND VGND VPWR VPWR _16348_/X sky130_fd_sc_hd__or2_4
XFILLER_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20284__A _20212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18161__B1 _18160_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16279_ _16243_/X _16279_/B VGND VGND VPWR VPWR _16279_/X sky130_fd_sc_hd__or2_4
X_19067_ _19065_/Y _19066_/Y _11513_/B VGND VGND VPWR VPWR _19067_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24301__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14282__A _14322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18018_ _24135_/Q _18017_/Y _17894_/D VGND VGND VPWR VPWR _18018_/X sky130_fd_sc_hd__o21a_4
XFILLER_12_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21599__B2 _21595_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20271__A1 _19953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19969_ _19968_/X VGND VGND VPWR VPWR _19969_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13626__A _13659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22012__A2 _22009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19413__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22980_ _22980_/A VGND VGND VPWR VPWR _23004_/B sky130_fd_sc_hd__buf_2
XANTENNA__12530__A _15032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16002__A _16002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21931_ _21938_/A VGND VGND VPWR VPWR _21931_/X sky130_fd_sc_hd__buf_2
XFILLER_83_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21771__B2 _21766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15841__A _13041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19313__A _19313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21862_ _21861_/X _21853_/X _23584_/Q _21787_/X VGND VGND VPWR VPWR _23584_/D sky130_fd_sc_hd__o22a_4
XFILLER_93_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23601_ _23473_/CLK _23601_/D VGND VGND VPWR VPWR _13174_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_3_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20813_ _20813_/A VGND VGND VPWR VPWR _20813_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15560__B _15560_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21793_ _21817_/A VGND VGND VPWR VPWR _21793_/X sky130_fd_sc_hd__buf_2
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21523__B2 _21515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23532_ _23794_/CLK _21948_/X VGND VGND VPWR VPWR _15410_/B sky130_fd_sc_hd__dfxtp_4
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20744_ _20673_/X _20730_/Y _20742_/X _20743_/Y _20692_/X VGND VGND VPWR VPWR _20744_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23463_ _23368_/CLK _23463_/D VGND VGND VPWR VPWR _23463_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20675_ _20699_/B VGND VGND VPWR VPWR _20675_/X sky130_fd_sc_hd__buf_2
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16672__A _16630_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22414_ _22413_/X _22404_/X _12758_/B _22411_/X VGND VGND VPWR VPWR _22414_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23394_ _24066_/CLK _23394_/D VGND VGND VPWR VPWR _15293_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16391__B _16391_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15288__A _14146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22345_ _22083_/X _22340_/X _16391_/B _22344_/X VGND VGND VPWR VPWR _23290_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12705__A _12705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21039__B1 _15818_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_30_0_HCLK clkbuf_7_30_0_HCLK/A VGND VGND VPWR VPWR _23073_/CLK sky130_fd_sc_hd__clkbuf_1
X_22276_ _22269_/A VGND VGND VPWR VPWR _22276_/X sky130_fd_sc_hd__buf_2
XFILLER_69_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20922__A HRDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_93_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR _23320_/CLK sky130_fd_sc_hd__clkbuf_1
X_24015_ _23983_/CLK _24015_/D VGND VGND VPWR VPWR _13513_/B sky130_fd_sc_hd__dfxtp_4
X_21227_ _21797_/A VGND VGND VPWR VPWR _21227_/X sky130_fd_sc_hd__buf_2
XFILLER_78_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21158_ _20958_/X _21154_/X _15210_/B _21115_/X VGND VGND VPWR VPWR _21158_/X sky130_fd_sc_hd__o22a_4
XFILLER_77_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20109_ _19934_/X _20108_/X _19380_/X _16964_/A VGND VGND VPWR VPWR _24113_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13536__A _13494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13980_ _13953_/A _23082_/Q VGND VGND VPWR VPWR _13982_/B sky130_fd_sc_hd__or2_4
XANTENNA__22003__A2 _22002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21089_ _21075_/A VGND VGND VPWR VPWR _21089_/X sky130_fd_sc_hd__buf_2
XFILLER_115_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14492__A2 _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12931_ _12655_/A _12927_/X _12930_/X VGND VGND VPWR VPWR _12931_/X sky130_fd_sc_hd__or3_4
XFILLER_74_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20565__A2 _20564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12862_ _12862_/A VGND VGND VPWR VPWR _12890_/A sky130_fd_sc_hd__buf_2
X_15650_ _15650_/A VGND VGND VPWR VPWR _15650_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11813_ _11818_/A _11813_/B VGND VGND VPWR VPWR _11815_/B sky130_fd_sc_hd__or2_4
X_14601_ _15006_/A _14674_/B VGND VGND VPWR VPWR _14601_/X sky130_fd_sc_hd__or2_4
X_15581_ _11977_/X _15558_/X _15565_/X _15572_/X _15580_/X VGND VGND VPWR VPWR _15581_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15470__B _23916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12793_ _12802_/A _23156_/Q VGND VGND VPWR VPWR _12793_/X sky130_fd_sc_hd__or2_4
XFILLER_37_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14367__A _14367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__A _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22711__B1 _15176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14500_/X _14532_/B VGND VGND VPWR VPWR _14532_/X sky130_fd_sc_hd__or2_4
X_17320_ _18655_/B _18658_/A VGND VGND VPWR VPWR _18662_/A sky130_fd_sc_hd__or2_4
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _13422_/A VGND VGND VPWR VPWR _16229_/A sky130_fd_sc_hd__buf_2
XFILLER_72_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19877__B _19877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14463_/A _14533_/B VGND VGND VPWR VPWR _14464_/C sky130_fd_sc_hd__or2_4
X_17251_ _17251_/A VGND VGND VPWR VPWR _17811_/A sky130_fd_sc_hd__buf_2
XFILLER_30_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _16180_/A VGND VGND VPWR VPWR _11675_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _13388_/A _13414_/B _13414_/C VGND VGND VPWR VPWR _13415_/C sky130_fd_sc_hd__and3_4
X_16202_ _16202_/A _23959_/Q VGND VGND VPWR VPWR _16203_/C sky130_fd_sc_hd__or2_4
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17182_ _17181_/X VGND VGND VPWR VPWR _17182_/Y sky130_fd_sc_hd__inv_2
X_14394_ _13844_/A VGND VGND VPWR VPWR _15618_/A sky130_fd_sc_hd__buf_2
XFILLER_70_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16133_ _16109_/A _16131_/X _16133_/C VGND VGND VPWR VPWR _16137_/B sky130_fd_sc_hd__and3_4
X_13345_ _12859_/A _13343_/X _13344_/X VGND VGND VPWR VPWR _13346_/C sky130_fd_sc_hd__and3_4
XANTENNA__15198__A _14215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19893__A _18752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16064_ _16064_/A _23704_/Q VGND VGND VPWR VPWR _16066_/B sky130_fd_sc_hd__or2_4
X_13276_ _13136_/X VGND VGND VPWR VPWR _13276_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21928__A _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15015_ _15015_/A _15015_/B _15015_/C VGND VGND VPWR VPWR _15015_/X sky130_fd_sc_hd__and3_4
X_12227_ _13054_/A VGND VGND VPWR VPWR _13017_/A sky130_fd_sc_hd__buf_2
XANTENNA__22242__A2 _22236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19823_ _19823_/A VGND VGND VPWR VPWR _21581_/A sky130_fd_sc_hd__buf_2
XFILLER_97_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12158_ _11746_/X _12154_/X _12157_/X VGND VGND VPWR VPWR _12158_/X sky130_fd_sc_hd__or3_4
XFILLER_69_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20270__C _20269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13446__A _13442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19754_ _19754_/A _19765_/B VGND VGND VPWR VPWR _19754_/X sky130_fd_sc_hd__and2_4
X_12089_ _12051_/X _12089_/B _12089_/C VGND VGND VPWR VPWR _12089_/X sky130_fd_sc_hd__or3_4
X_16966_ _16966_/A VGND VGND VPWR VPWR _17720_/A sky130_fd_sc_hd__inv_2
XANTENNA__12350__A _12350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18705_ _17117_/X VGND VGND VPWR VPWR _18705_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21202__B1 _14302_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15917_ _14267_/X _16841_/A VGND VGND VPWR VPWR _15917_/Y sky130_fd_sc_hd__nor2_4
X_19685_ _19661_/A VGND VGND VPWR VPWR _19873_/B sky130_fd_sc_hd__buf_2
XFILLER_37_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16897_ _16897_/A _12188_/Y VGND VGND VPWR VPWR _16897_/X sky130_fd_sc_hd__or2_4
XANTENNA__21753__B2 _21752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15661__A _12688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18636_ _18189_/A _18039_/Y VGND VGND VPWR VPWR _18636_/X sky130_fd_sc_hd__and2_4
X_15848_ _13546_/X _15848_/B VGND VGND VPWR VPWR _15848_/X sky130_fd_sc_hd__or2_4
XFILLER_92_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20279__A _20279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18567_ _18137_/A _18567_/B VGND VGND VPWR VPWR _18567_/X sky130_fd_sc_hd__and2_4
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15779_ _15778_/X VGND VGND VPWR VPWR _15780_/B sky130_fd_sc_hd__buf_2
XFILLER_55_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14277__A _13670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23171__CLK _23107_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21505__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24297__CLK _24299_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13181__A _15696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17518_ _18332_/A _17516_/Y _17517_/X VGND VGND VPWR VPWR _17518_/X sky130_fd_sc_hd__o21a_4
X_18498_ _18498_/A VGND VGND VPWR VPWR _18714_/A sky130_fd_sc_hd__inv_2
XFILLER_75_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17449_ _16569_/A _17467_/B VGND VGND VPWR VPWR _17449_/X sky130_fd_sc_hd__and2_4
XFILLER_21_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20460_ _20444_/X _20446_/Y _20457_/X _20458_/Y _20459_/X VGND VGND VPWR VPWR _20461_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_105_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21808__A2 _21805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19119_ _24298_/Q _19181_/A VGND VGND VPWR VPWR _19120_/B sky130_fd_sc_hd__and2_4
XFILLER_118_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17488__A2 _17013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20391_ _20484_/A _20391_/B VGND VGND VPWR VPWR _20391_/X sky130_fd_sc_hd__or2_4
XANTENNA__12525__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22481__A2 _22479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22130_ _22129_/X _22125_/X _13875_/B _22120_/X VGND VGND VPWR VPWR _23431_/D sky130_fd_sc_hd__o22a_4
XFILLER_106_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_17_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22061_ _21855_/X _22059_/X _14769_/B _22056_/X VGND VGND VPWR VPWR _22061_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15836__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14740__A _12883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19352__A2_N _18654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21012_ _21027_/A VGND VGND VPWR VPWR _21012_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15555__B _23595_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17660__A2 _17653_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22669__A _22668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18866__B _18866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22963_ _18430_/X _22950_/X VGND VGND VPWR VPWR _22963_/X sky130_fd_sc_hd__or2_4
XFILLER_114_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16667__A _16640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21744__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21914_ _21863_/X _21887_/A _23551_/Q _21869_/X VGND VGND VPWR VPWR _21914_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15571__A _15571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22894_ _22886_/X _18701_/X _22887_/X _22893_/X VGND VGND VPWR VPWR _22895_/A sky130_fd_sc_hd__a211o_4
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20952__C1 _20951_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21845_ _20819_/A VGND VGND VPWR VPWR _21845_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21776_ _21740_/A VGND VGND VPWR VPWR _21776_/X sky130_fd_sc_hd__buf_2
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12419__B _12316_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23515_ _23515_/CLK _23515_/D VGND VGND VPWR VPWR _23515_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20727_ HRDATA[11] _20821_/B VGND VGND VPWR VPWR _20727_/X sky130_fd_sc_hd__or2_4
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23446_ _23313_/CLK _23446_/D VGND VGND VPWR VPWR _12276_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20658_ _20654_/X _20655_/Y _20657_/X _19034_/Y _20473_/X VGND VGND VPWR VPWR _20658_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23377_ _23313_/CLK _23377_/D VGND VGND VPWR VPWR _13181_/B sky130_fd_sc_hd__dfxtp_4
X_20589_ _24208_/Q _20512_/X _20588_/Y VGND VGND VPWR VPWR _20590_/A sky130_fd_sc_hd__o21a_4
XANTENNA__12435__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13130_ _13130_/A _13046_/B VGND VGND VPWR VPWR _13131_/C sky130_fd_sc_hd__or2_4
XFILLER_87_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20483__A1 _24245_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22328_ _15269_/B VGND VGND VPWR VPWR _22328_/X sky130_fd_sc_hd__buf_2
XANTENNA__21748__A _21755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13061_ _13087_/A VGND VGND VPWR VPWR _13096_/A sky130_fd_sc_hd__buf_2
XANTENNA__15746__A _12957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22259_ _22075_/X _22258_/X _12123_/B _22255_/X VGND VGND VPWR VPWR _23357_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22224__A2 _22222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18122__A _17568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12012_ _16143_/A VGND VGND VPWR VPWR _12020_/A sky130_fd_sc_hd__buf_2
XFILLER_117_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15465__B _15465_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21983__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16820_ _12188_/Y _16819_/X _12187_/X VGND VGND VPWR VPWR _16820_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17961__A _17871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13266__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22579__A _22586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16751_ _16773_/A _23739_/Q VGND VGND VPWR VPWR _16751_/X sky130_fd_sc_hd__or2_4
XANTENNA__17680__B _17479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13963_ _12472_/X _24042_/Q VGND VGND VPWR VPWR _13964_/C sky130_fd_sc_hd__or2_4
XANTENNA__20538__A2 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15702_ _15820_/A _15698_/X _15701_/X VGND VGND VPWR VPWR _15702_/X sky130_fd_sc_hd__or3_4
X_12914_ _12914_/A _12914_/B _12913_/X VGND VGND VPWR VPWR _12914_/X sky130_fd_sc_hd__or3_4
X_19470_ _19458_/A _19469_/X HRDATA[10] _19462_/A VGND VGND VPWR VPWR _19471_/A sky130_fd_sc_hd__o22a_4
X_13894_ _13878_/A _13814_/B VGND VGND VPWR VPWR _13896_/B sky130_fd_sc_hd__or2_4
X_16682_ _16682_/A _16681_/Y VGND VGND VPWR VPWR _16682_/X sky130_fd_sc_hd__or2_4
X_18421_ _18421_/A _17380_/A VGND VGND VPWR VPWR _18421_/X sky130_fd_sc_hd__and2_4
X_12845_ _12842_/X _12845_/B VGND VGND VPWR VPWR _12845_/X sky130_fd_sc_hd__or2_4
X_15633_ _15633_/A _15577_/B VGND VGND VPWR VPWR _15634_/C sky130_fd_sc_hd__or2_4
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13713__B _13713_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19888__A _19933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18352_ _17699_/X _18352_/B VGND VGND VPWR VPWR _18383_/B sky130_fd_sc_hd__or2_4
X_12776_ _12421_/A VGND VGND VPWR VPWR _13087_/A sky130_fd_sc_hd__buf_2
X_15564_ _11911_/A _15562_/X _15563_/X VGND VGND VPWR VPWR _15565_/C sky130_fd_sc_hd__and3_4
XFILLER_15_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17297_/X _17309_/B VGND VGND VPWR VPWR _17306_/A sky130_fd_sc_hd__and2_4
XFILLER_42_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22160__B2 _22155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _12830_/A VGND VGND VPWR VPWR _11727_/X sky130_fd_sc_hd__buf_2
X_14515_ _14500_/X _14453_/B VGND VGND VPWR VPWR _14515_/X sky130_fd_sc_hd__or2_4
XFILLER_72_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15495_/A _15495_/B _15494_/X VGND VGND VPWR VPWR _15499_/B sky130_fd_sc_hd__and3_4
X_18283_ _18263_/X _18268_/Y _18273_/X _18281_/X _18282_/Y VGND VGND VPWR VPWR _18283_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14825__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17234_ _17825_/A _17230_/X _17817_/A _17233_/X VGND VGND VPWR VPWR _17234_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_35_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _11657_/X VGND VGND VPWR VPWR _11658_/X sky130_fd_sc_hd__buf_2
X_14446_ _12878_/A _14523_/B VGND VGND VPWR VPWR _14446_/X sky130_fd_sc_hd__or2_4
XFILLER_70_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _15604_/A _14377_/B _14377_/C VGND VGND VPWR VPWR _14388_/B sky130_fd_sc_hd__or3_4
X_17165_ _17164_/X VGND VGND VPWR VPWR _17165_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18667__A1 _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11589_ _17412_/A VGND VGND VPWR VPWR _17028_/A sky130_fd_sc_hd__buf_2
XFILLER_7_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22463__A2 _22416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20474__A1 _20425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13328_ _13300_/A _13328_/B VGND VGND VPWR VPWR _13328_/X sky130_fd_sc_hd__or2_4
X_16116_ _16087_/X _16116_/B _16116_/C VGND VGND VPWR VPWR _16121_/B sky130_fd_sc_hd__and3_4
XANTENNA__20474__B2 _20473_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17096_ _17081_/X _18180_/A _17096_/C _17095_/X VGND VGND VPWR VPWR _17097_/A sky130_fd_sc_hd__or4_4
XANTENNA__20562__A _20301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12064__B _23677_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15656__A _12286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13259_ _13211_/A _13255_/X _13258_/X VGND VGND VPWR VPWR _13259_/X sky130_fd_sc_hd__or3_4
X_16047_ _16047_/A _23960_/Q VGND VGND VPWR VPWR _16047_/X sky130_fd_sc_hd__or2_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14560__A _13747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19806_ _19612_/A _19759_/B _19806_/C _19805_/Y VGND VGND VPWR VPWR _19806_/X sky130_fd_sc_hd__or4_4
XFILLER_69_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17871__A _17871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23537__CLK _23155_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17998_ _18160_/A VGND VGND VPWR VPWR _17998_/X sky130_fd_sc_hd__buf_2
XFILLER_84_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19737_ _19724_/X _19733_/X _19534_/X _19736_/X VGND VGND VPWR VPWR _19737_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19919__B2 _20895_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16949_ _18234_/A VGND VGND VPWR VPWR _17673_/A sky130_fd_sc_hd__inv_2
X_19668_ _19800_/B _19624_/A VGND VGND VPWR VPWR _19668_/X sky130_fd_sc_hd__or2_4
XFILLER_93_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_8_0_HCLK clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18619_ _17103_/X _18078_/Y _17240_/X _18618_/X VGND VGND VPWR VPWR _18619_/X sky130_fd_sc_hd__a211o_4
XFILLER_111_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19599_ _19561_/A _19599_/B VGND VGND VPWR VPWR _19600_/B sky130_fd_sc_hd__or2_4
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21630_ _21574_/X _21626_/X _23713_/Q _21595_/A VGND VGND VPWR VPWR _21630_/X sky130_fd_sc_hd__o22a_4
XFILLER_90_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17158__A1 _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21561_ _21560_/X _21556_/X _23751_/Q _21551_/X VGND VGND VPWR VPWR _21561_/X sky130_fd_sc_hd__o22a_4
XFILLER_60_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18207__A _18266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23300_ _23363_/CLK _22326_/X VGND VGND VPWR VPWR _14682_/B sky130_fd_sc_hd__dfxtp_4
X_20512_ _20512_/A VGND VGND VPWR VPWR _20512_/X sky130_fd_sc_hd__buf_2
X_24280_ _24344_/CLK _24280_/D HRESETn VGND VGND VPWR VPWR _24280_/Q sky130_fd_sc_hd__dfrtp_4
X_21492_ _21282_/X _21491_/X _14632_/B _21488_/X VGND VGND VPWR VPWR _23780_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18654__A1_N _17742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23231_ _23889_/CLK _23231_/D VGND VGND VPWR VPWR _15052_/B sky130_fd_sc_hd__dfxtp_4
X_20443_ _20396_/X _20442_/X _24087_/Q _20374_/X VGND VGND VPWR VPWR _24087_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12255__A _12709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23162_ _23313_/CLK _23162_/D VGND VGND VPWR VPWR _16407_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21568__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20465__B2 _20374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20374_ _20202_/X VGND VGND VPWR VPWR _20374_/X sky130_fd_sc_hd__buf_2
XFILLER_101_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22113_ _22101_/A VGND VGND VPWR VPWR _22113_/X sky130_fd_sc_hd__buf_2
XANTENNA__19870__A3 _19869_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23093_ _23315_/CLK _23093_/D VGND VGND VPWR VPWR _12657_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17881__A2 _17775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20191__B _22017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22044_ _21826_/X _22038_/X _23471_/Q _22042_/X VGND VGND VPWR VPWR _22044_/X sky130_fd_sc_hd__o22a_4
XFILLER_114_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18877__A _18877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21965__B2 _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17781__A _18205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18830__A1 _17164_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22399__A _22386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23995_ _24092_/CLK _23995_/D VGND VGND VPWR VPWR _23995_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21717__B2 _21716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13814__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22946_ _22952_/A _22946_/B _22946_/C VGND VGND VPWR VPWR _22946_/X sky130_fd_sc_hd__and3_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21193__A2 _21190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22877_ _12116_/Y _22863_/X _19887_/X _22876_/X VGND VGND VPWR VPWR _22878_/B sky130_fd_sc_hd__o22a_4
XANTENNA__24404__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12630_ _12412_/A VGND VGND VPWR VPWR _13737_/A sky130_fd_sc_hd__buf_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13958__A1 _14172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21828_ _21543_/A VGND VGND VPWR VPWR _21828_/X sky130_fd_sc_hd__buf_2
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20647__A HRDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22142__B2 _22132_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _13770_/A VGND VGND VPWR VPWR _13083_/A sky130_fd_sc_hd__buf_2
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21759_ _21752_/A VGND VGND VPWR VPWR _21759_/X sky130_fd_sc_hd__buf_2
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18897__A1 _17194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14645__A _15105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11512_ _19065_/A _11512_/B VGND VGND VPWR VPWR _11513_/B sky130_fd_sc_hd__or2_4
X_14300_ _13597_/X _14274_/X _14281_/X _14291_/X _14299_/X VGND VGND VPWR VPWR _14300_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17021__A _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15280_ _11976_/A _15279_/X VGND VGND VPWR VPWR _15280_/X sky130_fd_sc_hd__and2_4
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12492_ _12905_/A _12628_/B VGND VGND VPWR VPWR _12493_/C sky130_fd_sc_hd__or2_4
X_24478_ _24229_/CLK _24478_/D HRESETn VGND VGND VPWR VPWR _19956_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14231_ _14252_/A _24041_/Q VGND VGND VPWR VPWR _14231_/X sky130_fd_sc_hd__or2_4
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23429_ _23973_/CLK _23429_/D VGND VGND VPWR VPWR _14520_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17956__A _17090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22445__A2 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18649__B2 _18648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12165__A _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24344__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14162_ _14737_/A _14162_/B _14161_/X VGND VGND VPWR VPWR _14163_/C sky130_fd_sc_hd__and3_4
XANTENNA__21653__B1 _12660_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13113_ _13096_/A _13111_/X _13113_/C VGND VGND VPWR VPWR _13113_/X sky130_fd_sc_hd__and3_4
XANTENNA__15476__A _12613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14093_ _11879_/A _24009_/Q VGND VGND VPWR VPWR _14093_/X sky130_fd_sc_hd__or2_4
X_18970_ _18956_/X _18969_/X _18956_/X _24344_/Q VGND VGND VPWR VPWR _18970_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_63_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13044_ _13017_/A _13044_/B _13043_/X VGND VGND VPWR VPWR _13048_/B sky130_fd_sc_hd__and3_4
X_17921_ _17921_/A VGND VGND VPWR VPWR _17921_/X sky130_fd_sc_hd__buf_2
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17852_ _17796_/X _17834_/X _17836_/X _17851_/X VGND VGND VPWR VPWR _17853_/A sky130_fd_sc_hd__o22a_4
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16803_ _16803_/A _23483_/Q VGND VGND VPWR VPWR _16805_/B sky130_fd_sc_hd__or2_4
XFILLER_43_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17783_ _17782_/Y VGND VGND VPWR VPWR _18442_/A sky130_fd_sc_hd__buf_2
XFILLER_94_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14995_ _14995_/A _14995_/B _14995_/C VGND VGND VPWR VPWR _14995_/X sky130_fd_sc_hd__or3_4
XANTENNA__21708__A1 _21536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21708__B2 _21702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19522_ _19866_/B _19521_/X VGND VGND VPWR VPWR _19522_/X sky130_fd_sc_hd__or2_4
XANTENNA__13724__A _15494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16734_ _11993_/A _23099_/Q VGND VGND VPWR VPWR _16736_/B sky130_fd_sc_hd__or2_4
X_13946_ _12509_/A _23530_/Q VGND VGND VPWR VPWR _13947_/C sky130_fd_sc_hd__or2_4
XFILLER_81_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21184__A2 _21183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22381__B2 _22344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19453_ _20224_/B _19545_/A _19712_/A HRDATA[15] VGND VGND VPWR VPWR _19453_/Y sky130_fd_sc_hd__a22oi_4
X_16665_ _16630_/X _23708_/Q VGND VGND VPWR VPWR _16665_/X sky130_fd_sc_hd__or2_4
XANTENNA__24145__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13877_ _13893_/A _13869_/X _13877_/C VGND VGND VPWR VPWR _13885_/B sky130_fd_sc_hd__or3_4
XFILLER_35_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18404_ _18216_/X _17377_/X _18397_/X _18398_/X _18403_/Y VGND VGND VPWR VPWR _18404_/X
+ sky130_fd_sc_hd__a32o_4
X_15616_ _15616_/A _15614_/X _15615_/X VGND VGND VPWR VPWR _15616_/X sky130_fd_sc_hd__and3_4
X_12828_ _12828_/A VGND VGND VPWR VPWR _12829_/A sky130_fd_sc_hd__buf_2
X_19384_ _19317_/A VGND VGND VPWR VPWR _19385_/A sky130_fd_sc_hd__buf_2
XFILLER_50_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16596_ _16596_/A VGND VGND VPWR VPWR _16596_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22133__B2 _22132_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12059__B _12132_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18335_ _18314_/X _18316_/X _18202_/X _18334_/X VGND VGND VPWR VPWR _18335_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15547_ _15574_/A _23435_/Q VGND VGND VPWR VPWR _15547_/X sky130_fd_sc_hd__or2_4
XANTENNA__18888__A1 _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12759_ _12605_/A VGND VGND VPWR VPWR _13065_/A sky130_fd_sc_hd__buf_2
XANTENNA__22684__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20695__A1 _24204_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18266_ _18266_/A _17500_/Y VGND VGND VPWR VPWR _18267_/D sky130_fd_sc_hd__and2_4
X_15478_ _12585_/A _15407_/B VGND VGND VPWR VPWR _15478_/X sky130_fd_sc_hd__or2_4
XFILLER_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24335__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17217_ _17132_/Y _17173_/X _15251_/X _17133_/X VGND VGND VPWR VPWR _17217_/X sky130_fd_sc_hd__o22a_4
X_14429_ _14336_/X _14429_/B VGND VGND VPWR VPWR _14430_/B sky130_fd_sc_hd__and2_4
X_18197_ _18129_/X _18196_/X _24469_/Q _18129_/X VGND VGND VPWR VPWR _24469_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12075__A _11994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22436__A2 _22428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21644__B1 _23707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17148_ _17147_/X VGND VGND VPWR VPWR _17148_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20998__A2 _20989_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17079_ _17079_/A _17224_/A _18728_/B VGND VGND VPWR VPWR _18025_/A sky130_fd_sc_hd__or3_4
XFILLER_116_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14290__A _11911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12803__A _12803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20090_ _20090_/A _20090_/B _20089_/X _20090_/D VGND VGND VPWR VPWR _20091_/A sky130_fd_sc_hd__or4_4
XANTENNA__18697__A _18697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21947__B2 _21942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22800_ _22792_/X _22800_/B VGND VGND VPWR VPWR HWDATA[8] sky130_fd_sc_hd__nor2_4
XANTENNA__13634__A _15436_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23780_ _23907_/CLK _23780_/D VGND VGND VPWR VPWR _14632_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20992_ _20403_/A _20991_/X _24255_/Q _20497_/A VGND VGND VPWR VPWR _20992_/X sky130_fd_sc_hd__o22a_4
XFILLER_65_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21175__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22731_ _22731_/A VGND VGND VPWR VPWR _22756_/A sky130_fd_sc_hd__inv_2
XFILLER_0_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13353__B _13282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19321__A _19328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22662_ _22460_/X _22657_/X _14962_/B _22626_/A VGND VGND VPWR VPWR _22662_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24401_ _23326_/CLK _24401_/D HRESETn VGND VGND VPWR VPWR _24401_/Q sky130_fd_sc_hd__dfrtp_4
X_21613_ _21543_/X _21612_/X _15656_/B _21609_/X VGND VGND VPWR VPWR _23726_/D sky130_fd_sc_hd__o22a_4
XFILLER_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18879__A1 _11837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22593_ _22586_/A VGND VGND VPWR VPWR _22593_/X sky130_fd_sc_hd__buf_2
XANTENNA__22675__A2 _22672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24332_ _23260_/CLK _24332_/D HRESETn VGND VGND VPWR VPWR _24332_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_90_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21544_ _21532_/A VGND VGND VPWR VPWR _21544_/X sky130_fd_sc_hd__buf_2
XANTENNA__21883__B1 _12271_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24263_ _24305_/CLK _19282_/X HRESETn VGND VGND VPWR VPWR _19212_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17776__A _18203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21475_ _21253_/X _21470_/X _13341_/B _21474_/X VGND VGND VPWR VPWR _21475_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16680__A _16596_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23214_ _23564_/CLK _23214_/D VGND VGND VPWR VPWR _15699_/B sky130_fd_sc_hd__dfxtp_4
X_20426_ _20426_/A _20519_/B VGND VGND VPWR VPWR _20426_/Y sky130_fd_sc_hd__nand2_4
X_24194_ _24199_/CLK _19409_/X HRESETn VGND VGND VPWR VPWR _24194_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23145_ _23145_/CLK _23145_/D VGND VGND VPWR VPWR _23145_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13809__A _15424_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15296__A _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20357_ _20280_/X _20356_/X _24091_/Q _20203_/X VGND VGND VPWR VPWR _20357_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12713__A _12713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23076_ _23812_/CLK _22708_/X VGND VGND VPWR VPWR _14703_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12679__A1 _12559_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20288_ _20515_/A VGND VGND VPWR VPWR _20288_/X sky130_fd_sc_hd__buf_2
XANTENNA__12432__B _12429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22027_ _21797_/X _22024_/X _23483_/Q _22021_/X VGND VGND VPWR VPWR _22027_/X sky130_fd_sc_hd__o22a_4
XFILLER_49_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13800_ _13800_/A _13798_/X _13800_/C VGND VGND VPWR VPWR _13800_/X sky130_fd_sc_hd__and3_4
XANTENNA__13544__A _13511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11992_ _11982_/X VGND VGND VPWR VPWR _11992_/X sky130_fd_sc_hd__buf_2
X_14780_ _12509_/A _14780_/B VGND VGND VPWR VPWR _14781_/C sky130_fd_sc_hd__or2_4
X_23978_ _23978_/CLK _23978_/D VGND VGND VPWR VPWR _23978_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22363__B2 _22358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13731_ _13731_/A _13725_/X _13730_/X VGND VGND VPWR VPWR _13731_/X sky130_fd_sc_hd__or3_4
XFILLER_75_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22929_ _22952_/A _22927_/X _22929_/C VGND VGND VPWR VPWR _22929_/X sky130_fd_sc_hd__and3_4
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16450_ _16464_/A _16383_/B VGND VGND VPWR VPWR _16453_/B sky130_fd_sc_hd__or2_4
X_13662_ _15430_/A _13662_/B VGND VGND VPWR VPWR _13662_/X sky130_fd_sc_hd__or2_4
X_15401_ _12450_/A _15401_/B _15401_/C VGND VGND VPWR VPWR _15401_/X sky130_fd_sc_hd__and3_4
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ _12613_/A VGND VGND VPWR VPWR _12948_/A sky130_fd_sc_hd__buf_2
X_13593_ _13590_/X _13593_/B VGND VGND VPWR VPWR _13593_/X sky130_fd_sc_hd__or2_4
X_16381_ _15997_/A _16381_/B VGND VGND VPWR VPWR _16382_/C sky130_fd_sc_hd__or2_4
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18120_ _18107_/X _18115_/Y _17240_/X _18119_/Y VGND VGND VPWR VPWR _18120_/X sky130_fd_sc_hd__a211o_4
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18334__A3 _18328_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12544_ _12540_/A _12542_/X _12544_/C VGND VGND VPWR VPWR _12549_/B sky130_fd_sc_hd__and3_4
X_15332_ _15332_/A _15273_/B VGND VGND VPWR VPWR _15332_/X sky130_fd_sc_hd__or2_4
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12607__B _12607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18051_ _17950_/X _18020_/Y _18022_/X _18050_/X VGND VGND VPWR VPWR _18051_/X sky130_fd_sc_hd__o22a_4
X_12475_ _12475_/A VGND VGND VPWR VPWR _13020_/A sky130_fd_sc_hd__buf_2
X_15263_ _14143_/A _15263_/B VGND VGND VPWR VPWR _15263_/X sky130_fd_sc_hd__or2_4
XANTENNA__16590__A _11903_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17002_ _17002_/A _17001_/X VGND VGND VPWR VPWR _17003_/A sky130_fd_sc_hd__and2_4
XANTENNA__20429__A1 _20425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14214_ _14205_/A _23977_/Q VGND VGND VPWR VPWR _14215_/C sky130_fd_sc_hd__or2_4
XANTENNA__20429__B2 _20253_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15194_ _11709_/A _23745_/Q VGND VGND VPWR VPWR _15195_/C sky130_fd_sc_hd__or2_4
X_14145_ _14145_/A _14145_/B _14144_/X VGND VGND VPWR VPWR _14145_/X sky130_fd_sc_hd__or3_4
XANTENNA__21001__A _21001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13719__A _15494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12623__A _12622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14076_ _14075_/X VGND VGND VPWR VPWR _14076_/Y sky130_fd_sc_hd__inv_2
X_18953_ _24346_/Q _11530_/X _18924_/Y VGND VGND VPWR VPWR _18953_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_4_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21929__B2 _21928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13027_ _12922_/A _13004_/X _13011_/X _13018_/X _13026_/X VGND VGND VPWR VPWR _13027_/X
+ sky130_fd_sc_hd__a32o_4
X_17904_ _18390_/A _17904_/B _17902_/X _17904_/D VGND VGND VPWR VPWR _17905_/A sky130_fd_sc_hd__or4_4
XANTENNA__15934__A _15956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18884_ _18891_/A VGND VGND VPWR VPWR _18884_/X sky130_fd_sc_hd__buf_2
XFILLER_45_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24397__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20601__A1 _20518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16749__B _16749_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17835_ _17256_/A VGND VGND VPWR VPWR _17836_/A sky130_fd_sc_hd__buf_2
XANTENNA__20601__B2 _20525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15653__B _15715_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13454__A _12865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17766_ _17766_/A _17274_/Y VGND VGND VPWR VPWR _17946_/A sky130_fd_sc_hd__or2_4
X_14978_ _15074_/A _14903_/B VGND VGND VPWR VPWR _14978_/X sky130_fd_sc_hd__or2_4
XANTENNA__21157__A2 _21154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19505_ _19598_/A VGND VGND VPWR VPWR _19744_/A sky130_fd_sc_hd__inv_2
XANTENNA__14269__B _14269_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16717_ _16698_/A _24059_/Q VGND VGND VPWR VPWR _16717_/X sky130_fd_sc_hd__or2_4
X_13929_ _11611_/A VGND VGND VPWR VPWR _15036_/A sky130_fd_sc_hd__buf_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17697_ _17697_/A VGND VGND VPWR VPWR _17698_/A sky130_fd_sc_hd__inv_2
XFILLER_39_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16765__A _16747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19436_ _24143_/Q _19432_/X HRDATA[17] _19435_/X VGND VGND VPWR VPWR _19436_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_90_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16648_ _16610_/A _23964_/Q VGND VGND VPWR VPWR _16649_/C sky130_fd_sc_hd__or2_4
XFILLER_91_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22106__B2 _22096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19367_ _19370_/A VGND VGND VPWR VPWR _19367_/X sky130_fd_sc_hd__buf_2
X_16579_ _16686_/A _23484_/Q VGND VGND VPWR VPWR _16581_/B sky130_fd_sc_hd__or2_4
X_18318_ _18264_/A _17517_/B VGND VGND VPWR VPWR _18321_/B sky130_fd_sc_hd__and2_4
XFILLER_17_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23725__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11702__A _11702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19298_ _22924_/A VGND VGND VPWR VPWR _23064_/B sky130_fd_sc_hd__buf_2
X_18249_ _18249_/A VGND VGND VPWR VPWR _18249_/X sky130_fd_sc_hd__buf_2
XANTENNA__22409__A2 _22404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21617__B1 _23723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21260_ _21258_/X _21259_/X _15729_/B _21254_/X VGND VGND VPWR VPWR _23918_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15828__B _15828_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23875__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19825__A3 _19822_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20211_ _20195_/D VGND VGND VPWR VPWR _20516_/A sky130_fd_sc_hd__inv_2
XANTENNA__13629__A _13645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21191_ _20637_/X _21190_/X _15748_/B _21187_/X VGND VGND VPWR VPWR _23950_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12533__A _12533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16005__A _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20840__A1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20142_ IRQ[11] VGND VGND VPWR VPWR _20142_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20840__B2 _20839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20750__A _20279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20073_ _12100_/X _12098_/A _18866_/D _11602_/X VGND VGND VPWR VPWR _20073_/X sky130_fd_sc_hd__or4_4
XFILLER_83_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21396__A2 _21369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23901_ _23515_/CLK _21306_/X VGND VGND VPWR VPWR _23901_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15563__B _23403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23832_ _24088_/CLK _23832_/D VGND VGND VPWR VPWR _23832_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21148__A2 _21147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23763_ _23986_/CLK _23763_/D VGND VGND VPWR VPWR _12858_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20975_ _22824_/B _20291_/X _20758_/X _20974_/Y VGND VGND VPWR VPWR _20976_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16675__A _16622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22714_ _19201_/X HREADY VGND VGND VPWR VPWR _22714_/X sky130_fd_sc_hd__and2_4
X_23694_ _23342_/CLK _23694_/D VGND VGND VPWR VPWR _15765_/B sky130_fd_sc_hd__dfxtp_4
X_22645_ _22430_/X _22643_/X _15821_/B _22640_/X VGND VGND VPWR VPWR _22645_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22648__A2 _22643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14195__A _14195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12708__A _12240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11612__A _13966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22576_ _22576_/A VGND VGND VPWR VPWR _22576_/X sky130_fd_sc_hd__buf_2
XFILLER_107_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21320__A2 _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21527_ _21527_/A VGND VGND VPWR VPWR _21527_/X sky130_fd_sc_hd__buf_2
X_24315_ _24290_/CLK _24315_/D HRESETn VGND VGND VPWR VPWR _24315_/Q sky130_fd_sc_hd__dfrtp_4
X_12260_ _15447_/A VGND VGND VPWR VPWR _12260_/X sky130_fd_sc_hd__buf_2
X_24246_ _24216_/CLK _19324_/X HRESETn VGND VGND VPWR VPWR _24246_/Q sky130_fd_sc_hd__dfrtp_4
X_21458_ _21225_/X _21456_/X _23804_/Q _21453_/X VGND VGND VPWR VPWR _23804_/D sky130_fd_sc_hd__o22a_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20409_ _20403_/X _20408_/X _24280_/Q _20327_/X VGND VGND VPWR VPWR _20409_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13539__A _15876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21084__B2 _21079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12191_ _15449_/A VGND VGND VPWR VPWR _15412_/A sky130_fd_sc_hd__buf_2
X_24177_ _23104_/CLK _19750_/Y HRESETn VGND VGND VPWR VPWR _11651_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22732__A1_N SYSTICKCLKDIV[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21389_ _21280_/X _21383_/X _14487_/B _21387_/X VGND VGND VPWR VPWR _23845_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12443__A _12443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23128_ _23313_/CLK _23128_/D VGND VGND VPWR VPWR _15981_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12162__B _12162_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15754__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15950_ _15959_/A VGND VGND VPWR VPWR _15984_/A sky130_fd_sc_hd__buf_2
X_23059_ _19925_/X _19306_/Y _22719_/X _23058_/X VGND VGND VPWR VPWR _23060_/A sky130_fd_sc_hd__a211o_4
XFILLER_118_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22584__A1 _22410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14901_ _14995_/A _14901_/B _14900_/X VGND VGND VPWR VPWR _14901_/X sky130_fd_sc_hd__or3_4
XANTENNA__22584__B2 _22583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15881_ _13529_/X _15881_/B _15880_/X VGND VGND VPWR VPWR _15882_/C sky130_fd_sc_hd__and3_4
XFILLER_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17620_ _18537_/B VGND VGND VPWR VPWR _17621_/D sky130_fd_sc_hd__inv_2
XANTENNA__13274__A _13135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14832_ _14816_/A _14828_/X _14831_/X VGND VGND VPWR VPWR _14832_/X sky130_fd_sc_hd__or3_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21139__A2 _21133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17551_ _18024_/B VGND VGND VPWR VPWR _18047_/A sky130_fd_sc_hd__inv_2
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14763_ _14763_/A _23811_/Q VGND VGND VPWR VPWR _14763_/X sky130_fd_sc_hd__or2_4
X_11975_ _13957_/A VGND VGND VPWR VPWR _11976_/A sky130_fd_sc_hd__buf_2
XFILLER_75_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16502_ _16203_/A _16502_/B _16501_/X VGND VGND VPWR VPWR _16503_/C sky130_fd_sc_hd__and3_4
XANTENNA__17212__B1 _14263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13714_ _13711_/X _13712_/X _13713_/X VGND VGND VPWR VPWR _13714_/X sky130_fd_sc_hd__and3_4
XFILLER_44_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17482_ _17481_/X VGND VGND VPWR VPWR _17484_/A sky130_fd_sc_hd__inv_2
X_14694_ _14397_/A _14690_/X _14693_/X VGND VGND VPWR VPWR _14694_/X sky130_fd_sc_hd__or3_4
XFILLER_16_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19221_ _24272_/Q _19220_/X VGND VGND VPWR VPWR _19263_/A sky130_fd_sc_hd__and2_4
XFILLER_60_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16433_ _16121_/A _16433_/B _16433_/C VGND VGND VPWR VPWR _16433_/X sky130_fd_sc_hd__or3_4
X_13645_ _13645_/A _13729_/B VGND VGND VPWR VPWR _13646_/C sky130_fd_sc_hd__or2_4
XANTENNA__22639__A2 _22636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19896__A _22978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12618__A _15491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19152_ _24312_/Q _19132_/X _19151_/Y VGND VGND VPWR VPWR _19152_/X sky130_fd_sc_hd__o21a_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16364_ _16364_/A _23481_/Q VGND VGND VPWR VPWR _16366_/B sky130_fd_sc_hd__or2_4
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _13575_/X VGND VGND VPWR VPWR _13577_/B sky130_fd_sc_hd__inv_2
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21311__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18103_ _18103_/A VGND VGND VPWR VPWR _18297_/A sky130_fd_sc_hd__buf_2
X_15315_ _14207_/A _15315_/B _15315_/C VGND VGND VPWR VPWR _15321_/B sky130_fd_sc_hd__and3_4
XFILLER_9_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12527_ _12466_/X _12525_/X _12527_/C VGND VGND VPWR VPWR _12528_/C sky130_fd_sc_hd__and3_4
X_19083_ _19083_/A VGND VGND VPWR VPWR _19083_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15929__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16295_ _11872_/X _16293_/X _16294_/X VGND VGND VPWR VPWR _16295_/X sky130_fd_sc_hd__and3_4
XANTENNA__14833__A _11766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18034_ _17244_/X _17198_/Y _17921_/A _17208_/Y VGND VGND VPWR VPWR _18034_/X sky130_fd_sc_hd__o22a_4
X_15246_ _14367_/A _15242_/X _15245_/X VGND VGND VPWR VPWR _15246_/X sky130_fd_sc_hd__or3_4
X_12458_ _12458_/A _12445_/X _12458_/C VGND VGND VPWR VPWR _12458_/X sky130_fd_sc_hd__or3_4
XANTENNA__13449__A _13448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12389_ _15889_/A _12389_/B _12389_/C VGND VGND VPWR VPWR _12390_/C sky130_fd_sc_hd__or3_4
X_15177_ _14165_/A _15177_/B VGND VGND VPWR VPWR _15177_/X sky130_fd_sc_hd__or2_4
XFILLER_119_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11563__A1 _24434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14128_ _14128_/A _14127_/X VGND VGND VPWR VPWR _14128_/X sky130_fd_sc_hd__and2_4
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21666__A _21659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19985_ _19985_/A VGND VGND VPWR VPWR _19985_/X sky130_fd_sc_hd__buf_2
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15664__A _15664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14059_ _11647_/A _23690_/Q VGND VGND VPWR VPWR _14059_/X sky130_fd_sc_hd__or2_4
X_18936_ _18935_/X VGND VGND VPWR VPWR _18971_/A sky130_fd_sc_hd__buf_2
XANTENNA__21378__A2 _21376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22575__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23278__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18867_ _12098_/A _20248_/A _19926_/B VGND VGND VPWR VPWR _18867_/X sky130_fd_sc_hd__or3_4
XANTENNA__19440__A1 _19545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13184__A _15695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17818_ _17817_/X VGND VGND VPWR VPWR _17818_/X sky130_fd_sc_hd__buf_2
XFILLER_55_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19991__A2 _19985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18798_ _14261_/X _18795_/X _20762_/A _18796_/X VGND VGND VPWR VPWR _18798_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22497__A _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17749_ _17704_/X _17749_/B VGND VGND VPWR VPWR _17749_/Y sky130_fd_sc_hd__nor2_4
XFILLER_78_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16006__A1 _11982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13912__A _13909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20760_ _20518_/A VGND VGND VPWR VPWR _20760_/X sky130_fd_sc_hd__buf_2
XFILLER_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19419_ _19419_/A VGND VGND VPWR VPWR _19419_/X sky130_fd_sc_hd__buf_2
XFILLER_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20691_ _24236_/Q VGND VGND VPWR VPWR _20691_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12528__A _12528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22430_ _20670_/A VGND VGND VPWR VPWR _22430_/X sky130_fd_sc_hd__buf_2
XFILLER_56_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22361_ _22354_/A VGND VGND VPWR VPWR _22361_/X sky130_fd_sc_hd__buf_2
XANTENNA__15839__A _13009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14743__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24100_ _24321_/CLK _24100_/D HRESETn VGND VGND VPWR VPWR _24100_/Q sky130_fd_sc_hd__dfrtp_4
X_21312_ _21319_/A VGND VGND VPWR VPWR _21312_/X sky130_fd_sc_hd__buf_2
X_22292_ _22134_/X _22286_/X _14501_/B _22290_/X VGND VGND VPWR VPWR _23333_/D sky130_fd_sc_hd__o22a_4
X_24031_ _23130_/CLK _24031_/D VGND VGND VPWR VPWR _15023_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_89_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21243_ _21241_/X _21235_/X _12614_/B _21242_/X VGND VGND VPWR VPWR _23925_/D sky130_fd_sc_hd__o22a_4
XFILLER_85_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21066__B2 _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22263__B1 _16383_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12263__A _15667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21576__A _21291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21174_ _20373_/X _21169_/X _23962_/Q _21173_/X VGND VGND VPWR VPWR _21174_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13078__B _24018_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24248__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20125_ _11622_/X _20124_/X VGND VGND VPWR VPWR _20125_/X sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_5_22_0_HCLK_A clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22015__B1 _23487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19046__A _19002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20056_ _20056_/A VGND VGND VPWR VPWR _20056_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20577__B1 _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18885__A _18892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12710__B _23156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11607__A _15015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19982__A2 _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23815_ _23816_/CLK _21436_/X VGND VGND VPWR VPWR _13815_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_38_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13822__A _12211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11819_/A _11760_/B VGND VGND VPWR VPWR _11760_/X sky130_fd_sc_hd__or2_4
XFILLER_60_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_53_0_HCLK clkbuf_6_26_0_HCLK/X VGND VGND VPWR VPWR _23819_/CLK sky130_fd_sc_hd__clkbuf_1
X_20958_ _21574_/A VGND VGND VPWR VPWR _20958_/X sky130_fd_sc_hd__buf_2
X_23746_ _23363_/CLK _23746_/D VGND VGND VPWR VPWR _15260_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _16039_/A VGND VGND VPWR VPWR _11691_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _20673_/X _20880_/Y _20887_/X _20888_/Y _20692_/X VGND VGND VPWR VPWR _20889_/X
+ sky130_fd_sc_hd__a32o_4
X_23677_ _23515_/CLK _21692_/X VGND VGND VPWR VPWR _23677_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12438__A _13925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _13427_/A _13502_/B VGND VGND VPWR VPWR _13430_/X sky130_fd_sc_hd__or2_4
XFILLER_35_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22628_ _22401_/X _22622_/X _16279_/B _22626_/X VGND VGND VPWR VPWR _23129_/D sky130_fd_sc_hd__o22a_4
XFILLER_74_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19498__A1 _20650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19498__B2 HRDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16856__A1_N _16840_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _13383_/A _23728_/Q VGND VGND VPWR VPWR _13362_/C sky130_fd_sc_hd__or2_4
X_22559_ _22454_/X _22557_/X _14794_/B _22554_/X VGND VGND VPWR VPWR _23171_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14653__A _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15100_ _15108_/A _15100_/B _15100_/C VGND VGND VPWR VPWR _15100_/X sky130_fd_sc_hd__or3_4
X_12312_ _12735_/A _12312_/B VGND VGND VPWR VPWR _12312_/X sky130_fd_sc_hd__or2_4
XFILLER_33_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13292_ _13283_/X _23760_/Q VGND VGND VPWR VPWR _13293_/C sky130_fd_sc_hd__or2_4
X_16080_ _16080_/A VGND VGND VPWR VPWR _16080_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12243_ _13048_/A _12230_/X _12242_/X VGND VGND VPWR VPWR _12243_/X sky130_fd_sc_hd__or3_4
X_15031_ _14617_/A _15029_/X _15031_/C VGND VGND VPWR VPWR _15032_/C sky130_fd_sc_hd__and3_4
XANTENNA__13269__A _11656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21057__B2 _21012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24229_ _24229_/CLK _24229_/D HRESETn VGND VGND VPWR VPWR _24229_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12174_ _11774_/A _23485_/Q VGND VGND VPWR VPWR _12174_/X sky130_fd_sc_hd__or2_4
XFILLER_64_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15484__A _15484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19770_ HRDATA[16] VGND VGND VPWR VPWR _19770_/X sky130_fd_sc_hd__buf_2
X_16982_ _16946_/Y _16981_/X VGND VGND VPWR VPWR _16982_/X sky130_fd_sc_hd__or2_4
XFILLER_96_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12901__A _12518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18721_ _18720_/X VGND VGND VPWR VPWR _22824_/B sky130_fd_sc_hd__inv_2
X_15933_ _15939_/A _23256_/Q VGND VGND VPWR VPWR _15936_/B sky130_fd_sc_hd__or2_4
XFILLER_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12620__B _12620_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18652_ _18652_/A VGND VGND VPWR VPWR _19994_/A sky130_fd_sc_hd__buf_2
XFILLER_114_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19973__A2 _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15864_ _13554_/A _15864_/B VGND VGND VPWR VPWR _15865_/C sky130_fd_sc_hd__or2_4
XFILLER_92_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17603_ _17422_/A _17603_/B VGND VGND VPWR VPWR _17621_/C sky130_fd_sc_hd__nand2_4
XFILLER_76_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21780__A2 _21776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14815_ _14815_/A _14815_/B _14815_/C VGND VGND VPWR VPWR _14815_/X sky130_fd_sc_hd__and3_4
X_18583_ _17792_/A _18583_/B VGND VGND VPWR VPWR _18583_/X sky130_fd_sc_hd__and2_4
X_15795_ _12444_/A _15795_/B VGND VGND VPWR VPWR _15796_/C sky130_fd_sc_hd__or2_4
XANTENNA__22110__A _20610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14828__A _13690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17534_ _17039_/X _17533_/X _17043_/X VGND VGND VPWR VPWR _17535_/A sky130_fd_sc_hd__o21a_4
XFILLER_83_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14746_ _13925_/A _14802_/B VGND VGND VPWR VPWR _14748_/B sky130_fd_sc_hd__or2_4
X_11958_ _12739_/A VGND VGND VPWR VPWR _13428_/A sky130_fd_sc_hd__buf_2
XFILLER_36_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19736__A1_N _19674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17465_ _17586_/C VGND VGND VPWR VPWR _17476_/C sky130_fd_sc_hd__inv_2
X_14677_ _14664_/X _14677_/B _14677_/C VGND VGND VPWR VPWR _14677_/X sky130_fd_sc_hd__and3_4
X_11889_ _14101_/A VGND VGND VPWR VPWR _11890_/A sky130_fd_sc_hd__inv_2
XFILLER_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12348__A _15774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19204_ _20190_/A _24255_/Q VGND VGND VPWR VPWR _19205_/B sky130_fd_sc_hd__and2_4
XFILLER_33_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16416_ _16400_/A _23610_/Q VGND VGND VPWR VPWR _16416_/X sky130_fd_sc_hd__or2_4
X_13628_ _12509_/A VGND VGND VPWR VPWR _13645_/A sky130_fd_sc_hd__buf_2
XANTENNA__19489__A1 _19536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17396_ _17395_/B VGND VGND VPWR VPWR _17396_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19135_ _24314_/Q _19134_/X VGND VGND VPWR VPWR _19135_/X sky130_fd_sc_hd__and2_4
X_16347_ _16185_/A _16279_/B VGND VGND VPWR VPWR _16347_/X sky130_fd_sc_hd__or2_4
XANTENNA__15659__A _12284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13559_ _13559_/A _13485_/B VGND VGND VPWR VPWR _13560_/C sky130_fd_sc_hd__or2_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24076__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14563__A _11656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19066_ _11512_/B VGND VGND VPWR VPWR _19066_/Y sky130_fd_sc_hd__inv_2
X_16278_ _15980_/A _16274_/X _16277_/X VGND VGND VPWR VPWR _16278_/X sky130_fd_sc_hd__or3_4
XFILLER_51_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18017_ _16986_/X VGND VGND VPWR VPWR _18017_/Y sky130_fd_sc_hd__inv_2
X_15229_ _15234_/A _15166_/B VGND VGND VPWR VPWR _15229_/X sky130_fd_sc_hd__or2_4
XANTENNA__17874__A _17874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13179__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21599__A2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13907__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19968_ _18653_/X _17769_/A _19934_/X _19967_/X VGND VGND VPWR VPWR _19968_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22548__B2 _22547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18919_ _15121_/X _18891_/A _20968_/A _18892_/A VGND VGND VPWR VPWR _24352_/D sky130_fd_sc_hd__o22a_4
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19413__B2 _17736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19899_ _19909_/A VGND VGND VPWR VPWR _19899_/X sky130_fd_sc_hd__buf_2
XFILLER_110_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21930_ _21802_/X _21924_/X _16260_/B _21928_/X VGND VGND VPWR VPWR _21930_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21220__B2 _21218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21771__A2 _21769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21861_ _21291_/A VGND VGND VPWR VPWR _21861_/X sky130_fd_sc_hd__buf_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22020__A _22035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20812_ _18570_/X _20653_/X _20758_/X _20811_/Y VGND VGND VPWR VPWR _20813_/A sky130_fd_sc_hd__a211o_4
X_23600_ _23635_/CLK _21825_/X VGND VGND VPWR VPWR _23600_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13642__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21792_ _21792_/A VGND VGND VPWR VPWR _21817_/A sky130_fd_sc_hd__buf_2
XANTENNA__13461__A1 _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21523__A2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22955__A _22985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20743_ _20743_/A VGND VGND VPWR VPWR _20743_/Y sky130_fd_sc_hd__inv_2
X_23531_ _24044_/CLK _23531_/D VGND VGND VPWR VPWR _23531_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12258__A _12742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23462_ _23781_/CLK _22057_/X VGND VGND VPWR VPWR _14317_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22470__A2_N _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20674_ _20642_/X VGND VGND VPWR VPWR _22821_/A sky130_fd_sc_hd__buf_2
XFILLER_56_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22413_ _22413_/A VGND VGND VPWR VPWR _22413_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15569__A _12441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22484__B1 _12667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23393_ _24032_/CLK _23393_/D VGND VGND VPWR VPWR _15166_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14473__A _13020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22344_ _22344_/A VGND VGND VPWR VPWR _22344_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22690__A _22683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21039__B2 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22275_ _22105_/X _22272_/X _13140_/B _22269_/X VGND VGND VPWR VPWR _23345_/D sky130_fd_sc_hd__o22a_4
XFILLER_30_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24014_ _24044_/CLK _21090_/X VGND VGND VPWR VPWR _15724_/B sky130_fd_sc_hd__dfxtp_4
X_21226_ _21225_/X _21223_/X _23932_/Q _21218_/X VGND VGND VPWR VPWR _21226_/X sky130_fd_sc_hd__o22a_4
XFILLER_3_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21157_ _20937_/X _21154_/X _15267_/B _21151_/X VGND VGND VPWR VPWR _23970_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13817__A _13794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12721__A _15689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22539__B2 _22533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20108_ _19931_/B _20107_/X _24451_/Q _19957_/X VGND VGND VPWR VPWR _20108_/X sky130_fd_sc_hd__o22a_4
XFILLER_115_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21088_ _20611_/X _21082_/X _13513_/B _21086_/X VGND VGND VPWR VPWR _24015_/D sky130_fd_sc_hd__o22a_4
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14492__A3 _14461_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12930_ _12982_/A _12930_/B _12929_/X VGND VGND VPWR VPWR _12930_/X sky130_fd_sc_hd__and3_4
X_20039_ _18433_/X _20033_/X _20038_/Y _20020_/X VGND VGND VPWR VPWR _20039_/X sky130_fd_sc_hd__o22a_4
XFILLER_86_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23026__A _22967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ _12861_/A VGND VGND VPWR VPWR _12862_/A sky130_fd_sc_hd__buf_2
XANTENNA__15751__B _15686_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14600_ _14617_/A _14598_/X _14600_/C VGND VGND VPWR VPWR _14604_/B sky130_fd_sc_hd__and3_4
XFILLER_27_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13552__A _13551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11812_ _11692_/X _11810_/X _11811_/X VGND VGND VPWR VPWR _11812_/X sky130_fd_sc_hd__and3_4
XFILLER_15_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15580_ _13682_/A _15579_/X VGND VGND VPWR VPWR _15580_/X sky130_fd_sc_hd__and2_4
XFILLER_76_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12792_ _12792_/A VGND VGND VPWR VPWR _12802_/A sky130_fd_sc_hd__buf_2
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22711__A1 _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22711__B2 _22668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14531_ _11664_/A _14514_/X _14531_/C VGND VGND VPWR VPWR _14531_/X sky130_fd_sc_hd__or3_4
XFILLER_18_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _13370_/A VGND VGND VPWR VPWR _13422_/A sky130_fd_sc_hd__buf_2
X_23729_ _23122_/CLK _23729_/D VGND VGND VPWR VPWR _13141_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17959__A _17779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17911_/A _17247_/Y _17249_/X VGND VGND VPWR VPWR _17250_/X sky130_fd_sc_hd__o21a_4
XFILLER_57_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _12441_/A _14532_/B VGND VGND VPWR VPWR _14462_/X sky130_fd_sc_hd__or2_4
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11673_/X VGND VGND VPWR VPWR _16180_/A sky130_fd_sc_hd__buf_2
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ _16201_/A _16124_/B VGND VGND VPWR VPWR _16201_/X sky130_fd_sc_hd__or2_4
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _13378_/X _13344_/B VGND VGND VPWR VPWR _13414_/C sky130_fd_sc_hd__or2_4
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17181_ _12841_/X VGND VGND VPWR VPWR _17181_/X sky130_fd_sc_hd__buf_2
XANTENNA__15479__A _12646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14393_ _15598_/A _14304_/B VGND VGND VPWR VPWR _14393_/X sky130_fd_sc_hd__or2_4
X_16132_ _16108_/A _16132_/B VGND VGND VPWR VPWR _16133_/C sky130_fd_sc_hd__or2_4
XANTENNA__11800__A _12392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13344_ _15785_/A _13344_/B VGND VGND VPWR VPWR _13344_/X sky130_fd_sc_hd__or2_4
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16063_ _16063_/A _16063_/B _16062_/X VGND VGND VPWR VPWR _16067_/B sky130_fd_sc_hd__and3_4
X_13275_ _13059_/Y _13274_/X VGND VGND VPWR VPWR _13277_/A sky130_fd_sc_hd__and2_4
XANTENNA__12715__B1 _12706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15014_ _15041_/A _23423_/Q VGND VGND VPWR VPWR _15015_/C sky130_fd_sc_hd__or2_4
X_12226_ _12556_/A _12214_/X _12225_/X VGND VGND VPWR VPWR _12226_/X sky130_fd_sc_hd__or3_4
XFILLER_100_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22105__A _20573_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12157_ _12169_/A _12155_/X _12157_/C VGND VGND VPWR VPWR _12157_/X sky130_fd_sc_hd__and3_4
X_19822_ _19822_/A _19829_/B VGND VGND VPWR VPWR _19822_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__13727__A _13735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12631__A _13737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12088_ _12088_/A _12088_/B _12088_/C VGND VGND VPWR VPWR _12089_/C sky130_fd_sc_hd__and3_4
X_16965_ _17734_/A _17735_/A _16965_/C VGND VGND VPWR VPWR _18642_/A sky130_fd_sc_hd__or3_4
X_19753_ _20939_/B _19496_/X _19752_/X _19616_/X VGND VGND VPWR VPWR _19753_/X sky130_fd_sc_hd__a211o_4
XFILLER_110_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15916_ _13776_/A _13922_/Y _13774_/X VGND VGND VPWR VPWR _16841_/A sky130_fd_sc_hd__o21ai_4
X_18704_ _17740_/X VGND VGND VPWR VPWR _18704_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15942__A _16095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21202__B2 _21201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19684_ _19637_/Y _19643_/B VGND VGND VPWR VPWR _19759_/B sky130_fd_sc_hd__and2_4
X_16896_ _12033_/X _12187_/X VGND VGND VPWR VPWR _16903_/B sky130_fd_sc_hd__nor2_4
XFILLER_49_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21753__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18635_ _18500_/X _18634_/Y _17305_/A VGND VGND VPWR VPWR _18635_/X sky130_fd_sc_hd__o21a_4
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15847_ _13550_/A _15847_/B _15847_/C VGND VGND VPWR VPWR _15851_/B sky130_fd_sc_hd__and3_4
XFILLER_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14558__A _13697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18566_ _18714_/A _17387_/X _17782_/Y VGND VGND VPWR VPWR _18566_/X sky130_fd_sc_hd__a21o_4
X_15778_ _12989_/A _15746_/X _15777_/X VGND VGND VPWR VPWR _15778_/X sky130_fd_sc_hd__and3_4
XFILLER_79_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14640__B1 _11594_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17517_ _17195_/Y _17517_/B VGND VGND VPWR VPWR _17517_/X sky130_fd_sc_hd__or2_4
XANTENNA__22702__B2 _22697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14729_ _14756_/A _14791_/B VGND VGND VPWR VPWR _14730_/C sky130_fd_sc_hd__or2_4
X_18497_ _17961_/X _18248_/Y _17856_/X _18496_/Y VGND VGND VPWR VPWR _18497_/X sky130_fd_sc_hd__a211o_4
XANTENNA__12078__A _11997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17448_ _17447_/X VGND VGND VPWR VPWR _18254_/A sky130_fd_sc_hd__inv_2
XANTENNA__20295__A _20556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23466__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16492__B _16423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21269__B2 _21266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17379_ _15909_/B _17377_/B VGND VGND VPWR VPWR _17380_/B sky130_fd_sc_hd__and2_4
XANTENNA__12806__A _12822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19118_ _24297_/Q _19118_/B VGND VGND VPWR VPWR _19181_/A sky130_fd_sc_hd__and2_4
XANTENNA__11710__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20390_ _24249_/Q _20283_/X _20389_/X VGND VGND VPWR VPWR _20391_/B sky130_fd_sc_hd__o21a_4
XFILLER_118_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19882__A1 _19554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19049_ _24362_/Q VGND VGND VPWR VPWR _19049_/Y sky130_fd_sc_hd__inv_2
X_22060_ _21852_/X _22059_/X _14624_/B _22056_/X VGND VGND VPWR VPWR _23460_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15836__B _15836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21011_ _21015_/A VGND VGND VPWR VPWR _21027_/A sky130_fd_sc_hd__inv_2
XFILLER_47_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13637__A _15411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21441__A1 _21282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21441__B2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12541__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18866__C _12068_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22962_ _22962_/A _22962_/B VGND VGND VPWR VPWR _22962_/Y sky130_fd_sc_hd__nand2_4
XFILLER_110_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21744__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21913_ _21861_/X _21908_/X _23552_/Q _21869_/X VGND VGND VPWR VPWR _21913_/X sky130_fd_sc_hd__o22a_4
XFILLER_3_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22893_ _18700_/X _22889_/X _22892_/X VGND VGND VPWR VPWR _22893_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14468__A _12460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20952__B1 _20640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21844_ _21843_/X _21841_/X _23592_/Q _21836_/X VGND VGND VPWR VPWR _23592_/D sky130_fd_sc_hd__o22a_4
XFILLER_110_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21775_ _21565_/X _21769_/X _14480_/B _21773_/X VGND VGND VPWR VPWR _23621_/D sky130_fd_sc_hd__o22a_4
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17779__A _18063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20726_ _20699_/B VGND VGND VPWR VPWR _20821_/B sky130_fd_sc_hd__buf_2
X_23514_ _23514_/CLK _23514_/D VGND VGND VPWR VPWR _16381_/B sky130_fd_sc_hd__dfxtp_4
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20657_ _20657_/A _20521_/B VGND VGND VPWR VPWR _20657_/X sky130_fd_sc_hd__or2_4
X_23445_ _23699_/CLK _23445_/D VGND VGND VPWR VPWR _12623_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19994__A _19994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12716__A _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18125__B2 _18124_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11620__A _11619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23376_ _23472_/CLK _22227_/X VGND VGND VPWR VPWR _13328_/B sky130_fd_sc_hd__dfxtp_4
X_20588_ _20588_/A _20588_/B VGND VGND VPWR VPWR _20588_/Y sky130_fd_sc_hd__nand2_4
XFILLER_87_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20483__A2 _20421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22209__B1 _12162_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22327_ _14742_/B VGND VGND VPWR VPWR _23299_/D sky130_fd_sc_hd__buf_2
XANTENNA__21680__B2 _21637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14931__A _14002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13060_ _12626_/A VGND VGND VPWR VPWR _13101_/A sky130_fd_sc_hd__buf_2
X_22258_ _22272_/A VGND VGND VPWR VPWR _22258_/X sky130_fd_sc_hd__buf_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12011_ _12011_/A _12011_/B _12011_/C VGND VGND VPWR VPWR _12017_/B sky130_fd_sc_hd__and3_4
XFILLER_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21209_ _20982_/X _21204_/X _14889_/B _21165_/X VGND VGND VPWR VPWR _23936_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13547__A _13546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21432__B2 _21430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22189_ _22129_/X _22186_/X _23399_/Q _22183_/X VGND VGND VPWR VPWR _22189_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12451__A _12494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20090__D _20090_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12170__B _23709_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16750_ _11758_/X VGND VGND VPWR VPWR _16773_/A sky130_fd_sc_hd__buf_2
XFILLER_59_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13962_ _13966_/A _23594_/Q VGND VGND VPWR VPWR _13964_/B sky130_fd_sc_hd__or2_4
XFILLER_86_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15701_ _12849_/A _15699_/X _15701_/C VGND VGND VPWR VPWR _15701_/X sky130_fd_sc_hd__and3_4
X_12913_ _12493_/A _12911_/X _12913_/C VGND VGND VPWR VPWR _12913_/X sky130_fd_sc_hd__and3_4
X_16681_ _16681_/A VGND VGND VPWR VPWR _16681_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18600__A2 _18576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13893_ _13893_/A _13889_/X _13893_/C VGND VGND VPWR VPWR _13893_/X sky130_fd_sc_hd__or3_4
XFILLER_74_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24367__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18420_ _18101_/A _17380_/B VGND VGND VPWR VPWR _18420_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13282__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15632_ _15632_/A _23691_/Q VGND VGND VPWR VPWR _15634_/B sky130_fd_sc_hd__or2_4
X_12844_ _12843_/X VGND VGND VPWR VPWR _12845_/B sky130_fd_sc_hd__inv_2
XFILLER_62_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18351_ _18344_/X _18351_/B VGND VGND VPWR VPWR _18352_/B sky130_fd_sc_hd__or2_4
X_15563_ _15556_/A _23403_/Q VGND VGND VPWR VPWR _15563_/X sky130_fd_sc_hd__or2_4
XFILLER_61_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17689__A _16945_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22696__B1 _23084_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12775_ _13563_/A _12775_/B _12775_/C VGND VGND VPWR VPWR _12775_/X sky130_fd_sc_hd__and3_4
XFILLER_37_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_23_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_46_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16593__A _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17302_/A VGND VGND VPWR VPWR _17309_/B sky130_fd_sc_hd__inv_2
X_14514_ _11670_/A _14504_/X _14513_/X VGND VGND VPWR VPWR _14514_/X sky130_fd_sc_hd__and3_4
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _15743_/A VGND VGND VPWR VPWR _12830_/A sky130_fd_sc_hd__buf_2
X_18282_ _18281_/A _18280_/X _18160_/X VGND VGND VPWR VPWR _18282_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15494_/A _23820_/Q VGND VGND VPWR VPWR _15494_/X sky130_fd_sc_hd__or2_4
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17233_ _17130_/X _17231_/X _17815_/A _17232_/X VGND VGND VPWR VPWR _17233_/X sky130_fd_sc_hd__o22a_4
X_14445_ _12460_/A _14441_/X _14445_/C VGND VGND VPWR VPWR _14445_/X sky130_fd_sc_hd__or3_4
XANTENNA__22448__B1 _14268_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _12989_/A VGND VGND VPWR VPWR _11657_/X sky130_fd_sc_hd__buf_2
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15002__A _14119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17164_ _16077_/X VGND VGND VPWR VPWR _17164_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _15631_/A _14373_/X _14376_/C VGND VGND VPWR VPWR _14377_/C sky130_fd_sc_hd__and3_4
XANTENNA__18667__A2 _18654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11588_ _17343_/A VGND VGND VPWR VPWR _17040_/A sky130_fd_sc_hd__buf_2
XANTENNA__19864__B2 _19775_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16115_ _16146_/A _23575_/Q VGND VGND VPWR VPWR _16116_/C sky130_fd_sc_hd__or2_4
X_13327_ _13281_/X _13325_/X _13326_/X VGND VGND VPWR VPWR _13327_/X sky130_fd_sc_hd__and3_4
XANTENNA__17875__B1 _17871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17095_ _17047_/Y _18421_/A VGND VGND VPWR VPWR _17095_/X sky130_fd_sc_hd__and2_4
XANTENNA__21671__B2 _21666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14841__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16046_ _16019_/A _23896_/Q VGND VGND VPWR VPWR _16046_/X sky130_fd_sc_hd__or2_4
X_13258_ _12350_/A _13256_/X _13258_/C VGND VGND VPWR VPWR _13258_/X sky130_fd_sc_hd__and3_4
XANTENNA__24114__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12209_ _12209_/A VGND VGND VPWR VPWR _13635_/A sky130_fd_sc_hd__buf_2
XANTENNA__13457__A _12477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13189_ _15707_/A VGND VGND VPWR VPWR _15785_/A sky130_fd_sc_hd__buf_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20631__C1 _20630_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19805_ _19877_/A _19804_/X VGND VGND VPWR VPWR _19805_/Y sky130_fd_sc_hd__nor2_4
XFILLER_97_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17997_ _18048_/A VGND VGND VPWR VPWR _18160_/A sky130_fd_sc_hd__buf_2
XFILLER_97_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15672__A _15695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16948_ _24128_/Q VGND VGND VPWR VPWR _16948_/Y sky130_fd_sc_hd__inv_2
X_19736_ _19674_/X _19734_/Y _20895_/B _19551_/A VGND VGND VPWR VPWR _19736_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_105_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR _23155_/CLK sky130_fd_sc_hd__clkbuf_1
X_16879_ _16851_/X _16876_/X _16879_/C _16879_/D VGND VGND VPWR VPWR _16879_/X sky130_fd_sc_hd__and4_4
X_19667_ _19667_/A _19667_/B VGND VGND VPWR VPWR _19667_/X sky130_fd_sc_hd__and2_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13192__A _15820_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11705__A _11803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18618_ _18216_/A _18075_/Y VGND VGND VPWR VPWR _18618_/X sky130_fd_sc_hd__and2_4
XFILLER_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19598_ _19598_/A VGND VGND VPWR VPWR _19800_/B sky130_fd_sc_hd__buf_2
XFILLER_53_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18549_ _18458_/X _18536_/Y _18485_/X _18548_/X VGND VGND VPWR VPWR _18549_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21560_ _20819_/A VGND VGND VPWR VPWR _21560_/X sky130_fd_sc_hd__buf_2
XFILLER_33_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20511_ _20511_/A VGND VGND VPWR VPWR _20511_/X sky130_fd_sc_hd__buf_2
X_21491_ _21455_/A VGND VGND VPWR VPWR _21491_/X sky130_fd_sc_hd__buf_2
XANTENNA__12536__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16008__A _16007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23230_ _23358_/CLK _22470_/X VGND VGND VPWR VPWR _12014_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20442_ _20442_/A VGND VGND VPWR VPWR _20442_/X sky130_fd_sc_hd__buf_2
XFILLER_88_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19855__A1 _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20753__A HRDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23161_ _23354_/CLK _23161_/D VGND VGND VPWR VPWR _16266_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20373_ _21799_/A VGND VGND VPWR VPWR _20373_/X sky130_fd_sc_hd__buf_2
XANTENNA__15847__A _13550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14751__A _14778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22112_ _22112_/A VGND VGND VPWR VPWR _22112_/X sky130_fd_sc_hd__buf_2
X_23092_ _23315_/CLK _23092_/D VGND VGND VPWR VPWR _12823_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15566__B _23467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22043_ _21823_/X _22038_/X _23472_/Q _22042_/X VGND VGND VPWR VPWR _22043_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21414__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12271__A _12240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21965__A2 _21938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16678__A _16077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23994_ _23699_/CLK _21124_/X VGND VGND VPWR VPWR _16398_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21717__A2 _21712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22945_ _18506_/X _22945_/B VGND VGND VPWR VPWR _22946_/C sky130_fd_sc_hd__or2_4
XFILLER_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19791__B1 _19429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22876_ _19893_/X _22818_/X _15910_/Y _22855_/A VGND VGND VPWR VPWR _22876_/X sky130_fd_sc_hd__o22a_4
X_21827_ _21826_/X _21817_/X _23599_/Q _21824_/X VGND VGND VPWR VPWR _21827_/X sky130_fd_sc_hd__o22a_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14926__A _13992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22142__A2 _22137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _11670_/A VGND VGND VPWR VPWR _13770_/A sky130_fd_sc_hd__buf_2
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21758_ _21536_/X _21755_/X _13190_/B _21752_/X VGND VGND VPWR VPWR _23633_/D sky130_fd_sc_hd__o22a_4
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11511_ _11511_/A _11511_/B VGND VGND VPWR VPWR _11512_/B sky130_fd_sc_hd__or2_4
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20709_ _20473_/A VGND VGND VPWR VPWR _20709_/X sky130_fd_sc_hd__buf_2
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _13009_/A VGND VGND VPWR VPWR _12905_/A sky130_fd_sc_hd__buf_2
X_24477_ _24229_/CLK _24477_/D HRESETn VGND VGND VPWR VPWR _24477_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21689_ _21683_/Y _21688_/X _21504_/X _21688_/X VGND VGND VPWR VPWR _23678_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _14218_/A VGND VGND VPWR VPWR _14252_/A sky130_fd_sc_hd__buf_2
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23428_ _23812_/CLK _22138_/X VGND VGND VPWR VPWR _14676_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21759__A _21752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14161_ _14161_/A _23625_/Q VGND VGND VPWR VPWR _14161_/X sky130_fd_sc_hd__or2_4
XFILLER_50_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23359_ _23487_/CLK _22249_/X VGND VGND VPWR VPWR _15097_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21653__B2 _21652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14661__A _15105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13112_ _13112_/A _13112_/B VGND VGND VPWR VPWR _13113_/C sky130_fd_sc_hd__or2_4
X_14092_ _14991_/A VGND VGND VPWR VPWR _14098_/A sky130_fd_sc_hd__buf_2
XFILLER_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13043_ _13016_/A _24082_/Q VGND VGND VPWR VPWR _13043_/X sky130_fd_sc_hd__or2_4
X_17920_ _17811_/A VGND VGND VPWR VPWR _17921_/A sky130_fd_sc_hd__buf_2
XFILLER_78_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12181__A _11675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17851_ _17837_/X _17844_/X _17846_/X _17850_/X VGND VGND VPWR VPWR _17851_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18282__B1 _18160_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16588__A _12020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16802_ _16598_/X _16798_/X _16802_/C VGND VGND VPWR VPWR _16802_/X sky130_fd_sc_hd__or3_4
X_17782_ _18101_/A VGND VGND VPWR VPWR _17782_/Y sky130_fd_sc_hd__inv_2
X_14994_ _14994_/A _14994_/B _14994_/C VGND VGND VPWR VPWR _14995_/C sky130_fd_sc_hd__and3_4
XFILLER_19_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22905__A1 _22886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21708__A2 _21705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16733_ _12051_/X _16729_/X _16732_/X VGND VGND VPWR VPWR _16733_/X sky130_fd_sc_hd__or3_4
X_19521_ _19458_/X _19520_/X HRDATA[6] _19462_/X VGND VGND VPWR VPWR _19521_/X sky130_fd_sc_hd__o22a_4
X_13945_ _13643_/A _22320_/A VGND VGND VPWR VPWR _13947_/B sky130_fd_sc_hd__or2_4
XANTENNA__19899__A _19909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22381__A2 _22354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19452_ _19416_/B VGND VGND VPWR VPWR _19712_/A sky130_fd_sc_hd__buf_2
X_16664_ _16652_/A _16662_/X _16664_/C VGND VGND VPWR VPWR _16668_/B sky130_fd_sc_hd__and3_4
X_13876_ _12617_/A _13873_/X _13876_/C VGND VGND VPWR VPWR _13877_/C sky130_fd_sc_hd__and3_4
XFILLER_90_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15615_ _15615_/A _23947_/Q VGND VGND VPWR VPWR _15615_/X sky130_fd_sc_hd__or2_4
X_18403_ _18428_/A _18402_/X _17434_/Y VGND VGND VPWR VPWR _18403_/Y sky130_fd_sc_hd__o21ai_4
X_12827_ _12827_/A _12827_/B VGND VGND VPWR VPWR _12830_/B sky130_fd_sc_hd__or2_4
X_19383_ _19377_/X _19382_/Y _19380_/X _24212_/Q VGND VGND VPWR VPWR _19383_/X sky130_fd_sc_hd__o22a_4
X_16595_ _11844_/X _11620_/X _16563_/X _11598_/X _16594_/X VGND VGND VPWR VPWR _16596_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14836__A _14050_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22133__A2 _22125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20557__B _20595_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18334_ _18317_/X _18322_/Y _18328_/X _18332_/X _18333_/Y VGND VGND VPWR VPWR _18334_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_91_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13740__A _11664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15546_ _15576_/A _23147_/Q VGND VGND VPWR VPWR _15546_/X sky130_fd_sc_hd__or2_4
XANTENNA__19351__A2_N _18648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12758_ _12808_/A _12758_/B VGND VGND VPWR VPWR _12758_/X sky130_fd_sc_hd__or2_4
XFILLER_37_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17569__D _17568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _11709_/A VGND VGND VPWR VPWR _11710_/A sky130_fd_sc_hd__buf_2
X_18265_ _18265_/A _17501_/X VGND VGND VPWR VPWR _18265_/Y sky130_fd_sc_hd__nor2_4
XFILLER_72_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21892__A1 _21823_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20695__A2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15477_ _15477_/A _15406_/B VGND VGND VPWR VPWR _15477_/X sky130_fd_sc_hd__or2_4
XANTENNA__21892__B2 _21891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12689_ _12556_/A _12689_/B _12689_/C VGND VGND VPWR VPWR _12689_/X sky130_fd_sc_hd__or3_4
XFILLER_15_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12356__A _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17216_ _17227_/A _17208_/Y _17251_/A _17215_/Y VGND VGND VPWR VPWR _17216_/X sky130_fd_sc_hd__o22a_4
X_14428_ _14428_/A VGND VGND VPWR VPWR _14429_/B sky130_fd_sc_hd__buf_2
XANTENNA__21669__A _21636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18196_ _18009_/X _18194_/X _18053_/X _18195_/X VGND VGND VPWR VPWR _18196_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20573__A _20573_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19366__A2_N _17004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17147_ _17141_/X _17142_/X _17163_/A _17146_/X VGND VGND VPWR VPWR _17147_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15667__A _15667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14359_ _14359_/A VGND VGND VPWR VPWR _15598_/A sky130_fd_sc_hd__buf_2
XFILLER_89_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21644__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18043__A _17259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23504__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17078_ _17046_/B VGND VGND VPWR VPWR _17081_/A sky130_fd_sc_hd__inv_2
XFILLER_118_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16029_ _16180_/A _16029_/B _16029_/C VGND VGND VPWR VPWR _16045_/B sky130_fd_sc_hd__and3_4
XANTENNA__13187__A _12737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21947__A2 _21945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13915__A _11740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19719_ _19719_/A _19880_/B VGND VGND VPWR VPWR _19720_/B sky130_fd_sc_hd__or2_4
X_20991_ _20255_/A _20990_/X _24351_/Q _18870_/X VGND VGND VPWR VPWR _20991_/X sky130_fd_sc_hd__o22a_4
XFILLER_26_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19773__B1 _19592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22730_ _24099_/Q VGND VGND VPWR VPWR _22730_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19602__A _19598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24350__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22661_ _22458_/X _22657_/X _15225_/B _22626_/A VGND VGND VPWR VPWR _23105_/D sky130_fd_sc_hd__o22a_4
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14746__A _13925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24400_ _23326_/CLK _24400_/D HRESETn VGND VGND VPWR VPWR _24400_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13650__A _13647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21612_ _21605_/A VGND VGND VPWR VPWR _21612_/X sky130_fd_sc_hd__buf_2
XFILLER_90_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22592_ _22425_/X _22586_/X _13456_/B _22590_/X VGND VGND VPWR VPWR _23151_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22963__A _18430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24331_ _23260_/CLK _24331_/D HRESETn VGND VGND VPWR VPWR _24331_/Q sky130_fd_sc_hd__dfstp_4
X_21543_ _21543_/A VGND VGND VPWR VPWR _21543_/X sky130_fd_sc_hd__buf_2
XANTENNA__21883__B2 _21877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21474_ _21467_/A VGND VGND VPWR VPWR _21474_/X sky130_fd_sc_hd__buf_2
X_24262_ _24305_/CLK _19284_/X HRESETn VGND VGND VPWR VPWR _19211_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19828__A1 _19429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20425_ _20425_/A VGND VGND VPWR VPWR _20425_/X sky130_fd_sc_hd__buf_2
X_23213_ _23564_/CLK _23213_/D VGND VGND VPWR VPWR _15831_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15577__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20438__A2 _20421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24193_ _24199_/CLK _24193_/D HRESETn VGND VGND VPWR VPWR _24193_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14481__A _12465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20356_ _21797_/A VGND VGND VPWR VPWR _20356_/X sky130_fd_sc_hd__buf_2
X_23144_ _23304_/CLK _23144_/D VGND VGND VPWR VPWR _13727_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_1_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13097__A _13097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23075_ _23907_/CLK _23075_/D VGND VGND VPWR VPWR _14776_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17792__A _17792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20287_ _20285_/X _20650_/A _20286_/X VGND VGND VPWR VPWR _20287_/X sky130_fd_sc_hd__a21o_4
XFILLER_27_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12679__A2 _12676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22026_ _21795_/X _22024_/X _23484_/Q _22021_/X VGND VGND VPWR VPWR _22026_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22060__A1 _21852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22060__B2 _22056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22203__A _22207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13825__A _13636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11991_ _16741_/A _11924_/X _11947_/X _11973_/X _11990_/X VGND VGND VPWR VPWR _11991_/X
+ sky130_fd_sc_hd__a32o_4
X_23977_ _23910_/CLK _23977_/D VGND VGND VPWR VPWR _23977_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22363__A2 _22361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13730_ _15491_/A _13730_/B _13729_/X VGND VGND VPWR VPWR _13730_/X sky130_fd_sc_hd__and3_4
XFILLER_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19512__A _19754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22928_ _18570_/X _22945_/B VGND VGND VPWR VPWR _22929_/C sky130_fd_sc_hd__or2_4
XFILLER_43_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13661_ _13641_/A VGND VGND VPWR VPWR _15430_/A sky130_fd_sc_hd__buf_2
X_22859_ _22854_/X _22801_/X _13685_/Y _22855_/X VGND VGND VPWR VPWR _22859_/X sky130_fd_sc_hd__o22a_4
XFILLER_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14656__A _15108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15400_ _13620_/A _15463_/B VGND VGND VPWR VPWR _15401_/C sky130_fd_sc_hd__or2_4
XFILLER_71_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13560__A _13511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12612_ _12612_/A VGND VGND VPWR VPWR _13118_/A sky130_fd_sc_hd__buf_2
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ _15959_/A _16380_/B VGND VGND VPWR VPWR _16380_/X sky130_fd_sc_hd__or2_4
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13592_ _13493_/X _13591_/X _13578_/Y VGND VGND VPWR VPWR _13593_/B sky130_fd_sc_hd__a21o_4
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15331_ _13991_/A _15331_/B _15330_/X VGND VGND VPWR VPWR _15347_/B sky130_fd_sc_hd__and3_4
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12543_ _12500_/X _24085_/Q VGND VGND VPWR VPWR _12544_/C sky130_fd_sc_hd__or2_4
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18050_ _18024_/X _18032_/Y _18044_/X _18047_/X _18049_/Y VGND VGND VPWR VPWR _18050_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15262_ _14113_/A _15262_/B VGND VGND VPWR VPWR _15262_/X sky130_fd_sc_hd__or2_4
X_12474_ _13799_/A VGND VGND VPWR VPWR _12475_/A sky130_fd_sc_hd__buf_2
XANTENNA__20393__A _20393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17001_ _17889_/A _18013_/B _17001_/C VGND VGND VPWR VPWR _17001_/X sky130_fd_sc_hd__and3_4
X_14213_ _14204_/A _23657_/Q VGND VGND VPWR VPWR _14215_/B sky130_fd_sc_hd__or2_4
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15487__A _15487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15193_ _14644_/A _15132_/B VGND VGND VPWR VPWR _15193_/X sky130_fd_sc_hd__or2_4
XANTENNA__12904__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14144_ _14117_/A _14144_/B _14144_/C VGND VGND VPWR VPWR _14144_/X sky130_fd_sc_hd__and3_4
XFILLER_113_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14075_ _14074_/A _14073_/X VGND VGND VPWR VPWR _14075_/X sky130_fd_sc_hd__or2_4
X_18952_ _18937_/X _18951_/X _18937_/X _11532_/A VGND VGND VPWR VPWR _24347_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21929__A2 _21924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13026_ _13026_/A _13026_/B VGND VGND VPWR VPWR _13026_/X sky130_fd_sc_hd__and2_4
X_17903_ _18443_/A _17278_/X VGND VGND VPWR VPWR _17904_/D sky130_fd_sc_hd__and2_4
XANTENNA__18255__B1 _18048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22051__B2 _22049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18883_ _16514_/X _18875_/X _18954_/A _18878_/X VGND VGND VPWR VPWR _24378_/D sky130_fd_sc_hd__o22a_4
XFILLER_79_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22113__A _22101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13735__A _13735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17834_ _17798_/X _17821_/X _17823_/X _17833_/X VGND VGND VPWR VPWR _17834_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16111__A _16139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21952__A _21919_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14977_ _14970_/A _23456_/Q VGND VGND VPWR VPWR _14979_/B sky130_fd_sc_hd__or2_4
X_17765_ _17765_/A _17648_/Y _17765_/C _17764_/Y VGND VGND VPWR VPWR _17765_/X sky130_fd_sc_hd__or4_4
X_19504_ _19599_/B _19719_/A VGND VGND VPWR VPWR _19535_/A sky130_fd_sc_hd__or2_4
XANTENNA__15950__A _15959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13928_ _14778_/A _13925_/X _13928_/C VGND VGND VPWR VPWR _13928_/X sky130_fd_sc_hd__and3_4
X_16716_ _16713_/A _23611_/Q VGND VGND VPWR VPWR _16718_/B sky130_fd_sc_hd__or2_4
X_17696_ _17696_/A _17696_/B VGND VGND VPWR VPWR _17754_/B sky130_fd_sc_hd__or2_4
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16647_ _16617_/A _23900_/Q VGND VGND VPWR VPWR _16649_/B sky130_fd_sc_hd__or2_4
X_19435_ _19435_/A VGND VGND VPWR VPWR _19435_/X sky130_fd_sc_hd__buf_2
X_13859_ _13878_/A _13859_/B VGND VGND VPWR VPWR _13859_/X sky130_fd_sc_hd__or2_4
XANTENNA__14566__A _14492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22106__A2 _22101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16578_ _16586_/A VGND VGND VPWR VPWR _16686_/A sky130_fd_sc_hd__buf_2
X_19366_ _19359_/X _17004_/X _19359_/X _24221_/Q VGND VGND VPWR VPWR _19366_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22783__A _15051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15529_ _12257_/A _23179_/Q VGND VGND VPWR VPWR _15529_/X sky130_fd_sc_hd__or2_4
X_18317_ _18204_/A _17495_/A VGND VGND VPWR VPWR _18317_/X sky130_fd_sc_hd__or2_4
XFILLER_31_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19297_ _20190_/A VGND VGND VPWR VPWR _22924_/A sky130_fd_sc_hd__buf_2
XFILLER_31_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18248_ _18248_/A VGND VGND VPWR VPWR _18248_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24452__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15397__A _15424_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18179_ _18297_/A _17472_/Y VGND VGND VPWR VPWR _18180_/D sky130_fd_sc_hd__and2_4
XFILLER_89_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21617__B2 _21616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20210_ _20210_/A _20209_/X VGND VGND VPWR VPWR _20210_/X sky130_fd_sc_hd__or2_4
XFILLER_85_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21190_ _21183_/A VGND VGND VPWR VPWR _21190_/X sky130_fd_sc_hd__buf_2
X_20141_ _24426_/Q VGND VGND VPWR VPWR _20141_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20072_ _20071_/X VGND VGND VPWR VPWR _20077_/B sky130_fd_sc_hd__inv_2
XFILLER_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22023__A _22052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18797__A1 _17171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23900_ _23931_/CLK _21307_/X VGND VGND VPWR VPWR _23900_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13645__A _13645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22958__A _18453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23831_ _23632_/CLK _21414_/X VGND VGND VPWR VPWR _16132_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13364__B _13291_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15860__A _13546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19746__B1 _19672_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18549__B2 _18548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19332__A _19328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23762_ _23314_/CLK _21535_/X VGND VGND VPWR VPWR _13075_/B sky130_fd_sc_hd__dfxtp_4
X_20974_ _20424_/A _20974_/B VGND VGND VPWR VPWR _20974_/Y sky130_fd_sc_hd__nor2_4
X_22713_ _21293_/A _22686_/A _23071_/Q _22668_/X VGND VGND VPWR VPWR _23071_/D sky130_fd_sc_hd__o22a_4
XFILLER_92_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23693_ _23826_/CLK _21664_/X VGND VGND VPWR VPWR _15838_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14476__A _13022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22644_ _22427_/X _22643_/X _15689_/B _22640_/X VGND VGND VPWR VPWR _22644_/X sky130_fd_sc_hd__o22a_4
XFILLER_41_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22693__A _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12708__B _23572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17787__A _18443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22575_ _22396_/X _22572_/X _16767_/B _22569_/X VGND VGND VPWR VPWR _23163_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21856__B2 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24314_ _24301_/CLK _19148_/X HRESETn VGND VGND VPWR VPWR _24314_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21526_ _20487_/A VGND VGND VPWR VPWR _21526_/X sky130_fd_sc_hd__buf_2
XFILLER_33_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21608__A1 _21536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24245_ _24032_/CLK _24245_/D HRESETn VGND VGND VPWR VPWR _24245_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21608__B2 _21602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21457_ _21221_/X _21456_/X _23805_/Q _21453_/X VGND VGND VPWR VPWR _21457_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12724__A _15688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17288__A1 _17283_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15100__A _15108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12190_ _13056_/A VGND VGND VPWR VPWR _12922_/A sky130_fd_sc_hd__buf_2
X_20408_ _20255_/X _20406_/X _24376_/Q _20407_/X VGND VGND VPWR VPWR _20408_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17288__B2 _17287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21084__A2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21388_ _21277_/X _21383_/X _14410_/B _21387_/X VGND VGND VPWR VPWR _21388_/X sky130_fd_sc_hd__o22a_4
X_24176_ _23104_/CLK _19760_/X HRESETn VGND VGND VPWR VPWR _14175_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22281__B2 _22276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_13_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR _24065_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__11572__A2 IRQ[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23127_ _23217_/CLK _23127_/D VGND VGND VPWR VPWR _16131_/B sky130_fd_sc_hd__dfxtp_4
X_20339_ _21795_/A VGND VGND VPWR VPWR _20339_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_76_0_HCLK clkbuf_6_38_0_HCLK/X VGND VGND VPWR VPWR _23324_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_89_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23058_ _23048_/A _23056_/X _23058_/C VGND VGND VPWR VPWR _23058_/X sky130_fd_sc_hd__and3_4
XANTENNA__22033__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15754__B _15689_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14900_ _13985_/A _14898_/X _14899_/X VGND VGND VPWR VPWR _14900_/X sky130_fd_sc_hd__and3_4
XANTENNA__22584__A2 _22579_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22009_ _22002_/A VGND VGND VPWR VPWR _22009_/X sky130_fd_sc_hd__buf_2
XANTENNA__13555__A _13500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15880_ _15892_/A _15818_/B VGND VGND VPWR VPWR _15880_/X sky130_fd_sc_hd__or2_4
XFILLER_40_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14831_ _12575_/A _14829_/X _14830_/X VGND VGND VPWR VPWR _14831_/X sky130_fd_sc_hd__and3_4
XFILLER_97_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17460__A1 _12338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17460__B2 _17459_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17550_ _17550_/A _17550_/B VGND VGND VPWR VPWR _18024_/B sky130_fd_sc_hd__or2_4
XFILLER_91_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14762_ _14758_/A _14762_/B VGND VGND VPWR VPWR _14762_/X sky130_fd_sc_hd__or2_4
X_11974_ _11974_/A VGND VGND VPWR VPWR _13957_/A sky130_fd_sc_hd__inv_2
XFILLER_99_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16501_ _16159_/X _16438_/B VGND VGND VPWR VPWR _16501_/X sky130_fd_sc_hd__or2_4
XANTENNA__17212__A1 _17182_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13713_ _13697_/X _13713_/B VGND VGND VPWR VPWR _13713_/X sky130_fd_sc_hd__or2_4
X_17481_ _13591_/X _17480_/X VGND VGND VPWR VPWR _17481_/X sky130_fd_sc_hd__or2_4
XFILLER_44_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14693_ _14664_/X _14691_/X _14692_/X VGND VGND VPWR VPWR _14693_/X sky130_fd_sc_hd__and3_4
XANTENNA__13290__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16432_ _16083_/A _16432_/B _16432_/C VGND VGND VPWR VPWR _16433_/C sky130_fd_sc_hd__and3_4
X_19220_ _19220_/A _19220_/B VGND VGND VPWR VPWR _19220_/X sky130_fd_sc_hd__and2_4
XANTENNA__11803__A _11803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13644_ _15443_/A _13727_/B VGND VGND VPWR VPWR _13644_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19151_ _19151_/A VGND VGND VPWR VPWR _19151_/Y sky130_fd_sc_hd__inv_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _13370_/A VGND VGND VPWR VPWR _16363_/X sky130_fd_sc_hd__buf_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _13574_/X VGND VGND VPWR VPWR _13575_/X sky130_fd_sc_hd__buf_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18102_ _18242_/A _18081_/A VGND VGND VPWR VPWR _18105_/C sky130_fd_sc_hd__nor2_4
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18712__A1 _18082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15314_ _15314_/A _15253_/B VGND VGND VPWR VPWR _15315_/C sky130_fd_sc_hd__or2_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12526_ _12905_/A _12643_/B VGND VGND VPWR VPWR _12527_/C sky130_fd_sc_hd__or2_4
X_19082_ _11509_/A _11508_/X _19077_/Y VGND VGND VPWR VPWR _19082_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_9_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16294_ _11959_/X _16294_/B VGND VGND VPWR VPWR _16294_/X sky130_fd_sc_hd__or2_4
XANTENNA__22108__A _22108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18033_ _17824_/A _17168_/Y _17811_/A _17185_/Y VGND VGND VPWR VPWR _18033_/X sky130_fd_sc_hd__o22a_4
X_15245_ _14246_/A _15245_/B _15245_/C VGND VGND VPWR VPWR _15245_/X sky130_fd_sc_hd__and3_4
XFILLER_9_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21012__A _21027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12457_ _12522_/A _12454_/X _12457_/C VGND VGND VPWR VPWR _12458_/C sky130_fd_sc_hd__and3_4
XANTENNA__12634__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15176_ _14992_/A _15176_/B VGND VGND VPWR VPWR _15178_/B sky130_fd_sc_hd__or2_4
X_12388_ _12388_/A _12388_/B _12388_/C VGND VGND VPWR VPWR _12389_/C sky130_fd_sc_hd__and3_4
XANTENNA__11563__A2 IRQ[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14127_ _14119_/X _14123_/X _14126_/X VGND VGND VPWR VPWR _14127_/X sky130_fd_sc_hd__or3_4
XFILLER_10_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19417__A _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19984_ _19983_/X VGND VGND VPWR VPWR _24135_/D sky130_fd_sc_hd__inv_2
XANTENNA__18321__A _18267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14058_ _14046_/A _14056_/X _14058_/C VGND VGND VPWR VPWR _14062_/B sky130_fd_sc_hd__and3_4
X_18935_ _18987_/A VGND VGND VPWR VPWR _18935_/X sky130_fd_sc_hd__buf_2
XFILLER_97_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18779__A1 _12430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13009_ _13009_/A _23282_/Q VGND VGND VPWR VPWR _13010_/C sky130_fd_sc_hd__or2_4
XANTENNA__13465__A _13437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22575__A2 _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18866_ _11599_/X _18866_/B _12068_/X _18866_/D VGND VGND VPWR VPWR _19926_/B sky130_fd_sc_hd__or4_4
XFILLER_41_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17817_ _17817_/A VGND VGND VPWR VPWR _17817_/X sky130_fd_sc_hd__buf_2
XANTENNA__17451__B2 _17664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18797_ _17171_/X _18795_/X _24426_/Q _18796_/X VGND VGND VPWR VPWR _18797_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16776__A _16800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15680__A _15812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17748_ _17748_/A _17714_/X _17747_/X VGND VGND VPWR VPWR _17748_/X sky130_fd_sc_hd__and3_4
XFILLER_93_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17203__A1 _12992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20889__A2 _20880_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17679_ _17681_/A _17487_/X VGND VGND VPWR VPWR _17757_/A sky130_fd_sc_hd__or2_4
XFILLER_36_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19418_ _19490_/A VGND VGND VPWR VPWR _19419_/A sky130_fd_sc_hd__buf_2
X_20690_ _18453_/X _20680_/X _20492_/X _20689_/Y VGND VGND VPWR VPWR _20690_/X sky130_fd_sc_hd__a211o_4
XFILLER_17_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19349_ _19347_/X _18606_/X _19347_/X _24229_/Q VGND VGND VPWR VPWR _24229_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23842__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22360_ _22110_/X _22354_/X _23279_/Q _22358_/X VGND VGND VPWR VPWR _22360_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15839__B _15839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20510__B2 _20488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21311_ _21232_/X _21305_/X _16272_/B _21309_/X VGND VGND VPWR VPWR _23897_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22291_ _22131_/X _22286_/X _14271_/B _22290_/X VGND VGND VPWR VPWR _22291_/X sky130_fd_sc_hd__o22a_4
XFILLER_11_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12544__A _12540_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21242_ _21242_/A VGND VGND VPWR VPWR _21242_/X sky130_fd_sc_hd__buf_2
X_24030_ _23774_/CLK _21066_/X VGND VGND VPWR VPWR _24030_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13359__B _13287_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12263__B _12263_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21173_ _21165_/X VGND VGND VPWR VPWR _21173_/X sky130_fd_sc_hd__buf_2
XFILLER_89_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15855__A _13546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12751__B2 _12750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20124_ _20076_/B _20123_/Y VGND VGND VPWR VPWR _20124_/X sky130_fd_sc_hd__or2_4
XANTENNA__18219__B1 _18082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22015__B2 _21970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15574__B _23787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13375__A _12837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20055_ _20042_/X _18349_/A _20048_/X _20054_/X VGND VGND VPWR VPWR _20056_/A sky130_fd_sc_hd__o22a_4
XFILLER_115_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20577__A1 _20229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24288__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23814_ _23910_/CLK _21438_/X VGND VGND VPWR VPWR _14309_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _23073_/CLK _21575_/X VGND VGND VPWR VPWR _23745_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _22458_/A VGND VGND VPWR VPWR _21574_/A sky130_fd_sc_hd__buf_2
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12719__A _12286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _16447_/A VGND VGND VPWR VPWR _16039_/A sky130_fd_sc_hd__buf_2
X_23676_ _23867_/CLK _23676_/D VGND VGND VPWR VPWR _23676_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _20888_/A VGND VGND VPWR VPWR _20888_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20936__A _22456_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22627_ _22398_/X _22622_/X _16489_/B _22626_/X VGND VGND VPWR VPWR _22627_/X sky130_fd_sc_hd__o22a_4
XFILLER_70_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20655__B _20595_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13360_ _12829_/A VGND VGND VPWR VPWR _13383_/A sky130_fd_sc_hd__buf_2
X_22558_ _22451_/X _22557_/X _14661_/B _22554_/X VGND VGND VPWR VPWR _23172_/D sky130_fd_sc_hd__o22a_4
X_12311_ _12745_/A VGND VGND VPWR VPWR _12735_/A sky130_fd_sc_hd__buf_2
X_21509_ _21506_/X _21508_/X _23773_/Q _21503_/X VGND VGND VPWR VPWR _21509_/X sky130_fd_sc_hd__o22a_4
X_13291_ _12546_/A _13291_/B VGND VGND VPWR VPWR _13291_/X sky130_fd_sc_hd__or2_4
X_22489_ _22420_/X _22486_/X _13188_/B _22483_/X VGND VGND VPWR VPWR _22489_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12454__A _12462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15030_ _15030_/A _23391_/Q VGND VGND VPWR VPWR _15031_/C sky130_fd_sc_hd__or2_4
X_12242_ _12695_/A _12236_/X _12241_/X VGND VGND VPWR VPWR _12242_/X sky130_fd_sc_hd__and3_4
X_24228_ _24229_/CLK _19351_/X HRESETn VGND VGND VPWR VPWR _20888_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21057__A2 _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15765__A _12792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12173_ _11824_/A _12169_/X _12172_/X VGND VGND VPWR VPWR _12181_/B sky130_fd_sc_hd__or3_4
X_24159_ _24293_/CLK _19889_/Y HRESETn VGND VGND VPWR VPWR _24159_/Q sky130_fd_sc_hd__dfrtp_4
X_16981_ _16947_/Y _16981_/B VGND VGND VPWR VPWR _16981_/X sky130_fd_sc_hd__or2_4
XFILLER_46_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18720_ _18390_/A _18712_/Y _18713_/X _18048_/A _18719_/X VGND VGND VPWR VPWR _18720_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15932_ _11884_/X VGND VGND VPWR VPWR _15939_/A sky130_fd_sc_hd__buf_2
XFILLER_81_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_6_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR _24473_/CLK sky130_fd_sc_hd__clkbuf_1
X_15863_ _13551_/X _15863_/B VGND VGND VPWR VPWR _15865_/B sky130_fd_sc_hd__or2_4
X_18651_ _18554_/X _18649_/X _20093_/A _18650_/X VGND VGND VPWR VPWR _24452_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14814_ _14845_/A _14743_/B VGND VGND VPWR VPWR _14815_/C sky130_fd_sc_hd__or2_4
X_17602_ _17595_/X _17602_/B VGND VGND VPWR VPWR _17602_/Y sky130_fd_sc_hd__nor2_4
X_15794_ _12851_/A _15855_/B VGND VGND VPWR VPWR _15796_/B sky130_fd_sc_hd__or2_4
X_18582_ _17336_/B _18581_/X VGND VGND VPWR VPWR _18582_/X sky130_fd_sc_hd__or2_4
XFILLER_29_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14745_ _13600_/A _14741_/X _14744_/X VGND VGND VPWR VPWR _14745_/X sky130_fd_sc_hd__or3_4
X_17533_ _17533_/A _17457_/B VGND VGND VPWR VPWR _17533_/X sky130_fd_sc_hd__and2_4
XANTENNA__21007__A _21007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11957_ _15707_/A VGND VGND VPWR VPWR _12739_/A sky130_fd_sc_hd__buf_2
XFILLER_79_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12629__A _12963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17464_ _18138_/B _17464_/B VGND VGND VPWR VPWR _17586_/C sky130_fd_sc_hd__or2_4
XANTENNA__15005__A _15028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19700__A HRDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14676_ _14714_/A _14676_/B VGND VGND VPWR VPWR _14677_/C sky130_fd_sc_hd__or2_4
X_11888_ _11888_/A _11705_/B VGND VGND VPWR VPWR _11904_/B sky130_fd_sc_hd__or2_4
XFILLER_18_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16415_ _11915_/A _16413_/X _16414_/X VGND VGND VPWR VPWR _16415_/X sky130_fd_sc_hd__and3_4
X_19203_ _19201_/X _19108_/B _19202_/Y VGND VGND VPWR VPWR _24287_/D sky130_fd_sc_hd__o21a_4
X_13627_ _13794_/A _13627_/B VGND VGND VPWR VPWR _13631_/B sky130_fd_sc_hd__or2_4
XFILLER_38_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17395_ _17179_/Y _17395_/B VGND VGND VPWR VPWR _17395_/X sky130_fd_sc_hd__or2_4
XANTENNA__14844__A _14021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16346_ _13422_/A _16342_/X _16346_/C VGND VGND VPWR VPWR _16354_/B sky130_fd_sc_hd__or3_4
X_19134_ _19134_/A _19151_/A VGND VGND VPWR VPWR _19134_/X sky130_fd_sc_hd__and2_4
X_13558_ _13558_/A _13484_/B VGND VGND VPWR VPWR _13558_/X sky130_fd_sc_hd__or2_4
XFILLER_34_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15659__B _15659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12509_ _12509_/A VGND VGND VPWR VPWR _13641_/A sky130_fd_sc_hd__buf_2
X_19065_ _19065_/A VGND VGND VPWR VPWR _19065_/Y sky130_fd_sc_hd__inv_2
X_16277_ _15936_/A _16275_/X _16277_/C VGND VGND VPWR VPWR _16277_/X sky130_fd_sc_hd__and3_4
X_13489_ _12910_/A _13487_/X _13489_/C VGND VGND VPWR VPWR _13490_/C sky130_fd_sc_hd__and3_4
XANTENNA__12364__A _13133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15228_ _14186_/A _15228_/B VGND VGND VPWR VPWR _15228_/X sky130_fd_sc_hd__or2_4
X_18016_ _18016_/A VGND VGND VPWR VPWR _18016_/X sky130_fd_sc_hd__buf_2
XANTENNA__22245__B2 _22240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23245__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12083__B _23901_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15675__A _12709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15159_ _14096_/X _15159_/B VGND VGND VPWR VPWR _15159_/X sky130_fd_sc_hd__or2_4
XFILLER_102_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19967_ _17885_/X _19961_/X _19966_/Y _19957_/X VGND VGND VPWR VPWR _19967_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22548__A2 _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13195__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18918_ _15249_/X _18912_/X _19098_/A _18913_/X VGND VGND VPWR VPWR _24353_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11708__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19413__A2 _24191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19898_ _22932_/A VGND VGND VPWR VPWR _19909_/A sky130_fd_sc_hd__buf_2
XFILLER_60_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18849_ _18842_/A VGND VGND VPWR VPWR _18849_/X sky130_fd_sc_hd__buf_2
XFILLER_110_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24310__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21860_ _21859_/X _21853_/X _23585_/Q _21787_/X VGND VGND VPWR VPWR _23585_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20811_ _20715_/A _20811_/B VGND VGND VPWR VPWR _20811_/Y sky130_fd_sc_hd__nor2_4
XFILLER_93_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21791_ _21791_/A VGND VGND VPWR VPWR _21791_/X sky130_fd_sc_hd__buf_2
XANTENNA__17188__B1 _15782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23530_ _23915_/CLK _23530_/D VGND VGND VPWR VPWR _23530_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20742_ _18506_/X _20680_/X _20731_/X _20741_/Y VGND VGND VPWR VPWR _20742_/X sky130_fd_sc_hd__a211o_4
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23461_ _23365_/CLK _23461_/D VGND VGND VPWR VPWR _14476_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20673_ _20444_/A VGND VGND VPWR VPWR _20673_/X sky130_fd_sc_hd__buf_2
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22412_ _22410_/X _22404_/X _12564_/B _22411_/X VGND VGND VPWR VPWR _23253_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22484__A1 _22410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23392_ _24032_/CLK _22198_/X VGND VGND VPWR VPWR _14899_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22484__B2 _22483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15569__B _23211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22343_ _22081_/X _22340_/X _16759_/B _22337_/X VGND VGND VPWR VPWR _23291_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12274__A _12710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14174__B1 _11594_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21039__A2 _21037_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21587__A _21602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22274_ _22103_/X _22272_/X _13069_/B _22269_/X VGND VGND VPWR VPWR _23346_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24170__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24013_ _23698_/CLK _21091_/X VGND VGND VPWR VPWR _15855_/B sky130_fd_sc_hd__dfxtp_4
X_21225_ _21795_/A VGND VGND VPWR VPWR _21225_/X sky130_fd_sc_hd__buf_2
XANTENNA__15585__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19057__A _19027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20798__A1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20798__B2 _20724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21156_ _20916_/X _21154_/X _14811_/B _21151_/X VGND VGND VPWR VPWR _23971_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22539__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20107_ _11626_/Y _20106_/X _11625_/X _18668_/Y VGND VGND VPWR VPWR _20107_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11618__A _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21087_ _20591_/X _21082_/X _24016_/Q _21086_/X VGND VGND VPWR VPWR _21087_/X sky130_fd_sc_hd__o22a_4
XFILLER_63_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21747__B1 _16368_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20038_ _24461_/Q VGND VGND VPWR VPWR _20038_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14929__A _13998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13833__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12860_ _12860_/A VGND VGND VPWR VPWR _12861_/A sky130_fd_sc_hd__buf_2
XFILLER_2_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11811_ _11717_/X _23838_/Q VGND VGND VPWR VPWR _11811_/X sky130_fd_sc_hd__or2_4
XFILLER_76_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12791_ _12791_/A VGND VGND VPWR VPWR _12792_/A sky130_fd_sc_hd__buf_2
XFILLER_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ _21816_/X _21988_/X _23507_/Q _21985_/X VGND VGND VPWR VPWR _21989_/X sky130_fd_sc_hd__o22a_4
XFILLER_42_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23118__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18915__A1 _17297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _12612_/A _14522_/X _14529_/X VGND VGND VPWR VPWR _14531_/C sky130_fd_sc_hd__and3_4
XANTENNA__22711__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11741_/X VGND VGND VPWR VPWR _13370_/A sky130_fd_sc_hd__buf_2
X_23728_ _23157_/CLK _21610_/X VGND VGND VPWR VPWR _23728_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12168__B _23805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _13056_/A _14438_/X _14445_/X _14452_/X _14460_/X VGND VGND VPWR VPWR _14461_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _12787_/A VGND VGND VPWR VPWR _11673_/X sky130_fd_sc_hd__buf_2
X_23659_ _23688_/CLK _23659_/D VGND VGND VPWR VPWR _23659_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14664__A _14246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _11666_/X _16200_/B _16200_/C VGND VGND VPWR VPWR _16232_/B sky130_fd_sc_hd__or3_4
XFILLER_74_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18136__A _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13376_/X _23696_/Q VGND VGND VPWR VPWR _13414_/B sky130_fd_sc_hd__or2_4
XANTENNA__17040__A _17040_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17180_ _17179_/Y _17161_/X _12676_/X _17157_/X VGND VGND VPWR VPWR _17180_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18679__B1 _18674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ _15592_/A _14390_/X _14392_/C VGND VGND VPWR VPWR _14392_/X sky130_fd_sc_hd__and3_4
XANTENNA__22475__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16131_ _16127_/A _16131_/B VGND VGND VPWR VPWR _16131_/X sky130_fd_sc_hd__or2_4
X_13343_ _15784_/A _23696_/Q VGND VGND VPWR VPWR _13343_/X sky130_fd_sc_hd__or2_4
XANTENNA__16154__A1 _11982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16062_ _16050_/A _23800_/Q VGND VGND VPWR VPWR _16062_/X sky130_fd_sc_hd__or2_4
XANTENNA__24327__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13274_ _13135_/X VGND VGND VPWR VPWR _13274_/X sky130_fd_sc_hd__buf_2
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17694__B _17367_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22227__B2 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15013_ _15013_/A _23135_/Q VGND VGND VPWR VPWR _15015_/B sky130_fd_sc_hd__or2_4
XANTENNA__12715__A1 _12682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12225_ _12688_/A _12222_/X _12224_/X VGND VGND VPWR VPWR _12225_/X sky130_fd_sc_hd__and3_4
XANTENNA__15495__A _15495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21986__B1 _12571_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19821_ _19670_/X _19817_/X _19820_/Y VGND VGND VPWR VPWR _19829_/B sky130_fd_sc_hd__o21a_4
XFILLER_64_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12156_ _11734_/A _24061_/Q VGND VGND VPWR VPWR _12157_/C sky130_fd_sc_hd__or2_4
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24139__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_46_0_HCLK clkbuf_5_23_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16103__B _16103_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19752_ _19712_/A HRDATA[2] VGND VGND VPWR VPWR _19752_/X sky130_fd_sc_hd__and2_4
X_12087_ _12065_/X _24061_/Q VGND VGND VPWR VPWR _12088_/C sky130_fd_sc_hd__or2_4
X_16964_ _16964_/A VGND VGND VPWR VPWR _16965_/C sky130_fd_sc_hd__inv_2
XFILLER_77_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18703_ _16933_/A _18700_/X _16931_/X _18702_/X VGND VGND VPWR VPWR _18703_/Y sky130_fd_sc_hd__a22oi_4
X_15915_ _15914_/A _15914_/B VGND VGND VPWR VPWR _15915_/X sky130_fd_sc_hd__or2_4
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21202__A2 _21197_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19683_ _19784_/B _19754_/A VGND VGND VPWR VPWR _19683_/X sky130_fd_sc_hd__or2_4
XFILLER_76_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16895_ _17054_/A VGND VGND VPWR VPWR _16907_/C sky130_fd_sc_hd__buf_2
XANTENNA__14839__A _14815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13743__A _13711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18634_ _18418_/A _17306_/A VGND VGND VPWR VPWR _18634_/Y sky130_fd_sc_hd__nor2_4
X_15846_ _12386_/X _23501_/Q VGND VGND VPWR VPWR _15847_/C sky130_fd_sc_hd__or2_4
XFILLER_18_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14558__B _14480_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18565_ _17103_/X _18141_/Y _17933_/A _18564_/Y VGND VGND VPWR VPWR _18565_/X sky130_fd_sc_hd__a211o_4
X_12989_ _12989_/A _12957_/X _12988_/X VGND VGND VPWR VPWR _12989_/X sky130_fd_sc_hd__and3_4
X_15777_ _12672_/A _15761_/X _15776_/X VGND VGND VPWR VPWR _15777_/X sky130_fd_sc_hd__or3_4
XFILLER_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12359__A _13243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22163__B1 _16424_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14640__A1 _11841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22702__A2 _22700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_HCLK clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17516_ _13575_/X _17480_/X VGND VGND VPWR VPWR _17516_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__19430__A _16997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14728_ _14158_/A _14790_/B VGND VGND VPWR VPWR _14728_/X sky130_fd_sc_hd__or2_4
XFILLER_75_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18496_ _17968_/X _18250_/X VGND VGND VPWR VPWR _18496_/Y sky130_fd_sc_hd__nor2_4
XFILLER_36_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20713__A1 _20518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20576__A _20285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20713__B2 _20525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12078__B _12140_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14659_ _13708_/A VGND VGND VPWR VPWR _14925_/A sky130_fd_sc_hd__buf_2
X_17447_ _17447_/A _17446_/X VGND VGND VPWR VPWR _17447_/X sky130_fd_sc_hd__or2_4
XANTENNA__21269__A2 _21259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17378_ _17377_/X VGND VGND VPWR VPWR _17380_/A sky130_fd_sc_hd__inv_2
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14293__B _14293_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19117_ _24296_/Q _19117_/B VGND VGND VPWR VPWR _19118_/B sky130_fd_sc_hd__and2_4
X_16329_ _16447_/A _16329_/B _16329_/C VGND VGND VPWR VPWR _16330_/C sky130_fd_sc_hd__and3_4
X_19048_ _24330_/Q _11515_/B _19042_/Y VGND VGND VPWR VPWR _19048_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_118_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13918__A _13918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12822__A _12822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21010_ _21009_/X VGND VGND VPWR VPWR _21015_/A sky130_fd_sc_hd__buf_2
XANTENNA__21441__A2 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19398__B2 _24202_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22961_ _22961_/A VGND VGND VPWR VPWR HADDR[13] sky130_fd_sc_hd__inv_2
XANTENNA__15852__B _15852_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22031__A _22031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14749__A _13959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21912_ _21859_/X _21908_/X _23553_/Q _21869_/X VGND VGND VPWR VPWR _21912_/X sky130_fd_sc_hd__o22a_4
X_22892_ _19901_/X _18681_/A _23048_/A VGND VGND VPWR VPWR _22892_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20952__A1 _18700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21870__A _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21843_ _21843_/A VGND VGND VPWR VPWR _21843_/X sky130_fd_sc_hd__buf_2
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12269__A _12269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19340__A _19336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21774_ _21562_/X _21769_/X _14324_/B _21773_/X VGND VGND VPWR VPWR _21774_/X sky130_fd_sc_hd__o22a_4
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20486__A _20486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23513_ _23514_/CLK _23513_/D VGND VGND VPWR VPWR _23513_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23410__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20725_ _20613_/X _20723_/X _24075_/Q _20724_/X VGND VGND VPWR VPWR _24075_/D sky130_fd_sc_hd__o22a_4
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14484__A _13620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23444_ _23699_/CLK _23444_/D VGND VGND VPWR VPWR _12711_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20656_ _20656_/A VGND VGND VPWR VPWR _20657_/A sky130_fd_sc_hd__inv_2
XANTENNA__22457__B2 _22447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19322__B2 _20414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23375_ _23311_/CLK _23375_/D VGND VGND VPWR VPWR _13552_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_20_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20587_ _20444_/X _20577_/Y _20585_/X _20586_/Y _20459_/X VGND VGND VPWR VPWR _20588_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23560__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22326_ _14682_/B VGND VGND VPWR VPWR _22326_/X sky130_fd_sc_hd__buf_2
XANTENNA__22209__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21680__A2 _21676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13828__A _15443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22257_ _22286_/A VGND VGND VPWR VPWR _22272_/A sky130_fd_sc_hd__buf_2
XFILLER_105_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12732__A _12706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12010_ _16536_/A _24094_/Q VGND VGND VPWR VPWR _12011_/C sky130_fd_sc_hd__or2_4
X_21208_ _20958_/X _21204_/X _15156_/B _21165_/X VGND VGND VPWR VPWR _23937_/D sky130_fd_sc_hd__o22a_4
XFILLER_117_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21432__A2 _21426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22188_ _22127_/X _22186_/X _23400_/Q _22183_/X VGND VGND VPWR VPWR _22188_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21139_ _20611_/X _21133_/X _13531_/B _21137_/X VGND VGND VPWR VPWR _23983_/D sky130_fd_sc_hd__o22a_4
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13961_ _13611_/A _13959_/X _13961_/C VGND VGND VPWR VPWR _13961_/X sky130_fd_sc_hd__and3_4
XFILLER_8_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23037__A _22968_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14659__A _13708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21196__B2 _21194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12912_ _12500_/X _12912_/B VGND VGND VPWR VPWR _12913_/C sky130_fd_sc_hd__or2_4
X_15700_ _12739_/A _15700_/B VGND VGND VPWR VPWR _15701_/C sky130_fd_sc_hd__or2_4
XFILLER_78_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16680_ _16596_/Y _16678_/X VGND VGND VPWR VPWR _16681_/A sky130_fd_sc_hd__or2_4
XFILLER_100_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13892_ _13880_/A _13892_/B _13892_/C VGND VGND VPWR VPWR _13893_/C sky130_fd_sc_hd__and3_4
XFILLER_73_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14378__B _14283_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12843_ _12752_/Y _12841_/X VGND VGND VPWR VPWR _12843_/X sky130_fd_sc_hd__or2_4
X_15631_ _15631_/A _15629_/X _15630_/X VGND VGND VPWR VPWR _15635_/B sky130_fd_sc_hd__and3_4
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13282__B _13282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15562_ _15536_/A _23371_/Q VGND VGND VPWR VPWR _15562_/X sky130_fd_sc_hd__or2_4
X_18350_ _18459_/A _18350_/B VGND VGND VPWR VPWR _18351_/B sky130_fd_sc_hd__or2_4
X_12774_ _12816_/A _12774_/B VGND VGND VPWR VPWR _12775_/C sky130_fd_sc_hd__or2_4
XANTENNA__17689__B _17469_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22696__B2 _22690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20396__A _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23090__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _11740_/A _14507_/X _14512_/X VGND VGND VPWR VPWR _14513_/X sky130_fd_sc_hd__or3_4
X_17301_ _17298_/Y _17010_/X _17018_/A _17300_/X VGND VGND VPWR VPWR _17302_/A sky130_fd_sc_hd__o22a_4
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _13214_/A VGND VGND VPWR VPWR _15743_/A sky130_fd_sc_hd__buf_2
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _15493_/A _15493_/B VGND VGND VPWR VPWR _15495_/B sky130_fd_sc_hd__or2_4
X_18281_ _18281_/A _18280_/X VGND VGND VPWR VPWR _18281_/X sky130_fd_sc_hd__or2_4
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12907__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11811__A _11717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _12862_/A _14444_/B _14444_/C VGND VGND VPWR VPWR _14445_/C sky130_fd_sc_hd__and3_4
X_17232_ _16376_/X _17100_/X _14723_/B _17065_/X VGND VGND VPWR VPWR _17232_/X sky130_fd_sc_hd__o22a_4
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11656_/A VGND VGND VPWR VPWR _12989_/A sky130_fd_sc_hd__buf_2
XANTENNA__22448__B2 _22447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18116__A2 _17982_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17163_ _17163_/A VGND VGND VPWR VPWR _17163_/X sky130_fd_sc_hd__buf_2
XFILLER_80_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14375_ _15637_/A _14296_/B VGND VGND VPWR VPWR _14376_/C sky130_fd_sc_hd__or2_4
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _11634_/A _11634_/B _17009_/A _17024_/B VGND VGND VPWR VPWR _11591_/C sky130_fd_sc_hd__or4_4
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21120__B2 _21116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16114_ _16091_/A _16181_/B VGND VGND VPWR VPWR _16116_/B sky130_fd_sc_hd__or2_4
XFILLER_10_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13326_ _13301_/A _13326_/B VGND VGND VPWR VPWR _13326_/X sky130_fd_sc_hd__or2_4
XFILLER_116_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17875__A1 _17874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17094_ _18103_/A VGND VGND VPWR VPWR _18421_/A sky130_fd_sc_hd__buf_2
XANTENNA__21671__A2 _21669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16045_ _16045_/A _16045_/B _16044_/X VGND VGND VPWR VPWR _16077_/B sky130_fd_sc_hd__or3_4
XANTENNA__21020__A _21012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13257_ _13257_/A _13257_/B VGND VGND VPWR VPWR _13258_/C sky130_fd_sc_hd__or2_4
XFILLER_89_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12208_ _13984_/A VGND VGND VPWR VPWR _12209_/A sky130_fd_sc_hd__buf_2
X_13188_ _15784_/A _13188_/B VGND VGND VPWR VPWR _13188_/X sky130_fd_sc_hd__or2_4
XANTENNA__22620__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19804_ _19813_/A _19802_/X _19803_/X VGND VGND VPWR VPWR _19804_/X sky130_fd_sc_hd__and3_4
X_12139_ _11827_/A _12139_/B VGND VGND VPWR VPWR _12139_/X sky130_fd_sc_hd__or2_4
XANTENNA__19425__A _19416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17996_ _17569_/A _17995_/X VGND VGND VPWR VPWR _17996_/X sky130_fd_sc_hd__or2_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19735_ HRDATA[20] VGND VGND VPWR VPWR _20895_/B sky130_fd_sc_hd__buf_2
X_16947_ _24129_/Q VGND VGND VPWR VPWR _16947_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19666_ _19607_/X _19657_/X _19663_/Y _19665_/X VGND VGND VPWR VPWR _19667_/B sky130_fd_sc_hd__a211o_4
X_16878_ _12680_/B _16826_/X _12680_/B _16826_/X VGND VGND VPWR VPWR _16879_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22786__A _17109_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18617_ _18614_/Y _18615_/X VGND VGND VPWR VPWR _18617_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__23433__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21690__A _21690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15829_ _12477_/X _15829_/B VGND VGND VPWR VPWR _15829_/X sky130_fd_sc_hd__or2_4
XFILLER_0_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19597_ _19597_/A VGND VGND VPWR VPWR _19876_/B sky130_fd_sc_hd__inv_2
XFILLER_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18548_ _18487_/X _18540_/Y _18541_/X _18543_/X _18547_/Y VGND VGND VPWR VPWR _18548_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_52_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22687__B2 _22683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18479_ _18435_/X _18478_/X _24459_/Q _18435_/X VGND VGND VPWR VPWR _18479_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12817__A _12754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20510_ _20396_/X _20509_/X _24084_/Q _20488_/X VGND VGND VPWR VPWR _24084_/D sky130_fd_sc_hd__o22a_4
XFILLER_53_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11721__A _13708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21490_ _21280_/X _21484_/X _14484_/B _21488_/X VGND VGND VPWR VPWR _23781_/D sky130_fd_sc_hd__o22a_4
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20441_ _20441_/A VGND VGND VPWR VPWR _20442_/A sky130_fd_sc_hd__buf_2
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19855__A2 _19689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14129__B1 _14118_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23160_ _23383_/CLK _23160_/D VGND VGND VPWR VPWR _15967_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_88_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20372_ _20372_/A VGND VGND VPWR VPWR _21799_/A sky130_fd_sc_hd__buf_2
XFILLER_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22111_ _22110_/X _22101_/X _13457_/B _22108_/X VGND VGND VPWR VPWR _22111_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13648__A _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23091_ _23859_/CLK _22687_/X VGND VGND VPWR VPWR _23091_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12552__A _13014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24373__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22042_ _22035_/A VGND VGND VPWR VPWR _22042_/X sky130_fd_sc_hd__buf_2
XFILLER_47_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21414__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13367__B _24016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22611__B2 _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12271__B _12271_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15863__A _13551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19335__A _19317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23993_ _23514_/CLK _23993_/D VGND VGND VPWR VPWR _23993_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14479__A _13022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21178__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22944_ _22962_/A _22944_/B VGND VGND VPWR VPWR _22946_/B sky130_fd_sc_hd__nand2_4
XFILLER_99_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20925__B2 _20449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14198__B _24009_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22875_ _22872_/A _22875_/B VGND VGND VPWR VPWR HWDATA[29] sky130_fd_sc_hd__nor2_4
XFILLER_83_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21826_ _21256_/A VGND VGND VPWR VPWR _21826_/X sky130_fd_sc_hd__buf_2
XANTENNA__22678__A1 _21802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22678__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21757_ _21534_/X _21755_/X _13046_/B _21752_/X VGND VGND VPWR VPWR _23634_/D sky130_fd_sc_hd__o22a_4
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12727__A _15664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11510_ _24325_/Q _11510_/B VGND VGND VPWR VPWR _11511_/B sky130_fd_sc_hd__or2_4
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20708_ _20708_/A _20708_/B VGND VGND VPWR VPWR _20708_/X sky130_fd_sc_hd__or2_4
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _13020_/A VGND VGND VPWR VPWR _13009_/A sky130_fd_sc_hd__buf_2
X_24476_ _24229_/CLK _24476_/D HRESETn VGND VGND VPWR VPWR _24476_/Q sky130_fd_sc_hd__dfrtp_4
X_21688_ _21687_/X VGND VGND VPWR VPWR _21688_/X sky130_fd_sc_hd__buf_2
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23427_ _23907_/CLK _22140_/X VGND VGND VPWR VPWR _14806_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20639_ _20421_/A VGND VGND VPWR VPWR _20639_/X sky130_fd_sc_hd__buf_2
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14942__A _15074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21102__B2 _21100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14160_ _15030_/A VGND VGND VPWR VPWR _14161_/A sky130_fd_sc_hd__buf_2
X_23358_ _23358_/CLK _22256_/X VGND VGND VPWR VPWR _11732_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22850__A1 _17283_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21653__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13111_ _13104_/A _13111_/B VGND VGND VPWR VPWR _13111_/X sky130_fd_sc_hd__or2_4
X_22309_ _23317_/Q VGND VGND VPWR VPWR _23317_/D sky130_fd_sc_hd__buf_2
X_14091_ _11606_/A VGND VGND VPWR VPWR _14991_/A sky130_fd_sc_hd__buf_2
XFILLER_4_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23289_ _23354_/CLK _22346_/X VGND VGND VPWR VPWR _16253_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23306__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12462__A _12462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_111_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR _23827_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_106_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13042_ _13015_/A _23474_/Q VGND VGND VPWR VPWR _13044_/B sky130_fd_sc_hd__or2_4
XFILLER_45_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22602__B2 _22597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15773__A _12795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17850_ _17812_/A _17250_/X _17800_/A _17849_/Y VGND VGND VPWR VPWR _17850_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16801_ _16616_/A _16799_/X _16800_/X VGND VGND VPWR VPWR _16802_/C sky130_fd_sc_hd__and3_4
XFILLER_8_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23456__CLK _23840_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17781_ _18205_/A _17781_/B VGND VGND VPWR VPWR _17789_/B sky130_fd_sc_hd__and2_4
X_14993_ _14997_/A _23711_/Q VGND VGND VPWR VPWR _14994_/C sky130_fd_sc_hd__or2_4
XANTENNA__14389__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19520_ _24148_/Q _19459_/X HRDATA[22] _19460_/X VGND VGND VPWR VPWR _19520_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13293__A _12540_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16732_ _12100_/X _16730_/X _16732_/C VGND VGND VPWR VPWR _16732_/X sky130_fd_sc_hd__and3_4
X_13944_ _13968_/A _13942_/X _13943_/X VGND VGND VPWR VPWR _13944_/X sky130_fd_sc_hd__and3_4
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19451_ HRDATA[31] VGND VGND VPWR VPWR _20224_/B sky130_fd_sc_hd__buf_2
X_13875_ _13910_/A _13875_/B VGND VGND VPWR VPWR _13876_/C sky130_fd_sc_hd__or2_4
X_16663_ _16651_/A _23804_/Q VGND VGND VPWR VPWR _16664_/C sky130_fd_sc_hd__or2_4
X_18402_ _17382_/B _18401_/X _17432_/X VGND VGND VPWR VPWR _18402_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12826_ _12826_/A VGND VGND VPWR VPWR _12827_/A sky130_fd_sc_hd__buf_2
X_15614_ _15614_/A _23883_/Q VGND VGND VPWR VPWR _15614_/X sky130_fd_sc_hd__or2_4
X_19382_ _19382_/A VGND VGND VPWR VPWR _19382_/Y sky130_fd_sc_hd__inv_2
X_16594_ _11992_/X _16570_/X _16577_/X _16585_/X _16593_/X VGND VGND VPWR VPWR _16594_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_91_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18333_ _18332_/A _18331_/X _18160_/X VGND VGND VPWR VPWR _18333_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21015__A _21015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12757_ _13129_/A VGND VGND VPWR VPWR _12808_/A sky130_fd_sc_hd__buf_2
X_15545_ _15578_/A _15543_/X _15545_/C VGND VGND VPWR VPWR _15545_/X sky130_fd_sc_hd__and3_4
XFILLER_72_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12082__A1 _12036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12637__A _12957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21341__A1 _21282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16109__A _16109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21341__B2 _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11708_/A VGND VGND VPWR VPWR _11709_/A sky130_fd_sc_hd__buf_2
X_15476_ _12613_/A _15472_/X _15475_/X VGND VGND VPWR VPWR _15476_/X sky130_fd_sc_hd__or3_4
X_18264_ _18264_/A _17515_/Y VGND VGND VPWR VPWR _18267_/B sky130_fd_sc_hd__and2_4
X_12688_ _12688_/A _12686_/X _12687_/X VGND VGND VPWR VPWR _12689_/C sky130_fd_sc_hd__and3_4
XANTENNA__21892__A2 _21887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ _15389_/A VGND VGND VPWR VPWR _14427_/Y sky130_fd_sc_hd__inv_2
X_17215_ _17151_/X _17211_/X _17160_/X _17214_/X VGND VGND VPWR VPWR _17215_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_106_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11639_ _13686_/A VGND VGND VPWR VPWR _15611_/A sky130_fd_sc_hd__buf_2
XFILLER_50_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15948__A _15948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18195_ _17756_/Y _18166_/X _17756_/Y _18166_/X VGND VGND VPWR VPWR _18195_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18253__A1_N _18189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14852__A _14851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ _14371_/A VGND VGND VPWR VPWR _15607_/A sky130_fd_sc_hd__buf_2
X_17146_ _17143_/X _17161_/A _17144_/Y _17145_/X VGND VGND VPWR VPWR _17146_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22841__A1 _14786_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21644__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15667__B _15667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13309_ _15667_/A _23568_/Q VGND VGND VPWR VPWR _13309_/X sky130_fd_sc_hd__or2_4
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13468__A _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20852__B1 _20844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17077_ _17077_/A _18203_/A VGND VGND VPWR VPWR _17077_/X sky130_fd_sc_hd__or2_4
X_14289_ _15556_/A _14289_/B VGND VGND VPWR VPWR _14290_/C sky130_fd_sc_hd__or2_4
XFILLER_115_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24231__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16028_ _11745_/X _16028_/B _16028_/C VGND VGND VPWR VPWR _16029_/C sky130_fd_sc_hd__or3_4
XANTENNA__12091__B _23837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16779__A _16624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15683__A _12240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19470__B1 HRDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_16_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_97_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17979_ _17926_/X _17976_/Y _17921_/X _17978_/Y VGND VGND VPWR VPWR _17979_/X sky130_fd_sc_hd__o22a_4
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14299__A _12269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18994__A _18994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19718_ _19718_/A _19718_/B VGND VGND VPWR VPWR _19880_/B sky130_fd_sc_hd__and2_4
X_20990_ _24383_/Q _20405_/A _11540_/A _20449_/A VGND VGND VPWR VPWR _20990_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19773__A1 _19722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19649_ HRDATA[25] VGND VGND VPWR VPWR _20400_/B sky130_fd_sc_hd__buf_2
XFILLER_4_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13931__A _13960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22660_ _22456_/X _22657_/X _15289_/B _22654_/X VGND VGND VPWR VPWR _23106_/D sky130_fd_sc_hd__o22a_4
XFILLER_94_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21611_ _21541_/X _21605_/X _13504_/B _21609_/X VGND VGND VPWR VPWR _23727_/D sky130_fd_sc_hd__o22a_4
X_22591_ _22422_/X _22586_/X _13311_/B _22590_/X VGND VGND VPWR VPWR _23152_/D sky130_fd_sc_hd__o22a_4
XFILLER_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21332__B2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24330_ _24330_/CLK _24330_/D HRESETn VGND VGND VPWR VPWR _24330_/Q sky130_fd_sc_hd__dfstp_4
X_21542_ _21541_/X _21532_/X _13435_/B _21539_/X VGND VGND VPWR VPWR _23759_/D sky130_fd_sc_hd__o22a_4
XFILLER_33_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24261_ _24305_/CLK _24261_/D HRESETn VGND VGND VPWR VPWR _24261_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_5_16_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15858__A _15882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21473_ _21251_/X _21470_/X _13254_/B _21467_/X VGND VGND VPWR VPWR _23793_/D sky130_fd_sc_hd__o22a_4
XFILLER_53_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23212_ _23404_/CLK _23212_/D VGND VGND VPWR VPWR _15511_/B sky130_fd_sc_hd__dfxtp_4
X_20424_ _20424_/A VGND VGND VPWR VPWR _20424_/X sky130_fd_sc_hd__buf_2
X_24192_ _24203_/CLK _24192_/D HRESETn VGND VGND VPWR VPWR _24192_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22832__A1 _15120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15577__B _15577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23143_ _23847_/CLK _22603_/X VGND VGND VPWR VPWR _13873_/B sky130_fd_sc_hd__dfxtp_4
X_20355_ _20355_/A VGND VGND VPWR VPWR _21797_/A sky130_fd_sc_hd__buf_2
XFILLER_84_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12282__A _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21595__A _21595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23074_ _23522_/CLK _23074_/D VGND VGND VPWR VPWR _15303_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23479__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20286_ _20286_/A VGND VGND VPWR VPWR _20286_/X sky130_fd_sc_hd__buf_2
XFILLER_103_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22025_ _21791_/X _22024_/X _23485_/Q _22021_/X VGND VGND VPWR VPWR _23485_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22060__A2 _22059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19461__B1 HRDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22348__B1 _15952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11990_ _11982_/X _11990_/B VGND VGND VPWR VPWR _11990_/X sky130_fd_sc_hd__and2_4
X_23976_ _24008_/CLK _23976_/D VGND VGND VPWR VPWR _13630_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14002__A _14002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22927_ _22998_/A _22927_/B VGND VGND VPWR VPWR _22927_/X sky130_fd_sc_hd__or2_4
XFILLER_84_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21571__B2 _21563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13660_ _15429_/A _13660_/B VGND VGND VPWR VPWR _13660_/X sky130_fd_sc_hd__or2_4
XANTENNA__17313__A _14429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22858_ _22813_/X _22858_/B VGND VGND VPWR VPWR HWDATA[24] sky130_fd_sc_hd__nor2_4
XFILLER_72_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_36_0_HCLK clkbuf_6_18_0_HCLK/X VGND VGND VPWR VPWR _23973_/CLK sky130_fd_sc_hd__clkbuf_1
X_12611_ _13901_/A VGND VGND VPWR VPWR _12612_/A sky130_fd_sc_hd__buf_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21809_ _20464_/A VGND VGND VPWR VPWR _21809_/X sky130_fd_sc_hd__buf_2
XFILLER_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13591_ _13577_/B VGND VGND VPWR VPWR _13591_/X sky130_fd_sc_hd__buf_2
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17032__B _17032_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22789_ _14493_/Y _22781_/X VGND VGND VPWR VPWR HWDATA[6] sky130_fd_sc_hd__nor2_4
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12457__A _12522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_99_0_HCLK clkbuf_6_49_0_HCLK/X VGND VGND VPWR VPWR _23313_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15330_ _14008_/A _15330_/B _15329_/X VGND VGND VPWR VPWR _15330_/X sky130_fd_sc_hd__or3_4
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12542_ _12497_/X _12542_/B VGND VGND VPWR VPWR _12542_/X sky130_fd_sc_hd__or2_4
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15261_ _11909_/A _15259_/X _15260_/X VGND VGND VPWR VPWR _15265_/B sky130_fd_sc_hd__and3_4
XANTENNA__15768__A _11680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12473_ _12472_/X VGND VGND VPWR VPWR _13799_/A sky130_fd_sc_hd__buf_2
X_24459_ _24126_/CLK _18479_/X HRESETn VGND VGND VPWR VPWR _24459_/Q sky130_fd_sc_hd__dfrtp_4
X_14212_ _14367_/A _14212_/B _14211_/X VGND VGND VPWR VPWR _14212_/X sky130_fd_sc_hd__or3_4
X_17000_ _17000_/A VGND VGND VPWR VPWR _17001_/C sky130_fd_sc_hd__inv_2
XANTENNA__21087__B1 _24016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15192_ _14642_/A _15188_/X _15192_/C VGND VGND VPWR VPWR _15200_/B sky130_fd_sc_hd__or3_4
XFILLER_32_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14391__B _14302_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_HCLK clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_3_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_14143_ _14143_/A _23401_/Q VGND VGND VPWR VPWR _14144_/C sky130_fd_sc_hd__or2_4
XFILLER_4_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12192__A _15412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13316__A1 _13491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14074_ _14074_/A _14073_/X VGND VGND VPWR VPWR _14074_/X sky130_fd_sc_hd__and2_4
X_18951_ _18941_/X _18949_/X _18950_/Y _18946_/X VGND VGND VPWR VPWR _18951_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22587__B1 _12945_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13025_ _13025_/A _13021_/X _13024_/X VGND VGND VPWR VPWR _13026_/B sky130_fd_sc_hd__or3_4
X_17902_ _18442_/A _17902_/B VGND VGND VPWR VPWR _17902_/X sky130_fd_sc_hd__and2_4
XFILLER_80_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18882_ _17277_/X _18875_/X _24379_/Q _18878_/X VGND VGND VPWR VPWR _24379_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12920__A _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22051__A2 _22045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17833_ _17824_/X _17829_/Y _17812_/A _17832_/Y VGND VGND VPWR VPWR _17833_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15008__A _14748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17764_ _17764_/A VGND VGND VPWR VPWR _17764_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14976_ _14642_/A _14976_/B _14976_/C VGND VGND VPWR VPWR _14984_/B sky130_fd_sc_hd__or3_4
XFILLER_82_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19503_ _19464_/Y VGND VGND VPWR VPWR _19719_/A sky130_fd_sc_hd__buf_2
XFILLER_63_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16715_ _16715_/A _16715_/B _16715_/C VGND VGND VPWR VPWR _16719_/B sky130_fd_sc_hd__and3_4
X_13927_ _13927_/A _23498_/Q VGND VGND VPWR VPWR _13928_/C sky130_fd_sc_hd__or2_4
X_17695_ _17699_/A _17375_/X VGND VGND VPWR VPWR _17696_/B sky130_fd_sc_hd__or2_4
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20365__A2 _20364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18319__A _18206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14847__A _14847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13751__A _12935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19434_ _19433_/Y VGND VGND VPWR VPWR _19435_/A sky130_fd_sc_hd__buf_2
X_16646_ _16045_/A _16646_/B _16646_/C VGND VGND VPWR VPWR _16646_/X sky130_fd_sc_hd__or3_4
XFILLER_63_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13858_ _14499_/A _13858_/B _13858_/C VGND VGND VPWR VPWR _13858_/X sky130_fd_sc_hd__and3_4
XFILLER_62_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14566__B _14565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13470__B _23823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12809_ _12816_/A _23956_/Q VGND VGND VPWR VPWR _12810_/C sky130_fd_sc_hd__or2_4
X_19365_ _19359_/X _19364_/X _19359_/X _24222_/Q VGND VGND VPWR VPWR _19365_/X sky130_fd_sc_hd__a2bb2o_4
X_16577_ _16689_/A _16577_/B _16577_/C VGND VGND VPWR VPWR _16577_/X sky130_fd_sc_hd__or3_4
XANTENNA__12367__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13789_ _15404_/A _13787_/X _13789_/C VGND VGND VPWR VPWR _13790_/C sky130_fd_sc_hd__and3_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21314__B2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18316_ _18233_/B _22979_/B _18233_/B _22979_/B VGND VGND VPWR VPWR _18316_/X sky130_fd_sc_hd__a2bb2o_4
X_15528_ _11859_/A _15524_/X _15527_/X VGND VGND VPWR VPWR _15528_/X sky130_fd_sc_hd__or3_4
X_19296_ _19205_/A _19205_/B _19295_/Y VGND VGND VPWR VPWR _24256_/D sky130_fd_sc_hd__o21a_4
X_18247_ _18040_/X _18246_/X _18183_/X _17963_/X VGND VGND VPWR VPWR _18248_/A sky130_fd_sc_hd__o22a_4
XFILLER_31_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15678__A _12744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15459_ _12585_/A _15459_/B VGND VGND VPWR VPWR _15459_/X sky130_fd_sc_hd__or2_4
XANTENNA__14582__A _15015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21078__B1 _12236_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21617__A2 _21612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18178_ _18242_/A _17473_/X VGND VGND VPWR VPWR _18180_/C sky130_fd_sc_hd__nor2_4
XFILLER_85_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13198__A _11912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17129_ _17135_/A VGND VGND VPWR VPWR _17130_/A sky130_fd_sc_hd__inv_2
XANTENNA__17893__A _17680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20140_ IRQ[13] VGND VGND VPWR VPWR _20140_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22578__B1 _16266_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20071_ _20071_/A _20071_/B VGND VGND VPWR VPWR _20071_/X sky130_fd_sc_hd__or2_4
XANTENNA__12830__A _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23830_ _23473_/CLK _21415_/X VGND VGND VPWR VPWR _12294_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23761_ _23122_/CLK _23761_/D VGND VGND VPWR VPWR _13145_/B sky130_fd_sc_hd__dfxtp_4
X_20973_ _20759_/X _20972_/X _24288_/Q _20769_/X VGND VGND VPWR VPWR _20974_/B sky130_fd_sc_hd__o22a_4
X_22712_ _21291_/A _22707_/X _14909_/B _22668_/X VGND VGND VPWR VPWR _23072_/D sky130_fd_sc_hd__o22a_4
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13661__A _13641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23692_ _23692_/CLK _23692_/D VGND VGND VPWR VPWR _15504_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22974__A _18375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22643_ _22636_/A VGND VGND VPWR VPWR _22643_/X sky130_fd_sc_hd__buf_2
XFILLER_53_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12277__A _12198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23151__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22574_ _22394_/X _22572_/X _16631_/B _22569_/X VGND VGND VPWR VPWR _23164_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21856__A2 _21853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20494__A _20494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24313_ _24301_/CLK _19150_/X HRESETn VGND VGND VPWR VPWR _19134_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21525_ _21524_/X _21520_/X _12229_/B _21515_/X VGND VGND VPWR VPWR _21525_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24244_ _24032_/CLK _19327_/X HRESETn VGND VGND VPWR VPWR _24244_/Q sky130_fd_sc_hd__dfrtp_4
X_21456_ _21470_/A VGND VGND VPWR VPWR _21456_/X sky130_fd_sc_hd__buf_2
XANTENNA__22805__A1 _17411_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21608__A2 _21605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18899__A _18877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20407_ _20407_/A VGND VGND VPWR VPWR _20407_/X sky130_fd_sc_hd__buf_2
XANTENNA__17288__A2 _17012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24175_ _24180_/CLK _24175_/D HRESETn VGND VGND VPWR VPWR _11737_/A sky130_fd_sc_hd__dfrtp_4
X_21387_ _21373_/A VGND VGND VPWR VPWR _21387_/X sky130_fd_sc_hd__buf_2
XANTENNA__22281__A2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23126_ _23217_/CLK _23126_/D VGND VGND VPWR VPWR _12293_/B sky130_fd_sc_hd__dfxtp_4
X_20338_ _20338_/A VGND VGND VPWR VPWR _21795_/A sky130_fd_sc_hd__buf_2
XFILLER_107_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23057_ _19953_/X _23038_/B VGND VGND VPWR VPWR _23058_/C sky130_fd_sc_hd__or2_4
XFILLER_62_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17308__A _17143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20269_ _20247_/X _20263_/X _20493_/A _20268_/X VGND VGND VPWR VPWR _20269_/X sky130_fd_sc_hd__a211o_4
XFILLER_7_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12740__A _12740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16212__A _16227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22008_ _21850_/X _22002_/X _14497_/B _22006_/X VGND VGND VPWR VPWR _23493_/D sky130_fd_sc_hd__o22a_4
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14830_ _14811_/A _14766_/B VGND VGND VPWR VPWR _14830_/X sky130_fd_sc_hd__or2_4
XANTENNA__23045__A _22898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15770__B _15697_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11973_ _12112_/A _11973_/B _11973_/C VGND VGND VPWR VPWR _11973_/X sky130_fd_sc_hd__or3_4
X_14761_ _11929_/A _14757_/X _14760_/X VGND VGND VPWR VPWR _14761_/X sky130_fd_sc_hd__or3_4
XFILLER_29_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23959_ _24084_/CLK _21178_/X VGND VGND VPWR VPWR _23959_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19365__A2_N _19364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18139__A _18267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16500_ _16158_/A _16437_/B VGND VGND VPWR VPWR _16502_/B sky130_fd_sc_hd__or2_4
X_13712_ _11648_/X _13712_/B VGND VGND VPWR VPWR _13712_/X sky130_fd_sc_hd__or2_4
X_14692_ _14666_/X _14692_/B VGND VGND VPWR VPWR _14692_/X sky130_fd_sc_hd__or2_4
X_17480_ _17477_/Y _17014_/A _17022_/A _17479_/X VGND VGND VPWR VPWR _17480_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22884__A _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16431_ _16146_/A _16508_/B VGND VGND VPWR VPWR _16432_/C sky130_fd_sc_hd__or2_4
XFILLER_108_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13643_ _13643_/A VGND VGND VPWR VPWR _15443_/A sky130_fd_sc_hd__buf_2
XFILLER_73_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19150_ _19134_/A _19151_/A _19149_/Y VGND VGND VPWR VPWR _19150_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13574_ _11657_/X _13574_/B _13574_/C VGND VGND VPWR VPWR _13574_/X sky130_fd_sc_hd__and3_4
X_16362_ _16355_/X _16358_/X _16361_/X VGND VGND VPWR VPWR _16362_/X sky130_fd_sc_hd__or3_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ _18101_/A VGND VGND VPWR VPWR _18242_/A sky130_fd_sc_hd__buf_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _12904_/A _12525_/B VGND VGND VPWR VPWR _12525_/X sky130_fd_sc_hd__or2_4
X_15313_ _13839_/A _15252_/B VGND VGND VPWR VPWR _15315_/B sky130_fd_sc_hd__or2_4
XANTENNA__15498__A _13737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16293_ _11884_/X _16293_/B VGND VGND VPWR VPWR _16293_/X sky130_fd_sc_hd__or2_4
X_19081_ _19074_/X _19080_/X _19074_/X _24325_/Q VGND VGND VPWR VPWR _24325_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12915__A _12915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18032_ _18032_/A VGND VGND VPWR VPWR _18032_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12456_ _12865_/A _12586_/B VGND VGND VPWR VPWR _12457_/C sky130_fd_sc_hd__or2_4
X_15244_ _14210_/A _23617_/Q VGND VGND VPWR VPWR _15245_/C sky130_fd_sc_hd__or2_4
XFILLER_51_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15175_ _14146_/X _15171_/X _15175_/C VGND VGND VPWR VPWR _15175_/X sky130_fd_sc_hd__or3_4
XFILLER_86_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15010__B _23903_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12387_ _12386_/X _12263_/B VGND VGND VPWR VPWR _12388_/C sky130_fd_sc_hd__or2_4
XFILLER_103_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18476__B2 _18475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23794__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14126_ _11608_/A _14124_/X _14125_/X VGND VGND VPWR VPWR _14126_/X sky130_fd_sc_hd__and3_4
XANTENNA__21480__B1 _23788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19983_ _19970_/X _17646_/A _19976_/X _19982_/X VGND VGND VPWR VPWR _19983_/X sky130_fd_sc_hd__o22a_4
XFILLER_113_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22124__A _20778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14057_ _14045_/A _23786_/Q VGND VGND VPWR VPWR _14058_/C sky130_fd_sc_hd__or2_4
X_18934_ _18934_/A VGND VGND VPWR VPWR _18987_/A sky130_fd_sc_hd__inv_2
XFILLER_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13746__A _12646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12650__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16122__A _11982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22206__A2_N _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13008_ _12915_/A _24018_/Q VGND VGND VPWR VPWR _13010_/B sky130_fd_sc_hd__or2_4
X_18865_ _12036_/X _12096_/A VGND VGND VPWR VPWR _18866_/D sky130_fd_sc_hd__or2_4
XFILLER_80_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22778__B _18752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17816_ _17814_/X _17158_/X _17815_/X _17180_/X VGND VGND VPWR VPWR _17816_/X sky130_fd_sc_hd__o22a_4
XFILLER_62_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19433__A _19433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18796_ _18789_/A VGND VGND VPWR VPWR _18796_/X sky130_fd_sc_hd__buf_2
X_17747_ _17716_/X _17747_/B _17746_/X VGND VGND VPWR VPWR _17747_/X sky130_fd_sc_hd__or3_4
X_14959_ _14937_/A _14892_/B VGND VGND VPWR VPWR _14959_/X sky130_fd_sc_hd__or2_4
XANTENNA__21535__A1 _21534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23174__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13481__A _13477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21535__B2 _21527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22732__B1 SYSTICKCLKDIV[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17678_ _17674_/A _17506_/X _17675_/B VGND VGND VPWR VPWR _17678_/X sky130_fd_sc_hd__a21bo_4
XFILLER_62_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12809__B _23956_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19417_ _19449_/A VGND VGND VPWR VPWR _19490_/A sky130_fd_sc_hd__inv_2
XFILLER_51_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12028__A1 _11992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16629_ _11754_/X VGND VGND VPWR VPWR _16629_/X sky130_fd_sc_hd__buf_2
XANTENNA__17888__A _18129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_2_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19348_ _19347_/X _18576_/X _19347_/X _20833_/A VGND VGND VPWR VPWR _19348_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_82_0_HCLK clkbuf_7_82_0_HCLK/A VGND VGND VPWR VPWR _24365_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18703__A2 _18700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19279_ _19214_/B VGND VGND VPWR VPWR _19279_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12825__A _12813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21310_ _21229_/X _21305_/X _16413_/B _21309_/X VGND VGND VPWR VPWR _21310_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15201__A _15201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22290_ _22269_/A VGND VGND VPWR VPWR _22290_/X sky130_fd_sc_hd__buf_2
XFILLER_50_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21241_ _20487_/A VGND VGND VPWR VPWR _21241_/X sky130_fd_sc_hd__buf_2
XFILLER_89_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19608__A _19481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18512__A _18381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20761__B _20595_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21172_ _20356_/X _21169_/X _23963_/Q _21166_/X VGND VGND VPWR VPWR _23963_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15855__B _15855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20123_ _20122_/X VGND VGND VPWR VPWR _20123_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18219__A1 _18216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13656__A _13630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22015__A2 _21988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12560__A _11670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22969__A _18407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21873__A _21887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20054_ _18511_/X _20033_/X _20053_/Y _20044_/X VGND VGND VPWR VPWR _20054_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21774__B2 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15871__A _13554_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19343__A _19336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16686__B _16749_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23813_ _23973_/CLK _21439_/X VGND VGND VPWR VPWR _14470_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14487__A _13623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11904__A _11875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13391__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23744_ _23073_/CLK _23744_/D VGND VGND VPWR VPWR _14864_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ _24193_/Q _20873_/X _20955_/Y VGND VGND VPWR VPWR _22458_/A sky130_fd_sc_hd__o21a_4
XANTENNA__24257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12719__B _23956_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_31_0_HCLK_A clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23707_/CLK _23675_/D VGND VGND VPWR VPWR _23675_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _18641_/Y _20680_/X _20731_/X _20886_/Y VGND VGND VPWR VPWR _20887_/X sky130_fd_sc_hd__a211o_4
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22626_ _22626_/A VGND VGND VPWR VPWR _22626_/X sky130_fd_sc_hd__buf_2
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22557_ _22521_/A VGND VGND VPWR VPWR _22557_/X sky130_fd_sc_hd__buf_2
XANTENNA__12735__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16207__A _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20501__A2 _20499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12310_ _15552_/A VGND VGND VPWR VPWR _12745_/A sky130_fd_sc_hd__buf_2
X_21508_ _21532_/A VGND VGND VPWR VPWR _21508_/X sky130_fd_sc_hd__buf_2
XANTENNA__15111__A _15107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13290_ _12503_/A _13285_/X _13289_/X VGND VGND VPWR VPWR _13290_/X sky130_fd_sc_hd__or3_4
X_22488_ _22418_/X _22486_/X _13045_/B _22483_/X VGND VGND VPWR VPWR _22488_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12241_ _12240_/X _12241_/B VGND VGND VPWR VPWR _12241_/X sky130_fd_sc_hd__or2_4
X_24227_ _24229_/CLK _19352_/X HRESETn VGND VGND VPWR VPWR _24227_/Q sky130_fd_sc_hd__dfrtp_4
X_21439_ _21280_/X _21433_/X _14470_/B _21437_/X VGND VGND VPWR VPWR _21439_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14950__A _15074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18422__A _18244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12172_ _11730_/X _12172_/B _12172_/C VGND VGND VPWR VPWR _12172_/X sky130_fd_sc_hd__and3_4
X_24158_ _24293_/CLK _24158_/D HRESETn VGND VGND VPWR VPWR _24158_/Q sky130_fd_sc_hd__dfrtp_4
X_23109_ _23557_/CLK _22656_/X VGND VGND VPWR VPWR _14539_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13566__A _13554_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16980_ _16948_/Y _16980_/B VGND VGND VPWR VPWR _16981_/B sky130_fd_sc_hd__or2_4
X_24089_ _23514_/CLK _24089_/D VGND VGND VPWR VPWR _16365_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12470__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19958__A1 _19985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15931_ _11872_/X VGND VGND VPWR VPWR _15936_/A sky130_fd_sc_hd__buf_2
XFILLER_88_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15781__A _15778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21765__B2 _21759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18650_ _18381_/A VGND VGND VPWR VPWR _18650_/X sky130_fd_sc_hd__buf_2
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15862_ _13522_/A _15862_/B _15862_/C VGND VGND VPWR VPWR _15862_/X sky130_fd_sc_hd__and3_4
XFILLER_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17601_ _17601_/A _17600_/X VGND VGND VPWR VPWR _17602_/B sky130_fd_sc_hd__and2_4
XFILLER_97_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14813_ _14813_/A _14742_/B VGND VGND VPWR VPWR _14815_/B sky130_fd_sc_hd__or2_4
X_18581_ _17307_/Y _18630_/A _17309_/X VGND VGND VPWR VPWR _18581_/X sky130_fd_sc_hd__o21a_4
X_15793_ _12859_/A _15791_/X _15793_/C VGND VGND VPWR VPWR _15793_/X sky130_fd_sc_hd__and3_4
XFILLER_92_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17532_ _17531_/X VGND VGND VPWR VPWR _17532_/Y sky130_fd_sc_hd__inv_2
X_14744_ _13800_/A _14744_/B _14744_/C VGND VGND VPWR VPWR _14744_/X sky130_fd_sc_hd__and3_4
X_11956_ _15533_/A VGND VGND VPWR VPWR _15707_/A sky130_fd_sc_hd__buf_2
X_17463_ _17156_/Y _17461_/B VGND VGND VPWR VPWR _17464_/B sky130_fd_sc_hd__and2_4
XFILLER_32_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11887_ _11886_/X VGND VGND VPWR VPWR _11888_/A sky130_fd_sc_hd__buf_2
X_14675_ _14210_/A VGND VGND VPWR VPWR _14714_/A sky130_fd_sc_hd__buf_2
X_19202_ _19108_/X VGND VGND VPWR VPWR _19202_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16414_ _16002_/A _23962_/Q VGND VGND VPWR VPWR _16414_/X sky130_fd_sc_hd__or2_4
X_13626_ _13659_/A VGND VGND VPWR VPWR _13794_/A sky130_fd_sc_hd__buf_2
X_17394_ _13685_/Y _17340_/X _17020_/A _17393_/X VGND VGND VPWR VPWR _17395_/B sky130_fd_sc_hd__o22a_4
XFILLER_32_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22119__A _20722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19133_ _24312_/Q _19132_/X VGND VGND VPWR VPWR _19151_/A sky130_fd_sc_hd__and2_4
XANTENNA__21023__A _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16345_ _16447_/A _16345_/B _16345_/C VGND VGND VPWR VPWR _16346_/C sky130_fd_sc_hd__and3_4
X_13557_ _13557_/A _13545_/X _13556_/X VGND VGND VPWR VPWR _13573_/B sky130_fd_sc_hd__and3_4
XANTENNA__12645__A _12964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15021__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12508_ _12472_/A VGND VGND VPWR VPWR _12509_/A sky130_fd_sc_hd__buf_2
X_19064_ _19060_/X _19063_/X _19060_/X _24328_/Q VGND VGND VPWR VPWR _19064_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13488_ _12874_/A _23855_/Q VGND VGND VPWR VPWR _13489_/C sky130_fd_sc_hd__or2_4
X_16276_ _16252_/X _24057_/Q VGND VGND VPWR VPWR _16277_/C sky130_fd_sc_hd__or2_4
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18015_ _24190_/Q VGND VGND VPWR VPWR _18016_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12439_ _12439_/A VGND VGND VPWR VPWR _15392_/A sky130_fd_sc_hd__buf_2
X_15227_ _14183_/A _15227_/B _15226_/X VGND VGND VPWR VPWR _15227_/X sky130_fd_sc_hd__and3_4
XANTENNA__15956__A _15956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22245__A2 _22243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15158_ _14138_/X _23585_/Q VGND VGND VPWR VPWR _15158_/X sky130_fd_sc_hd__or2_4
XFILLER_99_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14109_ _15045_/A VGND VGND VPWR VPWR _14994_/A sky130_fd_sc_hd__buf_2
XANTENNA__13476__A _13448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15089_ _11723_/A _15087_/X _15088_/X VGND VGND VPWR VPWR _15089_/X sky130_fd_sc_hd__and3_4
X_19966_ _24476_/Q VGND VGND VPWR VPWR _19966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22789__A _14493_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21205__B1 _14689_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18917_ _15379_/X _18912_/X _19094_/A _18913_/X VGND VGND VPWR VPWR _24354_/D sky130_fd_sc_hd__o22a_4
XFILLER_84_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16880__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19897_ _23027_/A VGND VGND VPWR VPWR _22932_/A sky130_fd_sc_hd__buf_2
XFILLER_60_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16787__A _11834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21756__A1 _21531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21756__B2 _21752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15691__A _15664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18848_ _18841_/A VGND VGND VPWR VPWR _18848_/X sky130_fd_sc_hd__buf_2
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18779_ _12430_/X _18774_/X _24438_/Q _18775_/X VGND VGND VPWR VPWR _24438_/D sky130_fd_sc_hd__o22a_4
XFILLER_3_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20810_ _20759_/X _20809_/X _24295_/Q _20769_/X VGND VGND VPWR VPWR _20811_/B sky130_fd_sc_hd__o22a_4
XANTENNA__11724__A _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21790_ _21783_/Y _21788_/X _21789_/X _21788_/X VGND VGND VPWR VPWR _21790_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14100__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17188__A1 _13591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22181__B2 _22176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20741_ _20630_/A _20741_/B VGND VGND VPWR VPWR _20741_/Y sky130_fd_sc_hd__nor2_4
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23460_ _23907_/CLK _23460_/D VGND VGND VPWR VPWR _14624_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17411__A _14174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20672_ _20613_/X _20671_/X _15829_/B _20592_/X VGND VGND VPWR VPWR _20672_/X sky130_fd_sc_hd__o22a_4
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22411_ _22423_/A VGND VGND VPWR VPWR _22411_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23391_ _23391_/CLK _23391_/D VGND VGND VPWR VPWR _23391_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22484__A2 _22479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12555__A _13017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22342_ _22079_/X _22340_/X _16620_/B _22337_/X VGND VGND VPWR VPWR _22342_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20194__D _20206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20495__B2 _20449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21692__B1 _23677_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21868__A _21901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15866__A _13507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22273_ _22100_/X _22272_/X _12928_/B _22269_/X VGND VGND VPWR VPWR _23347_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14770__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18242__A _18242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24012_ _23404_/CLK _21092_/X VGND VGND VPWR VPWR _15465_/B sky130_fd_sc_hd__dfxtp_4
X_21224_ _21221_/X _21223_/X _23933_/Q _21218_/X VGND VGND VPWR VPWR _23933_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21444__B1 _23809_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17112__A1 _17109_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17112__B2 _17111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20798__A2 _20797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21155_ _20893_/X _21154_/X _14680_/B _21151_/X VGND VGND VPWR VPWR _23972_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18860__A1 _15379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12290__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20106_ _20074_/Y _20105_/X _11622_/X VGND VGND VPWR VPWR _20106_/X sky130_fd_sc_hd__o21a_4
X_21086_ _21079_/A VGND VGND VPWR VPWR _21086_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21747__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20037_ _20037_/A VGND VGND VPWR VPWR _20037_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11810_ _11803_/A _11810_/B VGND VGND VPWR VPWR _11810_/X sky130_fd_sc_hd__or2_4
XANTENNA__13988__A1 _11976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15106__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21922__A2_N _21921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19801__A _19742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12790_ _13563_/A _12788_/X _12790_/C VGND VGND VPWR VPWR _12798_/B sky130_fd_sc_hd__and3_4
X_21988_ _21988_/A VGND VGND VPWR VPWR _21988_/X sky130_fd_sc_hd__buf_2
XFILLER_2_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14010__A _14010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _12613_/A VGND VGND VPWR VPWR _11741_/X sky130_fd_sc_hd__buf_2
X_20939_ _20844_/A _20939_/B VGND VGND VPWR VPWR _20939_/X sky130_fd_sc_hd__or2_4
X_23727_ _23983_/CLK _23727_/D VGND VGND VPWR VPWR _13504_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_42_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14945__A _11645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _13133_/A VGND VGND VPWR VPWR _12787_/A sky130_fd_sc_hd__buf_2
X_14460_ _12269_/A _14460_/B VGND VGND VPWR VPWR _14460_/X sky130_fd_sc_hd__and2_4
XFILLER_109_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23658_ _23978_/CLK _21718_/X VGND VGND VPWR VPWR _23658_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ _13351_/X _13411_/B _13410_/X VGND VGND VPWR VPWR _13415_/B sky130_fd_sc_hd__and3_4
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _15584_/A _14302_/B VGND VGND VPWR VPWR _14392_/C sky130_fd_sc_hd__or2_4
X_22609_ _22454_/X _22607_/X _23139_/Q _22604_/X VGND VGND VPWR VPWR _23139_/D sky130_fd_sc_hd__o22a_4
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23589_ _23365_/CLK _21851_/X VGND VGND VPWR VPWR _14535_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12465__A _12465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22475__A2 _22472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13342_ _12740_/A _13342_/B _13341_/X VGND VGND VPWR VPWR _13342_/X sky130_fd_sc_hd__and3_4
X_16130_ _16130_/A _16130_/B _16130_/C VGND VGND VPWR VPWR _16130_/X sky130_fd_sc_hd__or3_4
XFILLER_100_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13273_ _13272_/X VGND VGND VPWR VPWR _13273_/Y sky130_fd_sc_hd__inv_2
X_16061_ _16037_/A _23096_/Q VGND VGND VPWR VPWR _16063_/B sky130_fd_sc_hd__or2_4
XANTENNA__15776__A _13133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22227__A2 _22222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12224_ _12691_/A _12224_/B VGND VGND VPWR VPWR _12224_/X sky130_fd_sc_hd__or2_4
X_15012_ _15045_/A _15012_/B _15011_/X VGND VGND VPWR VPWR _15016_/B sky130_fd_sc_hd__and3_4
XFILLER_100_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19820_ _19819_/X VGND VGND VPWR VPWR _19820_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21986__B2 _21985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12155_ _11774_/A _23613_/Q VGND VGND VPWR VPWR _12155_/X sky130_fd_sc_hd__or2_4
XFILLER_69_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18851__A1 _14261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19751_ HRDATA[18] VGND VGND VPWR VPWR _20939_/B sky130_fd_sc_hd__buf_2
X_12086_ _12086_/A _23613_/Q VGND VGND VPWR VPWR _12088_/B sky130_fd_sc_hd__or2_4
X_16963_ _18681_/A VGND VGND VPWR VPWR _17735_/A sky130_fd_sc_hd__inv_2
X_18702_ _18701_/X _18609_/Y _18681_/X VGND VGND VPWR VPWR _18702_/X sky130_fd_sc_hd__a21o_4
X_15914_ _15914_/A _15914_/B _15914_/C _15914_/D VGND VGND VPWR VPWR _15914_/X sky130_fd_sc_hd__or4_4
X_19682_ _20445_/B _19551_/X _19681_/X _19616_/X VGND VGND VPWR VPWR _19682_/X sky130_fd_sc_hd__a211o_4
XFILLER_65_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16894_ _16894_/A VGND VGND VPWR VPWR _16916_/B sky130_fd_sc_hd__buf_2
XFILLER_76_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18633_ _17306_/X _18633_/B VGND VGND VPWR VPWR _18633_/X sky130_fd_sc_hd__or2_4
X_15845_ _12384_/X _15845_/B VGND VGND VPWR VPWR _15847_/B sky130_fd_sc_hd__or2_4
XFILLER_94_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24108__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18564_ _18082_/A _18146_/X VGND VGND VPWR VPWR _18564_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19711__A HRDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15776_ _13133_/A _15768_/X _15775_/X VGND VGND VPWR VPWR _15776_/X sky130_fd_sc_hd__and3_4
XFILLER_40_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12988_ _12392_/A _12988_/B _12988_/C VGND VGND VPWR VPWR _12988_/X sky130_fd_sc_hd__or3_4
XANTENNA__14640__A2 _13595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17515_ _17498_/X VGND VGND VPWR VPWR _17515_/Y sky130_fd_sc_hd__inv_2
X_14727_ _14727_/A _14725_/X _14727_/C VGND VGND VPWR VPWR _14727_/X sky130_fd_sc_hd__and3_4
XFILLER_55_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11939_ _11921_/X _21498_/A VGND VGND VPWR VPWR _11940_/C sky130_fd_sc_hd__or2_4
X_18495_ _17422_/C _18493_/X VGND VGND VPWR VPWR _18495_/X sky130_fd_sc_hd__or2_4
XANTENNA__18327__A _18327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21910__B2 _21905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20576__B _20576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17446_ _12992_/X _17524_/B VGND VGND VPWR VPWR _17446_/X sky130_fd_sc_hd__and2_4
X_14658_ _14658_/A VGND VGND VPWR VPWR _15115_/A sky130_fd_sc_hd__buf_2
XFILLER_21_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13609_ _15404_/A _13607_/X _13608_/X VGND VGND VPWR VPWR _13609_/X sky130_fd_sc_hd__and3_4
X_17377_ _15909_/B _17377_/B VGND VGND VPWR VPWR _17377_/X sky130_fd_sc_hd__or2_4
XFILLER_18_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14589_ _14588_/X VGND VGND VPWR VPWR _14725_/A sky130_fd_sc_hd__buf_2
X_19116_ _24295_/Q _19116_/B VGND VGND VPWR VPWR _19117_/B sky130_fd_sc_hd__and2_4
XANTENNA__20477__A1 _20293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16328_ _16365_/A _16267_/B VGND VGND VPWR VPWR _16329_/C sky130_fd_sc_hd__or2_4
XFILLER_118_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21688__A _21687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21674__B1 _14330_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20592__A _20488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12094__B _23421_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19047_ _19030_/X _19045_/X _19046_/X _24331_/Q VGND VGND VPWR VPWR _24331_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15686__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16259_ _16286_/A _16259_/B VGND VGND VPWR VPWR _16259_/X sky130_fd_sc_hd__or2_4
XANTENNA__22218__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19619__B1 HRDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18062__A _18062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14590__A _14725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19095__A1 _18965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21977__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11719__A _11692_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19949_ _17049_/B _19948_/Y VGND VGND VPWR VPWR _19949_/X sky130_fd_sc_hd__or2_4
XFILLER_101_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21729__B2 _21723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13934__A _15036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22960_ _22955_/X _18344_/X _22937_/X _22959_/X VGND VGND VPWR VPWR _22961_/A sky130_fd_sc_hd__a211o_4
XFILLER_68_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17406__A _17171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21911_ _21857_/X _21908_/X _15274_/B _21905_/X VGND VGND VPWR VPWR _23554_/D sky130_fd_sc_hd__o22a_4
XFILLER_83_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22891_ _23015_/A VGND VGND VPWR VPWR _23048_/A sky130_fd_sc_hd__buf_2
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21842_ _21840_/X _21841_/X _23593_/Q _21836_/X VGND VGND VPWR VPWR _21842_/X sky130_fd_sc_hd__o22a_4
XFILLER_58_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19555__C1 _19554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21773_ _21752_/A VGND VGND VPWR VPWR _21773_/X sky130_fd_sc_hd__buf_2
XFILLER_110_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24333__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20724_ _20488_/A VGND VGND VPWR VPWR _20724_/X sky130_fd_sc_hd__buf_2
X_23512_ _23539_/CLK _23512_/D VGND VGND VPWR VPWR _23512_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23443_ _23827_/CLK _22102_/X VGND VGND VPWR VPWR _23443_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20655_ _24397_/Q _20595_/B VGND VGND VPWR VPWR _20655_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22457__A2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12285__A _12284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19858__B1 _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_52_0_HCLK clkbuf_6_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23374_ _23342_/CLK _22230_/X VGND VGND VPWR VPWR _15757_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21598__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20586_ _24240_/Q VGND VGND VPWR VPWR _20586_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17333__A1 _15251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22325_ _22325_/A VGND VGND VPWR VPWR _23301_/D sky130_fd_sc_hd__buf_2
XFILLER_118_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22256_ _22250_/Y _22255_/X _22073_/X _22255_/X VGND VGND VPWR VPWR _22256_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21207_ _20937_/X _21204_/X _15283_/B _21201_/X VGND VGND VPWR VPWR _23938_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18833__A1 _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22090__B1 _15969_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22187_ _22124_/X _22186_/X _23401_/Q _22183_/X VGND VGND VPWR VPWR _23401_/D sky130_fd_sc_hd__o22a_4
X_21138_ _20591_/X _21133_/X _23984_/Q _21137_/X VGND VGND VPWR VPWR _23984_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22222__A _22222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19515__B _19481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_HCLK_A clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13960_ _13960_/A _23946_/Q VGND VGND VPWR VPWR _13961_/C sky130_fd_sc_hd__or2_4
X_21069_ _20315_/X _21068_/X _24029_/Q _21065_/X VGND VGND VPWR VPWR _24029_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16220__A _16227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21196__A2 _21190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22393__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12911_ _12497_/X _12983_/B VGND VGND VPWR VPWR _12911_/X sky130_fd_sc_hd__or2_4
X_13891_ _13879_/A _24039_/Q VGND VGND VPWR VPWR _13892_/C sky130_fd_sc_hd__or2_4
XANTENNA__24201__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15630_ _15618_/A _23787_/Q VGND VGND VPWR VPWR _15630_/X sky130_fd_sc_hd__or2_4
X_12842_ _12752_/Y _12841_/X VGND VGND VPWR VPWR _12842_/X sky130_fd_sc_hd__and2_4
XFILLER_74_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20677__A _20317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23235__CLK _23107_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23053__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15561_ _15534_/A _15559_/X _15560_/X VGND VGND VPWR VPWR _15561_/X sky130_fd_sc_hd__and3_4
X_12773_ _12808_/A _12773_/B VGND VGND VPWR VPWR _12775_/B sky130_fd_sc_hd__or2_4
XFILLER_64_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22696__A2 _22693_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18147__A _18392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14675__A _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17299_/Y _17286_/A VGND VGND VPWR VPWR _17300_/X sky130_fd_sc_hd__or2_4
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14494_/X _14509_/X _14512_/C VGND VGND VPWR VPWR _14512_/X sky130_fd_sc_hd__and3_4
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11724_ _12412_/A VGND VGND VPWR VPWR _13214_/A sky130_fd_sc_hd__buf_2
X_18280_ _18216_/X _17508_/X _18276_/X _18082_/X _18279_/Y VGND VGND VPWR VPWR _18280_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_14_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _13731_/A _15488_/X _15492_/C VGND VGND VPWR VPWR _15492_/X sky130_fd_sc_hd__or3_4
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17165_/Y _17137_/X _14565_/Y _17138_/X VGND VGND VPWR VPWR _17231_/X sky130_fd_sc_hd__o22a_4
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _13918_/A VGND VGND VPWR VPWR _11656_/A sky130_fd_sc_hd__buf_2
X_14443_ _12885_/A _14511_/B VGND VGND VPWR VPWR _14444_/C sky130_fd_sc_hd__or2_4
XFILLER_35_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19849__B1 _21007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22448__A2 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16890__A _16821_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17162_ _14723_/B _17161_/X _16376_/X _17157_/X VGND VGND VPWR VPWR _17162_/X sky130_fd_sc_hd__o22a_4
XFILLER_70_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11586_ _11633_/A VGND VGND VPWR VPWR _17024_/B sky130_fd_sc_hd__inv_2
X_14374_ _13844_/A VGND VGND VPWR VPWR _15637_/A sky130_fd_sc_hd__buf_2
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16113_ _16113_/A _16113_/B _16113_/C VGND VGND VPWR VPWR _16113_/X sky130_fd_sc_hd__or3_4
XANTENNA__21301__A _21316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13325_ _13286_/X _13325_/B VGND VGND VPWR VPWR _13325_/X sky130_fd_sc_hd__or2_4
X_17093_ _18656_/A VGND VGND VPWR VPWR _18103_/A sky130_fd_sc_hd__inv_2
XANTENNA__21408__B1 _23835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16044_ _16215_/A _16044_/B _16044_/C VGND VGND VPWR VPWR _16044_/X sky130_fd_sc_hd__and3_4
X_13256_ _13256_/A _13196_/B VGND VGND VPWR VPWR _13256_/X sky130_fd_sc_hd__or2_4
XFILLER_83_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12207_ _12880_/A VGND VGND VPWR VPWR _13984_/A sky130_fd_sc_hd__buf_2
X_13187_ _12737_/A _13185_/X _13187_/C VGND VGND VPWR VPWR _13187_/X sky130_fd_sc_hd__and3_4
XANTENNA__18824__A1 _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19706__A _19706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20631__A1 _18407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12138_ _11773_/X _12136_/X _12138_/C VGND VGND VPWR VPWR _12138_/X sky130_fd_sc_hd__and3_4
X_19803_ _19876_/B _19718_/B VGND VGND VPWR VPWR _19803_/X sky130_fd_sc_hd__or2_4
XFILLER_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17995_ _17989_/X _17547_/X _17991_/X _17874_/X _17994_/Y VGND VGND VPWR VPWR _17995_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22132__A _22108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13754__A _13754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12069_ _12093_/A _12146_/B VGND VGND VPWR VPWR _12069_/X sky130_fd_sc_hd__or2_4
X_16946_ _24130_/Q VGND VGND VPWR VPWR _16946_/Y sky130_fd_sc_hd__inv_2
X_19734_ HRDATA[4] VGND VGND VPWR VPWR _19734_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21971__A _21970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19665_ _19800_/B _19793_/B _19672_/D _19500_/X VGND VGND VPWR VPWR _19665_/X sky130_fd_sc_hd__and4_4
XFILLER_93_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16877_ _16519_/A _16829_/X _16519_/A _16829_/X VGND VGND VPWR VPWR _16879_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15391__D _16840_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18616_ _18614_/Y _18615_/X VGND VGND VPWR VPWR _18616_/X sky130_fd_sc_hd__or2_4
XFILLER_53_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15828_ _12904_/A _15828_/B VGND VGND VPWR VPWR _15828_/X sky130_fd_sc_hd__or2_4
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19596_ _19424_/A _19595_/X HRDATA[3] _19439_/X VGND VGND VPWR VPWR _19597_/A sky130_fd_sc_hd__o22a_4
XFILLER_92_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18547_ _18547_/A VGND VGND VPWR VPWR _18547_/Y sky130_fd_sc_hd__inv_2
X_15759_ _12765_/X _15759_/B _15758_/X VGND VGND VPWR VPWR _15759_/X sky130_fd_sc_hd__and3_4
XANTENNA__22687__A2 _22686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14585__A _14152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20698__A1 _20613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20698__B2 _20592_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21895__B1 _15674_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18478_ _18340_/X _18476_/X _18377_/X _18477_/X VGND VGND VPWR VPWR _18478_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17563__A1 _17560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17563__B2 _17653_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17429_ _17172_/Y _17407_/B _17422_/C _17428_/X VGND VGND VPWR VPWR _17429_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19304__A2 _17044_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20440_ _24215_/Q _20398_/X _20439_/X VGND VGND VPWR VPWR _20441_/A sky130_fd_sc_hd__o21a_4
XFILLER_53_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23878__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14129__A1 _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20371_ _24218_/Q _20282_/X _20370_/Y VGND VGND VPWR VPWR _20372_/A sky130_fd_sc_hd__o21a_4
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12833__A _12803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16305__A _16188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22110_ _20610_/A VGND VGND VPWR VPWR _22110_/X sky130_fd_sc_hd__buf_2
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23090_ _23794_/CLK _22688_/X VGND VGND VPWR VPWR _13119_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_66_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22041_ _21821_/X _22038_/X _23473_/Q _22035_/X VGND VGND VPWR VPWR _22041_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23108__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22611__A2 _22607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15863__B _15863_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22042__A _22035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13664__A _15432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23992_ _24084_/CLK _21127_/X VGND VGND VPWR VPWR _23992_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22943_ _22943_/A VGND VGND VPWR VPWR HADDR[10] sky130_fd_sc_hd__inv_2
XFILLER_25_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22874_ _16596_/Y _22863_/X _19887_/X _22873_/X VGND VGND VPWR VPWR _22875_/B sky130_fd_sc_hd__o22a_4
XANTENNA__20497__A _20497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16694__B _16759_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21825_ _21823_/X _21817_/X _23600_/Q _21824_/X VGND VGND VPWR VPWR _21825_/X sky130_fd_sc_hd__o22a_4
XFILLER_93_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14495__A _12383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22678__A2 _22672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11912__A _11912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21756_ _21531_/X _21755_/X _12912_/B _21752_/X VGND VGND VPWR VPWR _21756_/X sky130_fd_sc_hd__o22a_4
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21886__B1 _23572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17554__B2 _17652_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20707_ _20471_/A VGND VGND VPWR VPWR _20708_/B sky130_fd_sc_hd__buf_2
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15103__B _23775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21687_ _21702_/A VGND VGND VPWR VPWR _21687_/X sky130_fd_sc_hd__buf_2
X_24475_ _24473_/CLK _24475_/D HRESETn VGND VGND VPWR VPWR _19971_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20638_ _20613_/X _20637_/X _15697_/B _20592_/X VGND VGND VPWR VPWR _24078_/D sky130_fd_sc_hd__o22a_4
X_23426_ _23522_/CLK _23426_/D VGND VGND VPWR VPWR _15277_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21102__A2 _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14942__B _14883_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23357_ _23100_/CLK _23357_/D VGND VGND VPWR VPWR _12123_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13839__A _13839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20569_ _20376_/X _20555_/X _20515_/X _20568_/Y VGND VGND VPWR VPWR _20569_/X sky130_fd_sc_hd__a211o_4
XANTENNA__20310__B1 _20288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12743__A _12743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16215__A _16215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13110_ _13082_/A _13110_/B _13110_/C VGND VGND VPWR VPWR _13110_/X sky130_fd_sc_hd__or3_4
X_22308_ _12259_/B VGND VGND VPWR VPWR _22308_/X sky130_fd_sc_hd__buf_2
X_14090_ _12252_/A _14088_/X _14090_/C VGND VGND VPWR VPWR _14099_/B sky130_fd_sc_hd__and3_4
X_23288_ _23383_/CLK _23288_/D VGND VGND VPWR VPWR _15952_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13041_ _13041_/A _13041_/B _13041_/C VGND VGND VPWR VPWR _13041_/X sky130_fd_sc_hd__or3_4
X_22239_ _22129_/X _22236_/X _23367_/Q _22233_/X VGND VGND VPWR VPWR _22239_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18806__A1 _14851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22063__B1 _15240_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22602__A2 _22600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19526__A _19672_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_59_0_HCLK clkbuf_7_58_0_HCLK/A VGND VGND VPWR VPWR _23698_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23048__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21810__B1 _12289_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15773__B _15700_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16800_ _16800_/A _23867_/Q VGND VGND VPWR VPWR _16800_/X sky130_fd_sc_hd__or2_4
XANTENNA__17046__A _17007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13574__A _11657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17780_ _17900_/A VGND VGND VPWR VPWR _18205_/A sky130_fd_sc_hd__buf_2
X_14992_ _14992_/A _15056_/B VGND VGND VPWR VPWR _14994_/B sky130_fd_sc_hd__or2_4
XFILLER_59_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22887__A _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22366__B2 _22365_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16731_ _12065_/X _23643_/Q VGND VGND VPWR VPWR _16732_/C sky130_fd_sc_hd__or2_4
XFILLER_87_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21791__A _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13943_ _12472_/X _23978_/Q VGND VGND VPWR VPWR _13943_/X sky130_fd_sc_hd__or2_4
XANTENNA__24183__CLK _24187_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19450_ _19450_/A VGND VGND VPWR VPWR _19454_/A sky130_fd_sc_hd__buf_2
X_16662_ _16662_/A _23100_/Q VGND VGND VPWR VPWR _16662_/X sky130_fd_sc_hd__or2_4
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13874_ _13862_/A VGND VGND VPWR VPWR _13910_/A sky130_fd_sc_hd__buf_2
XFILLER_35_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22118__A1 _22117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18401_ _17382_/A _18400_/X _17431_/Y VGND VGND VPWR VPWR _18401_/X sky130_fd_sc_hd__o21a_4
XFILLER_62_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22118__B2 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15613_ _13886_/A _15613_/B _15613_/C VGND VGND VPWR VPWR _15645_/B sky130_fd_sc_hd__or3_4
X_12825_ _12813_/A _12825_/B _12824_/X VGND VGND VPWR VPWR _12831_/B sky130_fd_sc_hd__and3_4
X_19381_ _19377_/X _19378_/Y _19380_/X _24213_/Q VGND VGND VPWR VPWR _19381_/X sky130_fd_sc_hd__o22a_4
X_16593_ _11853_/X _16592_/X VGND VGND VPWR VPWR _16593_/X sky130_fd_sc_hd__and2_4
XFILLER_62_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12918__A _13015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18332_ _18332_/A _18331_/X VGND VGND VPWR VPWR _18332_/X sky130_fd_sc_hd__or2_4
XANTENNA__11822__A _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15544_ _11955_/A _23563_/Q VGND VGND VPWR VPWR _15545_/C sky130_fd_sc_hd__or2_4
X_12756_ _13088_/A VGND VGND VPWR VPWR _13129_/A sky130_fd_sc_hd__buf_2
XFILLER_61_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21341__A2 _21340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11707_/A VGND VGND VPWR VPWR _11708_/A sky130_fd_sc_hd__buf_2
X_18263_ _18204_/A _17502_/X VGND VGND VPWR VPWR _18263_/X sky130_fd_sc_hd__or2_4
XANTENNA__11541__B IRQ[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _13087_/A _15473_/X _15474_/X VGND VGND VPWR VPWR _15475_/X sky130_fd_sc_hd__and3_4
X_12687_ _12286_/X _12768_/B VGND VGND VPWR VPWR _12687_/X sky130_fd_sc_hd__or2_4
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20854__B _20556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _17152_/X _17212_/X _17163_/X _17213_/X VGND VGND VPWR VPWR _17214_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21629__B1 _15256_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14426_ _14336_/X _14428_/A VGND VGND VPWR VPWR _15389_/A sky130_fd_sc_hd__or2_4
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11638_ _11638_/A VGND VGND VPWR VPWR _13686_/A sky130_fd_sc_hd__buf_2
X_18194_ _18171_/X _19378_/A _18022_/X _18193_/X VGND VGND VPWR VPWR _18194_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22127__A _22127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17145_ _17145_/A VGND VGND VPWR VPWR _17145_/X sky130_fd_sc_hd__buf_2
XANTENNA__13749__A _13697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14357_ _15592_/A _14355_/X _14356_/X VGND VGND VPWR VPWR _14357_/X sky130_fd_sc_hd__and3_4
XFILLER_89_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11569_ _24446_/Q IRQ[31] VGND VGND VPWR VPWR _11569_/X sky130_fd_sc_hd__and2_4
X_13308_ _15685_/A _13308_/B VGND VGND VPWR VPWR _13308_/X sky130_fd_sc_hd__or2_4
XFILLER_116_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17076_ _18418_/A VGND VGND VPWR VPWR _18203_/A sky130_fd_sc_hd__buf_2
X_14288_ _11955_/A VGND VGND VPWR VPWR _15556_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16027_ _16063_/A _16027_/B _16026_/X VGND VGND VPWR VPWR _16028_/C sky130_fd_sc_hd__and3_4
XFILLER_115_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15964__A _11884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13239_ _13239_/A _23953_/Q VGND VGND VPWR VPWR _13240_/C sky130_fd_sc_hd__or2_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18340__A _18198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20604__A1 _18375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21801__B1 _23610_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15683__B _15748_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24123__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13484__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17978_ _17978_/A VGND VGND VPWR VPWR _17978_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22357__B2 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16929_ _17009_/A _16929_/B _11634_/A _17079_/A VGND VGND VPWR VPWR _16929_/X sky130_fd_sc_hd__or4_4
X_19717_ _19710_/X _19713_/X _19716_/X _12100_/X _19697_/X VGND VGND VPWR VPWR _19717_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_66_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16795__A _16624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20907__A2 _20906_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19648_ _19537_/A _19647_/X VGND VGND VPWR VPWR _19648_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22109__B2 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19579_ _19579_/A _19562_/X _19575_/X _19578_/X VGND VGND VPWR VPWR _19579_/X sky130_fd_sc_hd__or4_4
XFILLER_94_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12828__A _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21610_ _21538_/X _21605_/X _23728_/Q _21609_/X VGND VGND VPWR VPWR _21610_/X sky130_fd_sc_hd__o22a_4
X_22590_ _22583_/A VGND VGND VPWR VPWR _22590_/X sky130_fd_sc_hd__buf_2
XANTENNA__17536__A1 _16444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17536__B2 _17535_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21332__A2 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16019__B _16019_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21541_ _21256_/A VGND VGND VPWR VPWR _21541_/X sky130_fd_sc_hd__buf_2
XANTENNA__20540__B1 _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24260_ _24305_/CLK _24260_/D HRESETn VGND VGND VPWR VPWR _19209_/A sky130_fd_sc_hd__dfrtp_4
X_21472_ _21249_/X _21470_/X _13120_/B _21467_/X VGND VGND VPWR VPWR _21472_/X sky130_fd_sc_hd__o22a_4
XFILLER_18_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23211_ _23336_/CLK _22498_/X VGND VGND VPWR VPWR _23211_/Q sky130_fd_sc_hd__dfxtp_4
X_20423_ _20422_/X _20800_/A _20286_/X VGND VGND VPWR VPWR _20423_/X sky130_fd_sc_hd__a21o_4
XANTENNA__13659__A _13659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24191_ _24229_/CLK _24191_/D HRESETn VGND VGND VPWR VPWR _24191_/Q sky130_fd_sc_hd__dfrtp_4
X_23142_ _23781_/CLK _23142_/D VGND VGND VPWR VPWR _14373_/B sky130_fd_sc_hd__dfxtp_4
X_20354_ _24219_/Q _20282_/X _20353_/Y VGND VGND VPWR VPWR _20355_/A sky130_fd_sc_hd__o21a_4
XFILLER_49_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23073_ _23073_/CLK _23073_/D VGND VGND VPWR VPWR _15176_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_66_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15874__A _13557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20285_ _18757_/X VGND VGND VPWR VPWR _20285_/X sky130_fd_sc_hd__buf_2
X_22024_ _22031_/A VGND VGND VPWR VPWR _22024_/X sky130_fd_sc_hd__buf_2
XANTENNA__22596__B2 _22590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15593__B _24011_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19461__A1 _24154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23975_ _24008_/CLK _23975_/D VGND VGND VPWR VPWR _13792_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22500__A _22471_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20939__B _20939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19764__A2 _19789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22926_ _22968_/A VGND VGND VPWR VPWR _22998_/A sky130_fd_sc_hd__buf_2
XFILLER_57_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21571__A2 _21568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21116__A _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22857_ _17560_/Y _22814_/X _22853_/X _22856_/X VGND VGND VPWR VPWR _22858_/B sky130_fd_sc_hd__o22a_4
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20020__A _19996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12738__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12610_ _13083_/A _12588_/X _12609_/X VGND VGND VPWR VPWR _12610_/X sky130_fd_sc_hd__and3_4
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15114__A _15114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21808_ _21807_/X _21805_/X _23607_/Q _21800_/X VGND VGND VPWR VPWR _21808_/X sky130_fd_sc_hd__o22a_4
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ _13426_/X _13590_/B VGND VGND VPWR VPWR _13590_/X sky130_fd_sc_hd__or2_4
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22788_ _17298_/Y _22781_/X VGND VGND VPWR VPWR HWDATA[5] sky130_fd_sc_hd__nor2_4
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22520__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12541_ _12876_/A _12541_/B _12541_/C VGND VGND VPWR VPWR _12541_/X sky130_fd_sc_hd__or3_4
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21739_ _21733_/Y _21738_/X _21504_/X _21738_/X VGND VGND VPWR VPWR _21739_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14953__A _14243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18425__A _18425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15260_ _14318_/A _15260_/B VGND VGND VPWR VPWR _15260_/X sky130_fd_sc_hd__or2_4
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12472_ _12472_/A VGND VGND VPWR VPWR _12472_/X sky130_fd_sc_hd__buf_2
X_24458_ _24202_/CLK _24458_/D HRESETn VGND VGND VPWR VPWR _20053_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14211_ _14371_/A _14208_/X _14210_/X VGND VGND VPWR VPWR _14211_/X sky130_fd_sc_hd__and3_4
X_23409_ _23313_/CLK _23409_/D VGND VGND VPWR VPWR _13249_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21087__B2 _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22284__B1 _23339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_22_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15191_ _15203_/A _15189_/X _15191_/C VGND VGND VPWR VPWR _15192_/C sky130_fd_sc_hd__and3_4
X_24389_ _24425_/CLK _24389_/D HRESETn VGND VGND VPWR VPWR _20854_/A sky130_fd_sc_hd__dfrtp_4
X_14142_ _14113_/A _23369_/Q VGND VGND VPWR VPWR _14144_/B sky130_fd_sc_hd__or2_4
XFILLER_10_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15784__A _15784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14073_ _14073_/A _14039_/X _14073_/C VGND VGND VPWR VPWR _14073_/X sky130_fd_sc_hd__and3_4
X_18950_ _24379_/Q VGND VGND VPWR VPWR _18950_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22587__B2 _22583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13024_ _12465_/A _13024_/B _13024_/C VGND VGND VPWR VPWR _13024_/X sky130_fd_sc_hd__and3_4
X_17901_ _18264_/A _17278_/B VGND VGND VPWR VPWR _17904_/B sky130_fd_sc_hd__and2_4
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18881_ _17266_/X _18875_/X _24380_/Q _18878_/X VGND VGND VPWR VPWR _18881_/X sky130_fd_sc_hd__o22a_4
XFILLER_49_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17832_ _17911_/A _17830_/X _17806_/X _17831_/X VGND VGND VPWR VPWR _17832_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__11817__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17763_ _17659_/X _17660_/X _17651_/X _17762_/X VGND VGND VPWR VPWR _17764_/A sky130_fd_sc_hd__or4_4
XANTENNA__11536__B IRQ[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14975_ _14195_/A _14975_/B _14975_/C VGND VGND VPWR VPWR _14976_/C sky130_fd_sc_hd__and3_4
XANTENNA__22410__A _20486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16714_ _16714_/A _23963_/Q VGND VGND VPWR VPWR _16715_/C sky130_fd_sc_hd__or2_4
X_19502_ _19572_/C VGND VGND VPWR VPWR _19599_/B sky130_fd_sc_hd__buf_2
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13926_ _13951_/A VGND VGND VPWR VPWR _13927_/A sky130_fd_sc_hd__buf_2
XANTENNA__17504__A _13202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17694_ _17694_/A _17367_/X VGND VGND VPWR VPWR _17696_/A sky130_fd_sc_hd__and2_4
XFILLER_74_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19433_ _19433_/A VGND VGND VPWR VPWR _19433_/Y sky130_fd_sc_hd__inv_2
X_16645_ _16624_/X _16635_/X _16644_/X VGND VGND VPWR VPWR _16646_/C sky130_fd_sc_hd__and3_4
X_13857_ _13845_/A _23751_/Q VGND VGND VPWR VPWR _13858_/C sky130_fd_sc_hd__or2_4
XFILLER_90_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12648__A _12640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15024__A _15028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12808_ _12808_/A _23892_/Q VGND VGND VPWR VPWR _12810_/B sky130_fd_sc_hd__or2_4
X_19364_ _19361_/X _23056_/B _19306_/Y _19363_/Y VGND VGND VPWR VPWR _19364_/X sky130_fd_sc_hd__o22a_4
XFILLER_90_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16576_ _12011_/A _16576_/B _16575_/X VGND VGND VPWR VPWR _16577_/C sky130_fd_sc_hd__and3_4
XFILLER_95_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13788_ _12475_/A _13863_/B VGND VGND VPWR VPWR _13789_/C sky130_fd_sc_hd__or2_4
XANTENNA__21314__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18315_ _24126_/Q _18231_/Y _16979_/B VGND VGND VPWR VPWR _22979_/B sky130_fd_sc_hd__o21a_4
XANTENNA__22511__B2 _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15527_ _12307_/A _15525_/X _15526_/X VGND VGND VPWR VPWR _15527_/X sky130_fd_sc_hd__and3_4
XFILLER_37_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12739_ _12739_/A _12836_/B VGND VGND VPWR VPWR _12740_/C sky130_fd_sc_hd__or2_4
X_19295_ _19206_/B VGND VGND VPWR VPWR _19295_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15959__A _15959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18246_ _17837_/X _17917_/X _17846_/X _17923_/X VGND VGND VPWR VPWR _18246_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15458_ _15477_/A _15458_/B VGND VGND VPWR VPWR _15458_/X sky130_fd_sc_hd__or2_4
XFILLER_50_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14409_ _15632_/A _14330_/B VGND VGND VPWR VPWR _14411_/B sky130_fd_sc_hd__or2_4
XFILLER_117_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13479__A _13447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21078__B2 _21072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18177_ _18241_/A _17527_/B VGND VGND VPWR VPWR _18180_/B sky130_fd_sc_hd__nor2_4
XFILLER_89_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15389_ _15389_/A _14566_/X VGND VGND VPWR VPWR _15389_/X sky130_fd_sc_hd__and2_4
XANTENNA__12383__A _12383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17128_ _15050_/Y _17010_/A _17018_/A _17127_/Y VGND VGND VPWR VPWR _17135_/A sky130_fd_sc_hd__o22a_4
XANTENNA__24304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15694__A _12705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17059_ _17028_/A _11584_/A _19927_/A VGND VGND VPWR VPWR _17059_/X sky130_fd_sc_hd__a21o_4
X_20070_ _20070_/A VGND VGND VPWR VPWR _20090_/D sky130_fd_sc_hd__inv_2
XANTENNA__20589__B1 _20588_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11727__A _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_42_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR _23591_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21250__B2 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14103__A _14992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13942__A _13966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20972_ _20760_/X _20971_/X _24320_/Q _20767_/X VGND VGND VPWR VPWR _20972_/X sky130_fd_sc_hd__o22a_4
X_23760_ _23983_/CLK _21540_/X VGND VGND VPWR VPWR _23760_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22711_ _21574_/A _22707_/X _15176_/B _22668_/X VGND VGND VPWR VPWR _23073_/D sky130_fd_sc_hd__o22a_4
XFILLER_81_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23691_ _23688_/CLK _23691_/D VGND VGND VPWR VPWR _23691_/Q sky130_fd_sc_hd__dfxtp_4
X_22642_ _22425_/X _22636_/X _13547_/B _22640_/X VGND VGND VPWR VPWR _23119_/D sky130_fd_sc_hd__o22a_4
XFILLER_59_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22502__B2 _22497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22573_ _22390_/X _22572_/X _12139_/B _22569_/X VGND VGND VPWR VPWR _23165_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15869__A _13529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14773__A _13645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24312_ _24301_/CLK _19152_/X HRESETn VGND VGND VPWR VPWR _24312_/Q sky130_fd_sc_hd__dfrtp_4
X_21524_ _20464_/A VGND VGND VPWR VPWR _21524_/X sky130_fd_sc_hd__buf_2
XFILLER_33_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21455_ _21455_/A VGND VGND VPWR VPWR _21470_/A sky130_fd_sc_hd__buf_2
X_24243_ _24241_/CLK _24243_/D HRESETn VGND VGND VPWR VPWR _24243_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21069__B2 _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22266__B1 _23352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12293__A _12725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20406_ _24408_/Q _20405_/X _24440_/Q _20260_/X VGND VGND VPWR VPWR _20406_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12724__C _12723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24174_ _23812_/CLK _19783_/X HRESETn VGND VGND VPWR VPWR _13688_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21386_ _21275_/X _21383_/X _13906_/B _21380_/X VGND VGND VPWR VPWR _21386_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19682__A1 _20445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20337_ _24220_/Q _20282_/X _20336_/Y VGND VGND VPWR VPWR _20338_/A sky130_fd_sc_hd__o21a_4
X_23125_ _23699_/CLK _22634_/X VGND VGND VPWR VPWR _12647_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23596__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23056_ _23051_/A _23056_/B VGND VGND VPWR VPWR _23056_/X sky130_fd_sc_hd__or2_4
XFILLER_89_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20268_ _20268_/A _20494_/A VGND VGND VPWR VPWR _20268_/X sky130_fd_sc_hd__and2_4
XANTENNA__16212__B _16135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22007_ _21847_/X _22002_/X _14269_/B _22006_/X VGND VGND VPWR VPWR _23494_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20199_ _20199_/A _20199_/B VGND VGND VPWR VPWR _20199_/X sky130_fd_sc_hd__or2_4
XANTENNA__14013__A _14815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14948__A _15063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13852__A _13895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14760_ _13603_/A _14758_/X _14760_/C VGND VGND VPWR VPWR _14760_/X sky130_fd_sc_hd__and3_4
XFILLER_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11972_ _11966_/X _11969_/X _11972_/C VGND VGND VPWR VPWR _11973_/C sky130_fd_sc_hd__and3_4
X_23958_ _24084_/CLK _21179_/X VGND VGND VPWR VPWR _12287_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_79_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13711_ _13911_/A VGND VGND VPWR VPWR _13711_/X sky130_fd_sc_hd__buf_2
XFILLER_79_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22909_ _23027_/A _18643_/X VGND VGND VPWR VPWR _22909_/X sky130_fd_sc_hd__and2_4
XFILLER_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14691_ _11697_/A _14691_/B VGND VGND VPWR VPWR _14691_/X sky130_fd_sc_hd__or2_4
X_23889_ _23889_/CLK _23889_/D VGND VGND VPWR VPWR _13171_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12468__A _13019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22884__B _22924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16430_ _16091_/A _16430_/B VGND VGND VPWR VPWR _16432_/B sky130_fd_sc_hd__or2_4
X_13642_ _13632_/A _13640_/X _13642_/C VGND VGND VPWR VPWR _13647_/B sky130_fd_sc_hd__and3_4
XANTENNA__24221__CLK _24187_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16361_ _11727_/X _16361_/B _16361_/C VGND VGND VPWR VPWR _16361_/X sky130_fd_sc_hd__and3_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15779__A _15778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13573_ _11800_/X _13573_/B _13573_/C VGND VGND VPWR VPWR _13574_/C sky130_fd_sc_hd__or3_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18100_ _18241_/A _17564_/B VGND VGND VPWR VPWR _18100_/Y sky130_fd_sc_hd__nor2_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ _11841_/A _13595_/A _15281_/X _11594_/A _15311_/X VGND VGND VPWR VPWR _15312_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _12915_/A VGND VGND VPWR VPWR _12904_/A sky130_fd_sc_hd__buf_2
X_19080_ _19052_/X _19078_/X _19079_/Y _19057_/X VGND VGND VPWR VPWR _19080_/X sky130_fd_sc_hd__o22a_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _15980_/A _16292_/B _16291_/X VGND VGND VPWR VPWR _16292_/X sky130_fd_sc_hd__or3_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23049__A2 _17769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18031_ _18180_/A _18027_/Y _18031_/C _18030_/X VGND VGND VPWR VPWR _18032_/A sky130_fd_sc_hd__or4_4
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15243_ _14247_/A _15243_/B VGND VGND VPWR VPWR _15245_/B sky130_fd_sc_hd__or2_4
XANTENNA__13299__A _15696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12455_ _12852_/A VGND VGND VPWR VPWR _12865_/A sky130_fd_sc_hd__buf_2
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15174_ _14737_/A _15172_/X _15173_/X VGND VGND VPWR VPWR _15175_/C sky130_fd_sc_hd__and3_4
X_12386_ _12926_/A VGND VGND VPWR VPWR _12386_/X sky130_fd_sc_hd__buf_2
X_14125_ _14997_/A _23433_/Q VGND VGND VPWR VPWR _14125_/X sky130_fd_sc_hd__or2_4
XFILLER_119_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21480__B2 _21474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19982_ _18055_/X _19961_/X _19981_/Y _19972_/X VGND VGND VPWR VPWR _19982_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12931__A _12655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14056_ _14031_/A _23082_/Q VGND VGND VPWR VPWR _14056_/X sky130_fd_sc_hd__or2_4
X_18933_ _18932_/X VGND VGND VPWR VPWR _24349_/D sky130_fd_sc_hd__inv_2
X_13007_ _12887_/A _13005_/X _13006_/X VGND VGND VPWR VPWR _13007_/X sky130_fd_sc_hd__and3_4
XANTENNA__15019__A _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_29_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_58_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18864_ _17262_/A _17273_/A _18864_/C _17413_/A VGND VGND VPWR VPWR _20248_/A sky130_fd_sc_hd__or4_4
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17815_ _17815_/A VGND VGND VPWR VPWR _17815_/X sky130_fd_sc_hd__buf_2
X_18795_ _18788_/A VGND VGND VPWR VPWR _18795_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17746_ _17718_/X _17721_/X _17745_/X VGND VGND VPWR VPWR _17746_/X sky130_fd_sc_hd__and3_4
X_14958_ _14970_/A _23584_/Q VGND VGND VPWR VPWR _14960_/B sky130_fd_sc_hd__or2_4
XFILLER_63_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17739__B2 _17122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21535__A2 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13909_ _13909_/A _23463_/Q VGND VGND VPWR VPWR _13911_/B sky130_fd_sc_hd__or2_4
X_17677_ _17677_/A _17676_/Y VGND VGND VPWR VPWR _17677_/X sky130_fd_sc_hd__or2_4
X_14889_ _13984_/A _14889_/B VGND VGND VPWR VPWR _14889_/X sky130_fd_sc_hd__or2_4
XANTENNA__12378__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16628_ _11782_/A VGND VGND VPWR VPWR _16652_/A sky130_fd_sc_hd__buf_2
X_19416_ _22978_/A _19416_/B VGND VGND VPWR VPWR _19449_/A sky130_fd_sc_hd__or2_4
XFILLER_62_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16792__B _16792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15689__A _15689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16559_ _12024_/A _16559_/B VGND VGND VPWR VPWR _16560_/C sky130_fd_sc_hd__or2_4
X_19347_ _19336_/A VGND VGND VPWR VPWR _19347_/X sky130_fd_sc_hd__buf_2
XANTENNA__14593__A _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18065__A _18206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19361__B1 _18174_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19278_ _24265_/Q _19214_/B _19277_/Y VGND VGND VPWR VPWR _19278_/X sky130_fd_sc_hd__o21a_4
XFILLER_31_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18229_ _18129_/X _18227_/X _24468_/Q _18228_/X VGND VGND VPWR VPWR _18229_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22248__B1 _14898_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15201__B _15146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22799__A1 _17383_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21240_ _21239_/X _21235_/X _12270_/B _21230_/X VGND VGND VPWR VPWR _23926_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13002__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21171_ _20339_/X _21169_/X _23964_/Q _21166_/X VGND VGND VPWR VPWR _23964_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13937__A _13611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12751__A3 _12715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12841__A _11657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21471__B2 _21467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16313__A _13415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20122_ _20110_/Y _20121_/Y _20103_/X _18940_/A VGND VGND VPWR VPWR _20122_/X sky130_fd_sc_hd__a211o_4
XANTENNA__13656__B _13745_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20053_ _20053_/A VGND VGND VPWR VPWR _20053_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19967__A2 _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21774__A2 _21769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15871__B _15802_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14768__A _13600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13672__A _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23812_ _23812_/CLK _23812_/D VGND VGND VPWR VPWR _14696_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17144__A _16514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24244__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22985__A _22985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23743_ _23889_/CLK _23743_/D VGND VGND VPWR VPWR _23743_/Q sky130_fd_sc_hd__dfxtp_4
X_20955_ _20282_/A _20955_/B VGND VGND VPWR VPWR _20955_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12288__A _12688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16983__A _16945_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ _23706_/CLK _21696_/X VGND VGND VPWR VPWR _16472_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20825_/X _20886_/B VGND VGND VPWR VPWR _20886_/Y sky130_fd_sc_hd__nor2_4
XFILLER_39_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22625_ _22396_/X _22622_/X _16788_/B _22619_/X VGND VGND VPWR VPWR _23131_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22487__B1 _12983_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11920__A _11993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22556_ _22449_/X _22550_/X _14505_/B _22554_/X VGND VGND VPWR VPWR _22556_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21507_ _21556_/A VGND VGND VPWR VPWR _21532_/A sky130_fd_sc_hd__buf_2
X_22487_ _22415_/X _22486_/X _12983_/B _22483_/X VGND VGND VPWR VPWR _23219_/D sky130_fd_sc_hd__o22a_4
X_12240_ _12240_/A VGND VGND VPWR VPWR _12240_/X sky130_fd_sc_hd__buf_2
X_24226_ _24229_/CLK _19353_/X HRESETn VGND VGND VPWR VPWR _20932_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21438_ _21277_/X _21433_/X _14309_/B _21437_/X VGND VGND VPWR VPWR _21438_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12171_ _11829_/A _23869_/Q VGND VGND VPWR VPWR _12172_/C sky130_fd_sc_hd__or2_4
X_21369_ _21369_/A VGND VGND VPWR VPWR _21369_/X sky130_fd_sc_hd__buf_2
X_24157_ _24293_/CLK _24157_/D HRESETn VGND VGND VPWR VPWR _24157_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17319__A _17143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21462__B2 _21460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23108_ _23812_/CLK _23108_/D VGND VGND VPWR VPWR _14695_/B sky130_fd_sc_hd__dfxtp_4
X_24088_ _24088_/CLK _24088_/D VGND VGND VPWR VPWR _24088_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12470__B _24021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15930_ _15929_/X VGND VGND VPWR VPWR _16095_/A sky130_fd_sc_hd__buf_2
XFILLER_77_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23039_ _23018_/A _23037_/X _23039_/C VGND VGND VPWR VPWR _23039_/X sky130_fd_sc_hd__and3_4
XFILLER_103_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21765__A2 _21762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15861_ _13548_/X _15861_/B VGND VGND VPWR VPWR _15862_/C sky130_fd_sc_hd__or2_4
XANTENNA__23056__A _23051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17600_ _17416_/A _17599_/Y _17408_/Y _17419_/Y VGND VGND VPWR VPWR _17600_/X sky130_fd_sc_hd__a211o_4
XFILLER_97_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14812_ _13690_/A _14809_/X _14811_/X VGND VGND VPWR VPWR _14812_/X sky130_fd_sc_hd__and3_4
XFILLER_40_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18580_ _17335_/X _17308_/X VGND VGND VPWR VPWR _18630_/A sky130_fd_sc_hd__and2_4
X_15792_ _15785_/A _15792_/B VGND VGND VPWR VPWR _15793_/C sky130_fd_sc_hd__or2_4
XFILLER_79_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17531_ _18153_/A _17514_/Y _17522_/Y _17530_/Y VGND VGND VPWR VPWR _17531_/X sky130_fd_sc_hd__a211o_4
X_14743_ _13799_/A _14743_/B VGND VGND VPWR VPWR _14744_/C sky130_fd_sc_hd__or2_4
XANTENNA__17989__A _18216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11955_ _11955_/A VGND VGND VPWR VPWR _15533_/A sky130_fd_sc_hd__buf_2
XANTENNA__20725__B1 _24075_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12198__A _13631_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16893__A _16893_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17462_ _17461_/X VGND VGND VPWR VPWR _18138_/B sky130_fd_sc_hd__inv_2
X_14674_ _14341_/A _14674_/B VGND VGND VPWR VPWR _14677_/B sky130_fd_sc_hd__or2_4
XFILLER_60_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11886_ _16286_/A VGND VGND VPWR VPWR _11886_/X sky130_fd_sc_hd__buf_2
XFILLER_72_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16413_ _15999_/X _16413_/B VGND VGND VPWR VPWR _16413_/X sky130_fd_sc_hd__or2_4
X_19201_ _19108_/A VGND VGND VPWR VPWR _19201_/X sky130_fd_sc_hd__buf_2
XFILLER_32_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13625_ _13813_/A _13621_/X _13625_/C VGND VGND VPWR VPWR _13625_/X sky130_fd_sc_hd__or3_4
XANTENNA__22478__B1 _16289_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17393_ _18760_/C _17413_/B VGND VGND VPWR VPWR _17393_/X sky130_fd_sc_hd__or2_4
XANTENNA__12926__A _12926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19132_ _19132_/A _19132_/B VGND VGND VPWR VPWR _19132_/X sky130_fd_sc_hd__and2_4
XFILLER_38_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16344_ _16365_/A _24057_/Q VGND VGND VPWR VPWR _16345_/C sky130_fd_sc_hd__or2_4
XFILLER_92_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23761__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13556_ _13494_/X _13550_/X _13556_/C VGND VGND VPWR VPWR _13556_/X sky130_fd_sc_hd__or3_4
XFILLER_41_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12507_ _13031_/A _12620_/B VGND VGND VPWR VPWR _12507_/X sky130_fd_sc_hd__or2_4
X_19063_ _19052_/X _19061_/Y _19062_/Y _19057_/X VGND VGND VPWR VPWR _19063_/X sky130_fd_sc_hd__o22a_4
X_16275_ _16243_/X _23609_/Q VGND VGND VPWR VPWR _16275_/X sky130_fd_sc_hd__or2_4
X_13487_ _12497_/X _13487_/B VGND VGND VPWR VPWR _13487_/X sky130_fd_sc_hd__or2_4
X_18014_ _17646_/A _18014_/B VGND VGND VPWR VPWR _18014_/Y sky130_fd_sc_hd__nand2_4
X_15226_ _14182_/A _23809_/Q VGND VGND VPWR VPWR _15226_/X sky130_fd_sc_hd__or2_4
X_12438_ _13925_/A VGND VGND VPWR VPWR _12439_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24117__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13757__A _15494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15157_ _11909_/A _15157_/B _15156_/X VGND VGND VPWR VPWR _15161_/B sky130_fd_sc_hd__and3_4
X_12369_ _12381_/A _12271_/B VGND VGND VPWR VPWR _12370_/C sky130_fd_sc_hd__or2_4
XFILLER_5_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12661__A _12622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16133__A _16109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14108_ _14108_/A _14108_/B _14108_/C VGND VGND VPWR VPWR _14118_/B sky130_fd_sc_hd__and3_4
XANTENNA__21974__A _21988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15088_ _14068_/A _15088_/B VGND VGND VPWR VPWR _15088_/X sky130_fd_sc_hd__or2_4
X_19965_ _19964_/X VGND VGND VPWR VPWR _19965_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15972__A _11980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14039_ _14039_/A _14019_/X _14039_/C VGND VGND VPWR VPWR _14039_/X sky130_fd_sc_hd__or3_4
X_18916_ _14851_/X _18912_/X _19089_/A _18913_/X VGND VGND VPWR VPWR _24355_/D sky130_fd_sc_hd__o22a_4
XFILLER_86_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16880__B2 _16816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21205__B2 _21201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22402__B1 _16240_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19896_ _22978_/A VGND VGND VPWR VPWR _23027_/A sky130_fd_sc_hd__buf_2
XFILLER_110_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21756__A2 _21755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20413__C1 _20412_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18847_ _15646_/X _18841_/X _24395_/Q _18842_/X VGND VGND VPWR VPWR _24395_/D sky130_fd_sc_hd__o22a_4
XFILLER_7_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18778_ _16233_/X _18774_/X _20427_/A _18775_/X VGND VGND VPWR VPWR _24439_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20102__B _20090_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22705__B2 _22704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17729_ _16965_/C _17106_/X VGND VGND VPWR VPWR _17729_/X sky130_fd_sc_hd__or2_4
XANTENNA__17899__A _18203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22181__A2 _22179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20740_ _20732_/X _20738_/X _24298_/Q _20739_/X VGND VGND VPWR VPWR _20741_/B sky130_fd_sc_hd__o22a_4
XANTENNA__21214__A _21112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20671_ _21831_/A VGND VGND VPWR VPWR _20671_/X sky130_fd_sc_hd__buf_2
XFILLER_91_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11740__A _11740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24390__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22410_ _20486_/A VGND VGND VPWR VPWR _22410_/X sky130_fd_sc_hd__buf_2
XFILLER_91_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23390_ _23326_/CLK _22206_/X VGND VGND VPWR VPWR _11813_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21141__B1 _15667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22341_ _22075_/X _22340_/X _12132_/B _22337_/X VGND VGND VPWR VPWR _23293_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20495__A2 _20405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21692__B2 _21688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22272_ _22272_/A VGND VGND VPWR VPWR _22272_/X sky130_fd_sc_hd__buf_2
XANTENNA__22045__A _22031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21223_ _21247_/A VGND VGND VPWR VPWR _21223_/X sky130_fd_sc_hd__buf_2
X_24011_ _24011_/CLK _21094_/X VGND VGND VPWR VPWR _24011_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13667__A _15412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12571__A _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21444__B2 _21401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22641__B1 _13325_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21154_ _21118_/A VGND VGND VPWR VPWR _21154_/X sky130_fd_sc_hd__buf_2
XFILLER_105_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15123__A1 _15051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21884__A _21884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12290__B _24054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16978__A _17681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24356__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20105_ _20105_/A _20104_/X _19027_/A VGND VGND VPWR VPWR _20105_/X sky130_fd_sc_hd__and3_4
XANTENNA__15882__A _15882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19354__A _19317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21085_ _20574_/X _21082_/X _24017_/Q _21079_/X VGND VGND VPWR VPWR _24017_/D sky130_fd_sc_hd__o22a_4
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21747__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20036_ _20018_/X _18383_/A _20024_/X _20035_/X VGND VGND VPWR VPWR _20037_/A sky130_fd_sc_hd__o22a_4
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23634__CLK _23155_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_12_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11915__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19801__B _19775_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15106__B _23839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21987_ _21814_/X _21981_/X _23508_/Q _21985_/X VGND VGND VPWR VPWR _21987_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18376__B2 _18375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11740_/A VGND VGND VPWR VPWR _12613_/A sky130_fd_sc_hd__buf_2
X_23726_ _23922_/CLK _23726_/D VGND VGND VPWR VPWR _15656_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_15_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23784__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20872_/X _20937_/X _15297_/B _20839_/X VGND VGND VPWR VPWR _24066_/D sky130_fd_sc_hd__o22a_4
XFILLER_57_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11671_/A VGND VGND VPWR VPWR _13133_/A sky130_fd_sc_hd__buf_2
X_23657_ _23847_/CLK _23657_/D VGND VGND VPWR VPWR _23657_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _22134_/A VGND VGND VPWR VPWR _20870_/A sky130_fd_sc_hd__buf_2
XFILLER_39_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12746__A _12315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13383_/A _13341_/B VGND VGND VPWR VPWR _13410_/X sky130_fd_sc_hd__or2_4
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22608_ _22451_/X _22607_/X _14674_/B _22604_/X VGND VGND VPWR VPWR _23140_/D sky130_fd_sc_hd__o22a_4
X_14390_ _15614_/A _14301_/B VGND VGND VPWR VPWR _14390_/X sky130_fd_sc_hd__or2_4
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23588_ _23907_/CLK _23588_/D VGND VGND VPWR VPWR _14691_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13341_ _15697_/A _13341_/B VGND VGND VPWR VPWR _13341_/X sky130_fd_sc_hd__or2_4
X_22539_ _22420_/X _22536_/X _13144_/B _22533_/X VGND VGND VPWR VPWR _22539_/X sky130_fd_sc_hd__o22a_4
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16060_ _16215_/A _16060_/B _16060_/C VGND VGND VPWR VPWR _16076_/B sky130_fd_sc_hd__and3_4
X_13272_ _13202_/X _13272_/B VGND VGND VPWR VPWR _13272_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15011_ _15011_/A _23551_/Q VGND VGND VPWR VPWR _15011_/X sky130_fd_sc_hd__or2_4
X_12223_ _12211_/X VGND VGND VPWR VPWR _12691_/A sky130_fd_sc_hd__buf_2
X_24209_ _23522_/CLK _24209_/D HRESETn VGND VGND VPWR VPWR _24209_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13577__A _13493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21435__A1 _21273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21435__B2 _21430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22632__B1 _12293_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12481__A _12556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12154_ _11748_/X _12152_/X _12154_/C VGND VGND VPWR VPWR _12154_/X sky130_fd_sc_hd__and3_4
XFILLER_1_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15792__A _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19750_ _19447_/X _19749_/X _16677_/A _19493_/X VGND VGND VPWR VPWR _19750_/Y sky130_fd_sc_hd__a22oi_4
X_12085_ _12044_/X _12085_/B _12085_/C VGND VGND VPWR VPWR _12089_/B sky130_fd_sc_hd__and3_4
X_16962_ _24112_/Q VGND VGND VPWR VPWR _17734_/A sky130_fd_sc_hd__inv_2
XFILLER_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18701_ _17735_/A VGND VGND VPWR VPWR _18701_/X sky130_fd_sc_hd__buf_2
X_15913_ _15909_/X _15913_/B VGND VGND VPWR VPWR _15914_/D sky130_fd_sc_hd__nand2_4
X_16893_ _16893_/A VGND VGND VPWR VPWR _16894_/A sky130_fd_sc_hd__inv_2
X_19681_ _19553_/A HRDATA[7] VGND VGND VPWR VPWR _19681_/X sky130_fd_sc_hd__and2_4
XANTENNA__20203__A _20202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11825__A _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15844_ _12189_/X _12681_/X _15813_/X _12281_/X _15843_/X VGND VGND VPWR VPWR _15844_/X
+ sky130_fd_sc_hd__a32o_4
X_18632_ _17306_/X _18633_/B VGND VGND VPWR VPWR _18632_/Y sky130_fd_sc_hd__nand2_4
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15775_ _11741_/X _15771_/X _15774_/X VGND VGND VPWR VPWR _15775_/X sky130_fd_sc_hd__or3_4
X_18563_ _17422_/A _18561_/X VGND VGND VPWR VPWR _18563_/Y sky130_fd_sc_hd__nand2_4
XFILLER_80_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12987_ _13083_/A _12987_/B _12987_/C VGND VGND VPWR VPWR _12988_/C sky130_fd_sc_hd__and3_4
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19564__B1 HRDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14726_ _11894_/A _14788_/B VGND VGND VPWR VPWR _14727_/C sky130_fd_sc_hd__or2_4
X_17514_ _17476_/X _17514_/B VGND VGND VPWR VPWR _17514_/Y sky130_fd_sc_hd__nor2_4
X_11938_ _11993_/A _11749_/B VGND VGND VPWR VPWR _11940_/B sky130_fd_sc_hd__or2_4
X_18494_ _17422_/C _18493_/X VGND VGND VPWR VPWR _18494_/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21910__A2 _21908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17445_ _17444_/X VGND VGND VPWR VPWR _17447_/A sky130_fd_sc_hd__inv_2
XFILLER_21_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21034__A _21027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14657_ _11738_/A VGND VGND VPWR VPWR _14658_/A sky130_fd_sc_hd__buf_2
XFILLER_53_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11869_ _13624_/A VGND VGND VPWR VPWR _12465_/A sky130_fd_sc_hd__buf_2
XANTENNA__12656__A _13118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13608_ _13608_/A _13698_/B VGND VGND VPWR VPWR _13608_/X sky130_fd_sc_hd__or2_4
XANTENNA__15032__A _15032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17376_ _15910_/Y _17013_/A _17021_/A _17375_/X VGND VGND VPWR VPWR _17377_/B sky130_fd_sc_hd__o22a_4
XANTENNA__21969__A _22002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14588_ _15013_/A VGND VGND VPWR VPWR _14588_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20873__A _20512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16327_ _11713_/X VGND VGND VPWR VPWR _16365_/A sky130_fd_sc_hd__buf_2
X_19115_ _24294_/Q _19115_/B VGND VGND VPWR VPWR _19116_/B sky130_fd_sc_hd__and2_4
XFILLER_119_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13539_ _15876_/A _23887_/Q VGND VGND VPWR VPWR _13539_/X sky130_fd_sc_hd__or2_4
XANTENNA__15967__A _15959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21674__B2 _21673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23507__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19046_ _19002_/A VGND VGND VPWR VPWR _19046_/X sky130_fd_sc_hd__buf_2
X_16258_ _15936_/A _16256_/X _16257_/X VGND VGND VPWR VPWR _16258_/X sky130_fd_sc_hd__and3_4
XANTENNA__15686__B _15686_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15209_ _11708_/A VGND VGND VPWR VPWR _15234_/A sky130_fd_sc_hd__buf_2
XANTENNA__13487__A _12497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16189_ _16227_/A _16189_/B VGND VGND VPWR VPWR _16189_/X sky130_fd_sc_hd__or2_4
XFILLER_12_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12391__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21977__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19948_ _17631_/X VGND VGND VPWR VPWR _19948_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21729__A2 _21726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19879_ _19878_/X VGND VGND VPWR VPWR _19879_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21910_ _21855_/X _21908_/X _14803_/B _21905_/X VGND VGND VPWR VPWR _23555_/D sky130_fd_sc_hd__o22a_4
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22890_ _20196_/A VGND VGND VPWR VPWR _23015_/A sky130_fd_sc_hd__buf_2
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21841_ _21792_/A VGND VGND VPWR VPWR _21841_/X sky130_fd_sc_hd__buf_2
XFILLER_82_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21772_ _21560_/X _21769_/X _13825_/B _21766_/X VGND VGND VPWR VPWR _21772_/X sky130_fd_sc_hd__o22a_4
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23511_ _23635_/CLK _23511_/D VGND VGND VPWR VPWR _23511_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20723_ _21265_/A VGND VGND VPWR VPWR _20723_/X sky130_fd_sc_hd__buf_2
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12566__A _14002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19307__B1 _17040_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23442_ _23922_/CLK _23442_/D VGND VGND VPWR VPWR _13091_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20654_ _20425_/A VGND VGND VPWR VPWR _20654_/X sky130_fd_sc_hd__buf_2
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_3_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15877__A _15884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20585_ _18334_/X _20447_/X _20492_/X _20584_/Y VGND VGND VPWR VPWR _20585_/X sky130_fd_sc_hd__a211o_4
X_23373_ _23826_/CLK _22231_/X VGND VGND VPWR VPWR _15824_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21665__B2 _21659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14781__A _12217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22324_ _14287_/B VGND VGND VPWR VPWR _22324_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21417__B2 _21416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22255_ _22262_/A VGND VGND VPWR VPWR _22255_/X sky130_fd_sc_hd__buf_2
X_21206_ _20916_/X _21204_/X _14820_/B _21201_/X VGND VGND VPWR VPWR _21206_/X sky130_fd_sc_hd__o22a_4
X_22186_ _22153_/A VGND VGND VPWR VPWR _22186_/X sky130_fd_sc_hd__buf_2
XFILLER_79_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17636__A3 _17260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19084__A _18999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21137_ _21130_/A VGND VGND VPWR VPWR _21137_/X sky130_fd_sc_hd__buf_2
XANTENNA__16501__A _16159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18046__B1 _18425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21068_ _21075_/A VGND VGND VPWR VPWR _21068_/X sky130_fd_sc_hd__buf_2
XFILLER_24_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21119__A _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22393__A2 _22392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ _12910_/A _12910_/B _12910_/C VGND VGND VPWR VPWR _12914_/B sky130_fd_sc_hd__and3_4
X_20019_ _24465_/Q VGND VGND VPWR VPWR _20019_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11645__A _11645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15117__A _14040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19812__A _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13890_ _13890_/A _23591_/Q VGND VGND VPWR VPWR _13892_/B sky130_fd_sc_hd__or2_4
XFILLER_73_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14021__A _14021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20958__A _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12841_ _11657_/X _12841_/B _12841_/C VGND VGND VPWR VPWR _12841_/X sky130_fd_sc_hd__and3_4
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19546__B1 _19497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13860__A _14002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15560_ _15533_/A _15560_/B VGND VGND VPWR VPWR _15560_/X sky130_fd_sc_hd__or2_4
X_12772_ _12954_/A VGND VGND VPWR VPWR _13563_/A sky130_fd_sc_hd__buf_2
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14536_/A _14511_/B VGND VGND VPWR VPWR _14512_/C sky130_fd_sc_hd__or2_4
XFILLER_70_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11723_/A VGND VGND VPWR VPWR _12412_/A sky130_fd_sc_hd__buf_2
X_23709_ _23707_/CLK _23709_/D VGND VGND VPWR VPWR _23709_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15491_/A _15491_/B _15491_/C VGND VGND VPWR VPWR _15492_/C sky130_fd_sc_hd__and3_4
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__A _13020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_19_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR _24216_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17152_/X _17228_/X _17163_/X _17229_/X VGND VGND VPWR VPWR _17230_/X sky130_fd_sc_hd__o22a_4
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _12878_/A _14442_/B VGND VGND VPWR VPWR _14444_/B sky130_fd_sc_hd__or2_4
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _14073_/A VGND VGND VPWR VPWR _13918_/A sky130_fd_sc_hd__buf_2
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17161_ _17161_/A VGND VGND VPWR VPWR _17161_/X sky130_fd_sc_hd__buf_2
XANTENNA__15787__A _12443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21656__A1 _21531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14373_ _15601_/A _14373_/B VGND VGND VPWR VPWR _14373_/X sky130_fd_sc_hd__or2_4
XANTENNA__21656__B2 _21652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ _11585_/A VGND VGND VPWR VPWR _17009_/A sky130_fd_sc_hd__buf_2
XFILLER_11_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16112_ _16140_/A _16112_/B _16111_/X VGND VGND VPWR VPWR _16113_/C sky130_fd_sc_hd__and3_4
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _13483_/A _13320_/X _13324_/C VGND VGND VPWR VPWR _13324_/X sky130_fd_sc_hd__or3_4
X_17092_ _17057_/A _17073_/X VGND VGND VPWR VPWR _18656_/A sky130_fd_sc_hd__or2_4
XFILLER_10_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16043_ _11684_/X _16043_/B _16042_/X VGND VGND VPWR VPWR _16044_/C sky130_fd_sc_hd__or3_4
XANTENNA__21408__A1 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13255_ _13243_/A _13253_/X _13255_/C VGND VGND VPWR VPWR _13255_/X sky130_fd_sc_hd__and3_4
XANTENNA__21408__B2 _21402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12206_ _12553_/A _12206_/B VGND VGND VPWR VPWR _12206_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11539__B IRQ[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13186_ _12739_/A _24081_/Q VGND VGND VPWR VPWR _13187_/C sky130_fd_sc_hd__or2_4
XANTENNA__22413__A _22413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19802_ _19754_/A _19801_/X _19523_/A _19861_/A VGND VGND VPWR VPWR _19802_/X sky130_fd_sc_hd__a211o_4
XFILLER_96_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12137_ _12168_/A _23581_/Q VGND VGND VPWR VPWR _12138_/C sky130_fd_sc_hd__or2_4
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13649__A1 _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17994_ _18047_/A _17993_/X _17574_/Y VGND VGND VPWR VPWR _17994_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_97_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16411__A _11980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19733_ _19643_/A _19731_/X _19580_/X _19732_/X VGND VGND VPWR VPWR _19733_/X sky130_fd_sc_hd__a211o_4
X_12068_ _11966_/X VGND VGND VPWR VPWR _12068_/X sky130_fd_sc_hd__buf_2
X_16945_ _24131_/Q VGND VGND VPWR VPWR _16945_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18588__A1 _18500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15027__A _14151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19722__A _19722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19664_ _19599_/B VGND VGND VPWR VPWR _19793_/B sky130_fd_sc_hd__buf_2
X_16876_ _16876_/A _16872_/X _16876_/C _16876_/D VGND VGND VPWR VPWR _16876_/X sky130_fd_sc_hd__and4_4
XFILLER_4_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20395__B2 _20374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21592__B1 _23741_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18615_ _17792_/A _18578_/X _18189_/A _18581_/X VGND VGND VPWR VPWR _18615_/X sky130_fd_sc_hd__o22a_4
X_15827_ _12458_/A _15823_/X _15827_/C VGND VGND VPWR VPWR _15827_/X sky130_fd_sc_hd__or3_4
XFILLER_20_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19595_ _24145_/Q _19435_/X HRDATA[19] _19432_/X VGND VGND VPWR VPWR _19595_/X sky130_fd_sc_hd__o22a_4
XFILLER_111_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13770__A _13770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21353__A2_N _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15758_ _15751_/A _15758_/B VGND VGND VPWR VPWR _15758_/X sky130_fd_sc_hd__or2_4
X_18546_ _17397_/X _18544_/X _17878_/X _18545_/X VGND VGND VPWR VPWR _18547_/A sky130_fd_sc_hd__a211o_4
XFILLER_20_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21344__B1 _23873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14709_ _15589_/A _14705_/X _14708_/X VGND VGND VPWR VPWR _14709_/X sky130_fd_sc_hd__or3_4
X_15689_ _15689_/A _15689_/B VGND VGND VPWR VPWR _15691_/B sky130_fd_sc_hd__or2_4
X_18477_ _17703_/X _17750_/X _17703_/X _17750_/X VGND VGND VPWR VPWR _18477_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12386__A _12926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21895__B2 _21891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24455__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17428_ _17422_/D _17426_/X _17427_/X VGND VGND VPWR VPWR _17428_/X sky130_fd_sc_hd__o21a_4
XFILLER_21_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15697__A _15697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21647__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17359_ _17191_/X _17432_/B VGND VGND VPWR VPWR _17360_/A sky130_fd_sc_hd__or2_4
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20370_ _20370_/A _20369_/X VGND VGND VPWR VPWR _20370_/Y sky130_fd_sc_hd__nand2_4
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16305__B _23513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19029_ _19016_/X _19028_/X _19016_/X _11519_/A VGND VGND VPWR VPWR _19029_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14106__A _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22040_ _21819_/X _22038_/X _23474_/Q _22035_/X VGND VGND VPWR VPWR _22040_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13010__A _12917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22323__A _13794_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13945__A _13643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23991_ _23316_/CLK _23991_/D VGND VGND VPWR VPWR _23991_/Q sky130_fd_sc_hd__dfxtp_4
X_22942_ _22924_/X _18348_/A _22937_/X _22941_/X VGND VGND VPWR VPWR _22943_/A sky130_fd_sc_hd__a211o_4
XFILLER_116_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20778__A _20778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22873_ _19893_/X _22815_/X _15453_/Y _22855_/A VGND VGND VPWR VPWR _22873_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14776__A _13959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13680__A _15448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21824_ _21812_/A VGND VGND VPWR VPWR _21824_/X sky130_fd_sc_hd__buf_2
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22993__A _18283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21755_ _21755_/A VGND VGND VPWR VPWR _21755_/X sky130_fd_sc_hd__buf_2
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21886__B2 _21884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12296__A _12742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20706_ _20706_/A VGND VGND VPWR VPWR _20708_/A sky130_fd_sc_hd__inv_2
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24474_ _24473_/CLK _24474_/D HRESETn VGND VGND VPWR VPWR _19977_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21686_ _21690_/A VGND VGND VPWR VPWR _21702_/A sky130_fd_sc_hd__inv_2
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23425_ _23104_/CLK _23425_/D VGND VGND VPWR VPWR _15150_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23822__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21402__A _21401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20637_ _21543_/A VGND VGND VPWR VPWR _20637_/X sky130_fd_sc_hd__buf_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15400__A _13620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23356_ _23100_/CLK _22260_/X VGND VGND VPWR VPWR _16608_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20310__A1 _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20568_ _20568_/A VGND VGND VPWR VPWR _20568_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20018__A _19994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12743__B _23796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22307_ _22307_/A VGND VGND VPWR VPWR _23319_/D sky130_fd_sc_hd__buf_2
XANTENNA__20861__A2 _20860_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23287_ _23473_/CLK _23287_/D VGND VGND VPWR VPWR _16103_/B sky130_fd_sc_hd__dfxtp_4
X_20499_ _20494_/X _20498_/X _24340_/Q _20453_/X VGND VGND VPWR VPWR _20499_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20960__B HRDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13040_ _13017_/A _13040_/B _13040_/C VGND VGND VPWR VPWR _13041_/C sky130_fd_sc_hd__and3_4
XFILLER_4_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22238_ _22127_/X _22236_/X _13664_/B _22233_/X VGND VGND VPWR VPWR _23368_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22063__B2 _22020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22233__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13855__A _13710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22169_ _22169_/A VGND VGND VPWR VPWR _22169_/X sky130_fd_sc_hd__buf_2
XANTENNA__21810__B2 _21800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16231__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18019__B1 _18016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23202__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14991_ _14991_/A _14991_/B _14991_/C VGND VGND VPWR VPWR _14995_/B sky130_fd_sc_hd__and3_4
XANTENNA__22366__A2 _22361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13942_ _13966_/A _23658_/Q VGND VGND VPWR VPWR _13942_/X sky130_fd_sc_hd__or2_4
X_16730_ _12093_/A _16806_/B VGND VGND VPWR VPWR _16730_/X sky130_fd_sc_hd__or2_4
XFILLER_43_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20377__A1 _20285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16661_ _16624_/X _16661_/B _16660_/X VGND VGND VPWR VPWR _16661_/X sky130_fd_sc_hd__and3_4
XANTENNA__23064__A _22898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13873_ _13909_/A _13873_/B VGND VGND VPWR VPWR _13873_/X sky130_fd_sc_hd__or2_4
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22118__A2 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19519__B1 HRDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15612_ _15628_/A _15612_/B _15612_/C VGND VGND VPWR VPWR _15613_/C sky130_fd_sc_hd__and3_4
X_18400_ _18399_/Y _17423_/B _17429_/X VGND VGND VPWR VPWR _18400_/X sky130_fd_sc_hd__o21a_4
XFILLER_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12824_ _12800_/A _23796_/Q VGND VGND VPWR VPWR _12824_/X sky130_fd_sc_hd__or2_4
XANTENNA__17062__A _17062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16592_ _11924_/A _16592_/B _16592_/C VGND VGND VPWR VPWR _16592_/X sky130_fd_sc_hd__or3_4
X_19380_ _19379_/X VGND VGND VPWR VPWR _19380_/X sky130_fd_sc_hd__buf_2
XFILLER_34_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15543_ _15543_/A _23915_/Q VGND VGND VPWR VPWR _15543_/X sky130_fd_sc_hd__or2_4
X_18331_ _18216_/X _17481_/X _18329_/X _18082_/X _18330_/Y VGND VGND VPWR VPWR _18331_/X
+ sky130_fd_sc_hd__a32o_4
X_12755_ _13726_/A VGND VGND VPWR VPWR _13088_/A sky130_fd_sc_hd__buf_2
XANTENNA__17997__A _18048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11644_/A VGND VGND VPWR VPWR _11707_/A sky130_fd_sc_hd__inv_2
X_18262_ _18235_/A _22992_/B _18237_/A VGND VGND VPWR VPWR _18262_/X sky130_fd_sc_hd__o21a_4
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _15512_/A _15474_/B VGND VGND VPWR VPWR _15474_/X sky130_fd_sc_hd__or2_4
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12284_/X _12767_/B VGND VGND VPWR VPWR _12686_/X sky130_fd_sc_hd__or2_4
XANTENNA__22408__A _20463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _14425_/A VGND VGND VPWR VPWR _14428_/A sky130_fd_sc_hd__inv_2
X_17213_ _12676_/X _17137_/X _17179_/Y _17138_/X VGND VGND VPWR VPWR _17213_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21312__A _21319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _11737_/A VGND VGND VPWR VPWR _11638_/A sky130_fd_sc_hd__buf_2
X_18193_ _18176_/X _18181_/Y _18188_/X _18191_/X _18192_/Y VGND VGND VPWR VPWR _18193_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21629__B2 _21623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16406__A _13447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12934__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17144_ _16514_/X VGND VGND VPWR VPWR _17144_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15310__A _14172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _15584_/A _14276_/B VGND VGND VPWR VPWR _14356_/X sky130_fd_sc_hd__or2_4
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11568_ _11565_/X _11567_/X VGND VGND VPWR VPWR _20090_/B sky130_fd_sc_hd__or2_4
XFILLER_89_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13307_ _12503_/A _13302_/X _13306_/X VGND VGND VPWR VPWR _13307_/X sky130_fd_sc_hd__or3_4
XFILLER_13_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17075_ _18498_/A VGND VGND VPWR VPWR _18418_/A sky130_fd_sc_hd__buf_2
X_14287_ _15536_/A _14287_/B VGND VGND VPWR VPWR _14290_/B sky130_fd_sc_hd__or2_4
XANTENNA__18621__A _18137_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16026_ _16050_/A _15952_/B VGND VGND VPWR VPWR _16026_/X sky130_fd_sc_hd__or2_4
XANTENNA__22054__A1 _21843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13238_ _12791_/A _13171_/B VGND VGND VPWR VPWR _13240_/B sky130_fd_sc_hd__or2_4
XANTENNA__22054__B2 _22049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22143__A _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13169_ _15812_/A _13168_/X VGND VGND VPWR VPWR _13169_/X sky130_fd_sc_hd__and2_4
XANTENNA__21801__B2 _21800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17977_ _17818_/X _17839_/X _17813_/X _17830_/X VGND VGND VPWR VPWR _17978_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22357__A2 _22354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19758__B1 _19481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19716_ _19597_/A _19714_/X _19581_/X _19715_/Y VGND VGND VPWR VPWR _19716_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15980__A _15980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19452__A _19416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16928_ _17285_/A VGND VGND VPWR VPWR _16929_/B sky130_fd_sc_hd__buf_2
XFILLER_61_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19647_ _19862_/A _19857_/C _19578_/X _19646_/X VGND VGND VPWR VPWR _19647_/X sky130_fd_sc_hd__a211o_4
X_16859_ _15051_/X _15119_/X _15123_/Y _15385_/X VGND VGND VPWR VPWR _16859_/X sky130_fd_sc_hd__a211o_4
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22109__A2 _22101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19701__A2_N _19699_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19578_ _19722_/A _19536_/A _19537_/B VGND VGND VPWR VPWR _19578_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21317__B1 _12639_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18529_ _18458_/X _18518_/Y _18485_/X _18528_/X VGND VGND VPWR VPWR _18529_/X sky130_fd_sc_hd__o22a_4
XFILLER_80_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13005__A _12879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21540_ _21538_/X _21532_/X _23760_/Q _21539_/X VGND VGND VPWR VPWR _21540_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20540__A1 _20229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21471_ _21246_/X _21470_/X _12974_/B _21467_/X VGND VGND VPWR VPWR _21471_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_65_0_HCLK clkbuf_7_65_0_HCLK/A VGND VGND VPWR VPWR _24290_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16316__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23210_ _23561_/CLK _23210_/D VGND VGND VPWR VPWR _14066_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15220__A _14195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20422_ _18757_/X VGND VGND VPWR VPWR _20422_/X sky130_fd_sc_hd__buf_2
XANTENNA__23995__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24190_ _24187_/CLK _24190_/D HRESETn VGND VGND VPWR VPWR _24190_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23141_ _23557_/CLK _22606_/X VGND VGND VPWR VPWR _14518_/B sky130_fd_sc_hd__dfxtp_4
X_20353_ _20370_/A _20353_/B VGND VGND VPWR VPWR _20353_/Y sky130_fd_sc_hd__nand2_4
X_20284_ _20212_/X VGND VGND VPWR VPWR _20284_/X sky130_fd_sc_hd__buf_2
X_23072_ _24180_/CLK _23072_/D VGND VGND VPWR VPWR _14909_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_115_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22596__A2 _22593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22023_ _22052_/A VGND VGND VPWR VPWR _22031_/A sky130_fd_sc_hd__buf_2
XFILLER_114_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22988__A _18309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_25_0_HCLK_A clkbuf_5_24_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22348__A2 _22347_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15890__A _13557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23974_ _23845_/CLK _23974_/D VGND VGND VPWR VPWR _14379_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22925_ _23048_/A VGND VGND VPWR VPWR _22952_/A sky130_fd_sc_hd__buf_2
XFILLER_21_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20301__A _20301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22856_ _22854_/X _22798_/X _17383_/Y _22855_/X VGND VGND VPWR VPWR _22856_/X sky130_fd_sc_hd__o22a_4
XFILLER_71_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21807_ _20442_/A VGND VGND VPWR VPWR _21807_/X sky130_fd_sc_hd__buf_2
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22787_ _14786_/Y _22782_/X VGND VGND VPWR VPWR HWDATA[4] sky130_fd_sc_hd__nor2_4
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18724__B2 _18723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12540_ _12540_/A _12540_/B _12540_/C VGND VGND VPWR VPWR _12541_/C sky130_fd_sc_hd__and3_4
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21738_ _21737_/X VGND VGND VPWR VPWR _21738_/X sky130_fd_sc_hd__buf_2
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12471_ _12880_/A VGND VGND VPWR VPWR _12472_/A sky130_fd_sc_hd__buf_2
X_24457_ _24203_/CLK _24457_/D HRESETn VGND VGND VPWR VPWR _20058_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21669_ _21636_/A VGND VGND VPWR VPWR _21669_/X sky130_fd_sc_hd__buf_2
XANTENNA__12754__A _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16226__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14210_ _14210_/A _23433_/Q VGND VGND VPWR VPWR _14210_/X sky130_fd_sc_hd__or2_4
XANTENNA__24000__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23408_ _23472_/CLK _22177_/X VGND VGND VPWR VPWR _13329_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21087__A2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15190_ _15190_/A _23713_/Q VGND VGND VPWR VPWR _15191_/C sky130_fd_sc_hd__or2_4
X_24388_ _24425_/CLK _24388_/D HRESETn VGND VGND VPWR VPWR _24388_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22284__B2 _22283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14141_ _14108_/A _14141_/B _14141_/C VGND VGND VPWR VPWR _14145_/B sky130_fd_sc_hd__and3_4
X_23339_ _24011_/CLK _22284_/X VGND VGND VPWR VPWR _23339_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20834__A2 _20824_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14072_ _14040_/X _14072_/B _14072_/C VGND VGND VPWR VPWR _14073_/C sky130_fd_sc_hd__or3_4
XFILLER_84_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22036__B2 _22035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15784__B _15845_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24150__CLK _24162_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13023_ _12512_/A _13091_/B VGND VGND VPWR VPWR _13024_/C sky130_fd_sc_hd__or2_4
X_17900_ _17900_/A VGND VGND VPWR VPWR _18264_/A sky130_fd_sc_hd__buf_2
XANTENNA__22587__A2 _22586_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17057__A _17057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18880_ _12184_/X _18875_/X _18930_/A _18878_/X VGND VGND VPWR VPWR _24381_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20598__A1 _20425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22898__A _22898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20598__B2 _20473_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17831_ _17826_/X _17196_/X _17815_/X _17187_/X VGND VGND VPWR VPWR _17831_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17762_ _17755_/A _17692_/Y _18164_/A _17761_/X VGND VGND VPWR VPWR _17762_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14974_ _11709_/A _23840_/Q VGND VGND VPWR VPWR _14975_/C sky130_fd_sc_hd__or2_4
XANTENNA__21547__B1 _15792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19501_ _19477_/A VGND VGND VPWR VPWR _19572_/C sky130_fd_sc_hd__inv_2
XFILLER_75_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16713_ _16713_/A _23899_/Q VGND VGND VPWR VPWR _16715_/B sky130_fd_sc_hd__or2_4
XFILLER_78_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13925_ _13925_/A _13995_/B VGND VGND VPWR VPWR _13925_/X sky130_fd_sc_hd__or2_4
X_17693_ _17694_/A _17367_/X VGND VGND VPWR VPWR _17697_/A sky130_fd_sc_hd__or2_4
XANTENNA__12929__A _12640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19432_ _19431_/X VGND VGND VPWR VPWR _19432_/X sky130_fd_sc_hd__buf_2
XANTENNA__11833__A _11782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13856_ _13887_/A _13784_/B VGND VGND VPWR VPWR _13858_/B sky130_fd_sc_hd__or2_4
X_16644_ _16599_/X _16639_/X _16643_/X VGND VGND VPWR VPWR _16644_/X sky130_fd_sc_hd__or3_4
X_12807_ _11665_/X _12807_/B _12807_/C VGND VGND VPWR VPWR _12841_/B sky130_fd_sc_hd__or3_4
XFILLER_16_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19363_ _19361_/X VGND VGND VPWR VPWR _19363_/Y sky130_fd_sc_hd__inv_2
X_13787_ _13651_/A _13859_/B VGND VGND VPWR VPWR _13787_/X sky130_fd_sc_hd__or2_4
X_16575_ _16583_/A _16658_/B VGND VGND VPWR VPWR _16575_/X sky130_fd_sc_hd__or2_4
XANTENNA__18715__A1 _17782_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22511__A2 _22507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18314_ _18171_/A VGND VGND VPWR VPWR _18314_/X sky130_fd_sc_hd__buf_2
XFILLER_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12738_ _12738_/A _23220_/Q VGND VGND VPWR VPWR _12740_/B sky130_fd_sc_hd__or2_4
X_15526_ _15553_/A _23723_/Q VGND VGND VPWR VPWR _15526_/X sky130_fd_sc_hd__or2_4
X_19294_ _24257_/Q _19206_/B _19293_/Y VGND VGND VPWR VPWR _19294_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20522__A1 _20425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20522__B2 _20473_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15457_ _12578_/A VGND VGND VPWR VPWR _15477_/A sky130_fd_sc_hd__buf_2
X_18245_ _18245_/A VGND VGND VPWR VPWR _18245_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12669_ _12947_/A _12667_/X _12669_/C VGND VGND VPWR VPWR _12669_/X sky130_fd_sc_hd__and3_4
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14408_ _15607_/A _14406_/X _14407_/X VGND VGND VPWR VPWR _14408_/X sky130_fd_sc_hd__and3_4
X_15388_ _14724_/X _14855_/Y _15386_/X _14724_/B _15387_/X VGND VGND VPWR VPWR _15388_/X
+ sky130_fd_sc_hd__o32a_4
X_18176_ _18239_/A _18152_/A VGND VGND VPWR VPWR _18176_/X sky130_fd_sc_hd__or2_4
XANTENNA__22275__B2 _22269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14339_ _14371_/A VGND VGND VPWR VPWR _15623_/A sky130_fd_sc_hd__buf_2
X_17127_ _17126_/X VGND VGND VPWR VPWR _17127_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17058_ _17052_/X _17088_/A _11631_/A _17072_/A VGND VGND VPWR VPWR _17058_/X sky130_fd_sc_hd__a211o_4
XFILLER_48_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16009_ _16023_/A _23256_/Q VGND VGND VPWR VPWR _16009_/X sky130_fd_sc_hd__or2_4
XFILLER_98_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22578__A2 _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13495__A _12958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20589__A1 _24208_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_HCLK clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__20105__B _20104_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21250__A2 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17206__A1 _13278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21217__A _21242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20971_ _20468_/A _20970_/Y _19205_/A _20325_/X VGND VGND VPWR VPWR _20971_/X sky130_fd_sc_hd__o22a_4
XFILLER_96_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12839__A _12787_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22710_ _21287_/A _22707_/X _15303_/B _22704_/X VGND VGND VPWR VPWR _23074_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19910__A _22723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23690_ _23978_/CLK _21668_/X VGND VGND VPWR VPWR _23690_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22641_ _22422_/X _22636_/X _13325_/B _22640_/X VGND VGND VPWR VPWR _23120_/D sky130_fd_sc_hd__o22a_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22502__A2 _22500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22572_ _22586_/A VGND VGND VPWR VPWR _22572_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14773__B _14773_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24311_ _24299_/CLK _24311_/D HRESETn VGND VGND VPWR VPWR _19132_/A sky130_fd_sc_hd__dfrtp_4
X_21523_ _21522_/X _21520_/X _16171_/B _21515_/X VGND VGND VPWR VPWR _21523_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12574__A _14009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24242_ _24065_/CLK _19330_/X HRESETn VGND VGND VPWR VPWR _24242_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21887__A _21887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21454_ _21447_/Y _21453_/X _21219_/X _21453_/X VGND VGND VPWR VPWR _23806_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24173__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12293__B _12293_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11557__A2 IRQ[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20405_ _20405_/A VGND VGND VPWR VPWR _20405_/X sky130_fd_sc_hd__buf_2
XANTENNA__15885__A _13550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24173_ _24065_/CLK _19792_/X HRESETn VGND VGND VPWR VPWR _11644_/A sky130_fd_sc_hd__dfrtp_4
X_21385_ _21273_/X _21383_/X _13760_/B _21380_/X VGND VGND VPWR VPWR _21385_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17142__B1 _16814_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23124_ _23699_/CLK _22635_/X VGND VGND VPWR VPWR _23124_/Q sky130_fd_sc_hd__dfxtp_4
X_20336_ _20370_/A _20335_/X VGND VGND VPWR VPWR _20336_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__11918__A _11886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23055_ _23055_/A VGND VGND VPWR VPWR HADDR[30] sky130_fd_sc_hd__inv_2
X_20267_ _20518_/A VGND VGND VPWR VPWR _20494_/A sky130_fd_sc_hd__buf_2
X_22006_ _21985_/A VGND VGND VPWR VPWR _22006_/X sky130_fd_sc_hd__buf_2
X_20198_ _21866_/D VGND VGND VPWR VPWR _20199_/B sky130_fd_sc_hd__buf_2
XANTENNA__15109__B _15033_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11971_ _11971_/A _23550_/Q VGND VGND VPWR VPWR _11972_/C sky130_fd_sc_hd__or2_4
X_23957_ _24021_/CLK _21181_/X VGND VGND VPWR VPWR _12640_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13710_ _13710_/A VGND VGND VPWR VPWR _13911_/A sky130_fd_sc_hd__buf_2
XFILLER_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11653__A _11652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22908_ _22889_/X VGND VGND VPWR VPWR _22908_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15125__A _12202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14690_ _14673_/A _14690_/B _14689_/X VGND VGND VPWR VPWR _14690_/X sky130_fd_sc_hd__and3_4
X_23888_ _23920_/CLK _21324_/X VGND VGND VPWR VPWR _13318_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13641_ _13641_/A _23560_/Q VGND VGND VPWR VPWR _13642_/C sky130_fd_sc_hd__or2_4
XFILLER_112_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22884__C _22932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22839_ _13059_/Y _22825_/X _22831_/X _22838_/X VGND VGND VPWR VPWR _22840_/A sky130_fd_sc_hd__a211o_4
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14964__A _15063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ _11715_/A _16297_/B VGND VGND VPWR VPWR _16361_/C sky130_fd_sc_hd__or2_4
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17340__A _17012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13572_ _13572_/A _13572_/B _13572_/C VGND VGND VPWR VPWR _13573_/C sky130_fd_sc_hd__and3_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15311_ _12267_/X _15288_/X _15295_/X _15302_/X _15310_/X VGND VGND VPWR VPWR _15311_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _13019_/A VGND VGND VPWR VPWR _12915_/A sky130_fd_sc_hd__buf_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16291_ _15936_/A _16291_/B _16290_/X VGND VGND VPWR VPWR _16291_/X sky130_fd_sc_hd__and3_4
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12484__A _13643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15242_ _15203_/A _15242_/B _15241_/X VGND VGND VPWR VPWR _15242_/X sky130_fd_sc_hd__and3_4
X_18030_ _18137_/A _17550_/A VGND VGND VPWR VPWR _18030_/X sky130_fd_sc_hd__and2_4
X_12454_ _12462_/A _12580_/B VGND VGND VPWR VPWR _12454_/X sky130_fd_sc_hd__or2_4
XFILLER_51_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15173_ _14161_/A _23617_/Q VGND VGND VPWR VPWR _15173_/X sky130_fd_sc_hd__or2_4
XANTENNA__15795__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12385_ _12384_/X _12259_/B VGND VGND VPWR VPWR _12388_/B sky130_fd_sc_hd__or2_4
XANTENNA__18171__A _18171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14124_ _14992_/A _23145_/Q VGND VGND VPWR VPWR _14124_/X sky130_fd_sc_hd__or2_4
XFILLER_10_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19981_ _19981_/A VGND VGND VPWR VPWR _19981_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21480__A2 _21477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20206__A _20206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14055_ _14055_/A _14055_/B _14055_/C VGND VGND VPWR VPWR _14072_/B sky130_fd_sc_hd__and3_4
X_18932_ _18927_/A _18926_/X _18928_/Y _18931_/X VGND VGND VPWR VPWR _18932_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11828__A _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19103__A1_N _18971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13006_ _12886_/A _13075_/B VGND VGND VPWR VPWR _13006_/X sky130_fd_sc_hd__or2_4
XANTENNA__17436__A1 _15782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13170__A1 _12682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18863_ _15119_/X _18834_/A _24383_/Q _18835_/A VGND VGND VPWR VPWR _24383_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15019__B _23871_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17814_ _17826_/A VGND VGND VPWR VPWR _17814_/X sky130_fd_sc_hd__buf_2
XFILLER_67_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18794_ _15646_/X _18788_/X _20706_/A _18789_/X VGND VGND VPWR VPWR _24427_/D sky130_fd_sc_hd__o22a_4
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20991__A1 _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21037__A _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17745_ _17745_/A _17745_/B _17745_/C VGND VGND VPWR VPWR _17745_/X sky130_fd_sc_hd__or3_4
X_14957_ _13998_/A _14955_/X _14956_/X VGND VGND VPWR VPWR _14961_/B sky130_fd_sc_hd__and3_4
XANTENNA__12659__A _12963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15035__A _14748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13908_ _13908_/A _13904_/X _13907_/X VGND VGND VPWR VPWR _13908_/X sky130_fd_sc_hd__or3_4
XANTENNA__19730__A _19730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17676_ _17684_/A VGND VGND VPWR VPWR _17676_/Y sky130_fd_sc_hd__inv_2
X_14888_ _13983_/A _23872_/Q VGND VGND VPWR VPWR _14890_/B sky130_fd_sc_hd__or2_4
XANTENNA__21940__B1 _23538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_30_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19415_ _19430_/B VGND VGND VPWR VPWR _19416_/B sky130_fd_sc_hd__buf_2
XFILLER_51_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16627_ _16616_/A _16627_/B _16627_/C VGND VGND VPWR VPWR _16635_/B sky130_fd_sc_hd__and3_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13839_ _13839_/A VGND VGND VPWR VPWR _13847_/A sky130_fd_sc_hd__buf_2
XANTENNA__14874__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20595__B _20595_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19346_ _19343_/X _18572_/X _19343_/X _24231_/Q VGND VGND VPWR VPWR _24231_/D sky130_fd_sc_hd__a2bb2o_4
X_16558_ _16586_/A _16631_/B VGND VGND VPWR VPWR _16558_/X sky130_fd_sc_hd__or2_4
XANTENNA__22496__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15689__B _15689_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15509_ _15497_/A _15437_/B VGND VGND VPWR VPWR _15509_/X sky130_fd_sc_hd__or2_4
X_19277_ _19215_/B VGND VGND VPWR VPWR _19277_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12394__A _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16489_ _16464_/A _16489_/B VGND VGND VPWR VPWR _16489_/X sky130_fd_sc_hd__or2_4
X_18228_ _18129_/A VGND VGND VPWR VPWR _18228_/X sky130_fd_sc_hd__buf_2
XANTENNA__22248__B2 _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18159_ _17476_/C _18158_/X VGND VGND VPWR VPWR _18159_/X sky130_fd_sc_hd__or2_4
XFILLER_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21170_ _20315_/X _21169_/X _23965_/Q _21166_/X VGND VGND VPWR VPWR _21170_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21471__A2 _21470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20121_ _11565_/X _20119_/X _20120_/Y VGND VGND VPWR VPWR _20121_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__11738__A _11738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20052_ _20051_/X VGND VGND VPWR VPWR _20052_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23811_ _23494_/CLK _21442_/X VGND VGND VPWR VPWR _23811_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22184__B1 _23403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23742_ _23320_/CLK _21589_/X VGND VGND VPWR VPWR _23742_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20954_ _20283_/X _20945_/Y _20952_/X _20953_/Y _20459_/A VGND VGND VPWR VPWR _20955_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_96_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _23770_/CLK _23673_/D VGND VGND VPWR VPWR _16256_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _20732_/X _20884_/X _19113_/A _20739_/X VGND VGND VPWR VPWR _20886_/B sky130_fd_sc_hd__o22a_4
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22624_ _22394_/X _22622_/X _16654_/B _22619_/X VGND VGND VPWR VPWR _22624_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15599__B _23563_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22487__B2 _22483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24379__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22555_ _22446_/X _22550_/X _14275_/B _22554_/X VGND VGND VPWR VPWR _22555_/X sky130_fd_sc_hd__o22a_4
X_21506_ _21791_/A VGND VGND VPWR VPWR _21506_/X sky130_fd_sc_hd__buf_2
XANTENNA__22239__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22239__B2 _22233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22486_ _22486_/A VGND VGND VPWR VPWR _22486_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_35_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24225_ _24250_/CLK _19357_/X HRESETn VGND VGND VPWR VPWR _24225_/Q sky130_fd_sc_hd__dfrtp_4
X_21437_ _21416_/A VGND VGND VPWR VPWR _21437_/X sky130_fd_sc_hd__buf_2
XANTENNA__21998__B1 _15455_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12170_ _11827_/A _23709_/Q VGND VGND VPWR VPWR _12172_/B sky130_fd_sc_hd__or2_4
X_24156_ _24293_/CLK _24156_/D HRESETn VGND VGND VPWR VPWR _24156_/Q sky130_fd_sc_hd__dfrtp_4
X_21368_ _21244_/X _21362_/X _23860_/Q _21366_/X VGND VGND VPWR VPWR _21368_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23107_ _23107_/CLK _23107_/D VGND VGND VPWR VPWR _14762_/B sky130_fd_sc_hd__dfxtp_4
X_20319_ _20492_/A VGND VGND VPWR VPWR _20319_/X sky130_fd_sc_hd__buf_2
X_24087_ _24088_/CLK _24087_/D VGND VGND VPWR VPWR _24087_/Q sky130_fd_sc_hd__dfxtp_4
X_21299_ _21299_/A VGND VGND VPWR VPWR _21300_/A sky130_fd_sc_hd__buf_2
XANTENNA__14024__A _12598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23038_ _18000_/X _23038_/B VGND VGND VPWR VPWR _23039_/C sky130_fd_sc_hd__or2_4
XANTENNA__18615__B1 _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13863__A _13879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15860_ _13546_/X _15805_/B VGND VGND VPWR VPWR _15862_/B sky130_fd_sc_hd__or2_4
XFILLER_49_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14811_ _14811_/A _14811_/B VGND VGND VPWR VPWR _14811_/X sky130_fd_sc_hd__or2_4
XFILLER_76_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15791_ _12443_/A _15852_/B VGND VGND VPWR VPWR _15791_/X sky130_fd_sc_hd__or2_4
XANTENNA__12479__A _12466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18918__A1 _15249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17530_ _17530_/A VGND VGND VPWR VPWR _17530_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19550__A HRDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11954_ _11954_/A VGND VGND VPWR VPWR _11955_/A sky130_fd_sc_hd__buf_2
X_14742_ _15413_/A _14742_/B VGND VGND VPWR VPWR _14744_/B sky130_fd_sc_hd__or2_4
XFILLER_79_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20725__A1 _20613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20725__B2 _20724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20696__A _20696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14673_ _14673_/A _14671_/X _14673_/C VGND VGND VPWR VPWR _14678_/B sky130_fd_sc_hd__and3_4
X_17461_ _17156_/Y _17461_/B VGND VGND VPWR VPWR _17461_/X sky130_fd_sc_hd__or2_4
XFILLER_72_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11885_ _11884_/X VGND VGND VPWR VPWR _16286_/A sky130_fd_sc_hd__buf_2
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19200_ _24288_/Q _19108_/X _19199_/Y VGND VGND VPWR VPWR _19200_/X sky130_fd_sc_hd__o21a_4
XFILLER_18_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13624_ _13624_/A _13624_/B _13624_/C VGND VGND VPWR VPWR _13625_/C sky130_fd_sc_hd__and3_4
X_16412_ _11852_/X _16386_/X _16393_/X _16403_/X _16411_/X VGND VGND VPWR VPWR _16412_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_38_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23906__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_117_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR _23316_/CLK sky130_fd_sc_hd__clkbuf_1
X_17392_ _17262_/A VGND VGND VPWR VPWR _18760_/C sky130_fd_sc_hd__inv_2
XFILLER_38_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19131_ _24310_/Q _19157_/A VGND VGND VPWR VPWR _19132_/B sky130_fd_sc_hd__and2_4
XFILLER_73_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13555_ _13500_/X _13555_/B _13555_/C VGND VGND VPWR VPWR _13556_/C sky130_fd_sc_hd__and3_4
X_16343_ _16364_/A _23609_/Q VGND VGND VPWR VPWR _16345_/B sky130_fd_sc_hd__or2_4
XANTENNA__21150__B2 _21144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12506_ _12920_/A _12506_/B _12506_/C VGND VGND VPWR VPWR _12515_/B sky130_fd_sc_hd__and3_4
XANTENNA__13103__A _12957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16274_ _16151_/A _16272_/X _16273_/X VGND VGND VPWR VPWR _16274_/X sky130_fd_sc_hd__and3_4
X_19062_ _19062_/A VGND VGND VPWR VPWR _19062_/Y sky130_fd_sc_hd__inv_2
X_13486_ _12466_/X _13486_/B _13485_/X VGND VGND VPWR VPWR _13486_/X sky130_fd_sc_hd__and3_4
XANTENNA__22416__A _22416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15225_ _14225_/A _15225_/B VGND VGND VPWR VPWR _15227_/B sky130_fd_sc_hd__or2_4
X_18013_ _18012_/X _18013_/B VGND VGND VPWR VPWR _18014_/B sky130_fd_sc_hd__or2_4
X_12437_ _15013_/A VGND VGND VPWR VPWR _13925_/A sky130_fd_sc_hd__buf_2
XANTENNA__17106__B1 _13594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16414__A _16002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15156_ _11954_/A _15156_/B VGND VGND VPWR VPWR _15156_/X sky130_fd_sc_hd__or2_4
X_12368_ _12360_/A _12270_/B VGND VGND VPWR VPWR _12368_/X sky130_fd_sc_hd__or2_4
XFILLER_47_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14107_ _14318_/A _23977_/Q VGND VGND VPWR VPWR _14108_/C sky130_fd_sc_hd__or2_4
XANTENNA__21014__A2_N _21013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15087_ _12341_/A _23871_/Q VGND VGND VPWR VPWR _15087_/X sky130_fd_sc_hd__or2_4
X_19964_ _18653_/X _16937_/X _19934_/X _19963_/X VGND VGND VPWR VPWR _19964_/X sky130_fd_sc_hd__o22a_4
XFILLER_4_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12299_ _12255_/X _12297_/X _12298_/X VGND VGND VPWR VPWR _12299_/X sky130_fd_sc_hd__and3_4
XANTENNA__18756__A2_N _18755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14038_ _14055_/A _14038_/B _14038_/C VGND VGND VPWR VPWR _14039_/C sky130_fd_sc_hd__and3_4
X_18915_ _17297_/X _18912_/X _19083_/A _18913_/X VGND VGND VPWR VPWR _24356_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21205__A2 _21204_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19895_ _19884_/X _20875_/A _19894_/X VGND VGND VPWR VPWR _24158_/D sky130_fd_sc_hd__o21ai_4
XFILLER_68_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13773__A _13685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18846_ _17191_/X _18841_/X _24396_/Q _18842_/X VGND VGND VPWR VPWR _18846_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18777_ _17164_/X _18774_/X _24440_/Q _18775_/X VGND VGND VPWR VPWR _24440_/D sky130_fd_sc_hd__o22a_4
X_15989_ _15997_/A VGND VGND VPWR VPWR _16097_/A sky130_fd_sc_hd__buf_2
XFILLER_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18909__A1 _17178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12389__A _15889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22166__B1 _23416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22705__A2 _22700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17728_ _17726_/X _17300_/X VGND VGND VPWR VPWR _17732_/B sky130_fd_sc_hd__and2_4
XANTENNA__19460__A _19433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20716__A1 _18475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17659_ _17659_/A _17658_/Y VGND VGND VPWR VPWR _17659_/X sky130_fd_sc_hd__or2_4
XFILLER_23_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20670_ _20670_/A VGND VGND VPWR VPWR _21831_/A sky130_fd_sc_hd__buf_2
XFILLER_51_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12836__B _12836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19329_ _19325_/X _18258_/X _19328_/X _24243_/Q VGND VGND VPWR VPWR _24243_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21141__B2 _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13013__A _13032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22340_ _22354_/A VGND VGND VPWR VPWR _22340_/X sky130_fd_sc_hd__buf_2
XANTENNA__21692__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21230__A _21230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22271_ _22098_/X _22265_/X _12767_/B _22269_/X VGND VGND VPWR VPWR _22271_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12852__A _12852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16324__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24010_ _24011_/CLK _24010_/D VGND VGND VPWR VPWR _24010_/Q sky130_fd_sc_hd__dfxtp_4
X_21222_ _21271_/A VGND VGND VPWR VPWR _21247_/A sky130_fd_sc_hd__buf_2
XANTENNA__21444__A2 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22641__B2 _22640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12571__B _12571_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21153_ _20870_/X _21147_/X _14447_/B _21151_/X VGND VGND VPWR VPWR _21153_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15123__A2 _15119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20104_ _20097_/Y _20101_/Y _11572_/X _20103_/X VGND VGND VPWR VPWR _20104_/X sky130_fd_sc_hd__a211o_4
X_21084_ _20553_/X _21082_/X _24018_/Q _21079_/X VGND VGND VPWR VPWR _21084_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14779__A _13966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20035_ _18411_/X _20033_/X _20034_/Y _20020_/X VGND VGND VPWR VPWR _20035_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12893__B1 _12876_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22996__A _22995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12299__A _12255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16994__A _24190_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19370__A _19370_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21986_ _21811_/X _21981_/X _12571_/B _21985_/X VGND VGND VPWR VPWR _21986_/X sky130_fd_sc_hd__o22a_4
XFILLER_76_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _23922_/CLK _21614_/X VGND VGND VPWR VPWR _15849_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21405__A _21419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ _21287_/A VGND VGND VPWR VPWR _20937_/X sky130_fd_sc_hd__buf_2
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__A _13025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15403__A _13623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11670_/A VGND VGND VPWR VPWR _11671_/A sky130_fd_sc_hd__buf_2
X_23656_ _23304_/CLK _21721_/X VGND VGND VPWR VPWR _13627_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _24197_/Q _20751_/X _20867_/X VGND VGND VPWR VPWR _22134_/A sky130_fd_sc_hd__o21a_4
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12746__B _23860_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22607_ _22600_/A VGND VGND VPWR VPWR _22607_/X sky130_fd_sc_hd__buf_2
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23587_ _23270_/CLK _23587_/D VGND VGND VPWR VPWR _14758_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20799_ HRDATA[8] _20753_/B VGND VGND VPWR VPWR _20799_/X sky130_fd_sc_hd__or2_4
XANTENNA__14019__A _14071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21132__B2 _21130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13340_ _12738_/A _13340_/B VGND VGND VPWR VPWR _13342_/B sky130_fd_sc_hd__or2_4
X_22538_ _22418_/X _22536_/X _13005_/B _22533_/X VGND VGND VPWR VPWR _22538_/X sky130_fd_sc_hd__o22a_4
XFILLER_13_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22880__A1 _12031_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22236__A _22207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21140__A _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20891__B1 _20890_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13271_ _13270_/X VGND VGND VPWR VPWR _13272_/B sky130_fd_sc_hd__inv_2
X_22469_ _22476_/A VGND VGND VPWR VPWR _22469_/X sky130_fd_sc_hd__buf_2
XANTENNA__16234__A _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15010_ _15010_/A _23903_/Q VGND VGND VPWR VPWR _15012_/B sky130_fd_sc_hd__or2_4
X_12222_ _12221_/X _12222_/B VGND VGND VPWR VPWR _12222_/X sky130_fd_sc_hd__or2_4
X_24208_ _24208_/CLK _19390_/X HRESETn VGND VGND VPWR VPWR _24208_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21435__A2 _21433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12153_ _12153_/A _23965_/Q VGND VGND VPWR VPWR _12154_/C sky130_fd_sc_hd__or2_4
X_24139_ _24229_/CLK _19965_/Y HRESETn VGND VGND VPWR VPWR _24139_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19545__A _19545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12084_ _12091_/A _23965_/Q VGND VGND VPWR VPWR _12085_/C sky130_fd_sc_hd__or2_4
X_16961_ _22907_/B VGND VGND VPWR VPWR _17726_/A sky130_fd_sc_hd__inv_2
XANTENNA__15792__B _15792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21199__A1 _20797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21199__B2 _21194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18700_ _18487_/X _18692_/X _18693_/Y _18695_/X _18699_/Y VGND VGND VPWR VPWR _18700_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_46_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15912_ _15910_/Y _15911_/X VGND VGND VPWR VPWR _15913_/B sky130_fd_sc_hd__or2_4
X_19680_ HRDATA[23] VGND VGND VPWR VPWR _20445_/B sky130_fd_sc_hd__buf_2
X_16892_ _17052_/A VGND VGND VPWR VPWR _16916_/A sky130_fd_sc_hd__buf_2
XANTENNA__20946__B2 _20449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18631_ _17858_/X _18656_/B _18629_/Y _18424_/X _18630_/Y VGND VGND VPWR VPWR _18633_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15843_ _12716_/X _15820_/X _15827_/X _15834_/X _15842_/X VGND VGND VPWR VPWR _15843_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22148__B1 _23423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18562_ _17422_/A _18561_/X VGND VGND VPWR VPWR _18562_/X sky130_fd_sc_hd__or2_4
XANTENNA__22389__A2_N _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12986_ _12948_/A _12982_/X _12985_/X VGND VGND VPWR VPWR _12987_/C sky130_fd_sc_hd__or3_4
X_15774_ _15774_/A _15772_/X _15773_/X VGND VGND VPWR VPWR _15774_/X sky130_fd_sc_hd__and3_4
XANTENNA__22699__B2 _22697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17513_ _17513_/A _18332_/A _18281_/A _18307_/A VGND VGND VPWR VPWR _17514_/B sky130_fd_sc_hd__or4_4
XFILLER_79_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14725_ _14725_/A _14787_/B VGND VGND VPWR VPWR _14725_/X sky130_fd_sc_hd__or2_4
XFILLER_75_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11937_ _11936_/X VGND VGND VPWR VPWR _11999_/A sky130_fd_sc_hd__buf_2
X_18493_ _18142_/A _17416_/A _18489_/X _18398_/X _18492_/Y VGND VGND VPWR VPWR _18493_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12937__A _12937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16409__A _13442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21371__B2 _21366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11841__A _11841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15313__A _13839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17444_ _12992_/X _17524_/B VGND VGND VPWR VPWR _17444_/X sky130_fd_sc_hd__or2_4
X_11868_ _13654_/A VGND VGND VPWR VPWR _13624_/A sky130_fd_sc_hd__buf_2
X_14656_ _15108_/A _14656_/B _14655_/X VGND VGND VPWR VPWR _14656_/X sky130_fd_sc_hd__or3_4
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13607_ _15399_/A _13696_/B VGND VGND VPWR VPWR _13607_/X sky130_fd_sc_hd__or2_4
XANTENNA__11560__B IRQ[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17375_ _17363_/A _17374_/X VGND VGND VPWR VPWR _17375_/X sky130_fd_sc_hd__or2_4
XFILLER_18_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11799_ _11799_/A VGND VGND VPWR VPWR _12392_/A sky130_fd_sc_hd__buf_2
X_14587_ _14146_/X _14581_/X _14586_/X VGND VGND VPWR VPWR _14587_/X sky130_fd_sc_hd__or3_4
X_19114_ _19114_/A _19113_/X VGND VGND VPWR VPWR _19115_/B sky130_fd_sc_hd__and2_4
XANTENNA__24188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24362__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16326_ _16364_/A _16266_/B VGND VGND VPWR VPWR _16329_/B sky130_fd_sc_hd__or2_4
X_13538_ _11665_/X _13538_/B _13538_/C VGND VGND VPWR VPWR _13574_/B sky130_fd_sc_hd__or3_4
XANTENNA__22871__A1 _17272_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21674__A2 _21669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15967__B _15967_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19045_ _19024_/X _19043_/X _19044_/Y _19027_/X VGND VGND VPWR VPWR _19045_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13768__A _15491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13469_ _13437_/X _13547_/B VGND VGND VPWR VPWR _13469_/X sky130_fd_sc_hd__or2_4
X_16257_ _16252_/X _23993_/Q VGND VGND VPWR VPWR _16257_/X sky130_fd_sc_hd__or2_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12672__A _12672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24234__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15208_ _15201_/A _23649_/Q VGND VGND VPWR VPWR _15208_/X sky130_fd_sc_hd__or2_4
XANTENNA__21985__A _21985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16188_ _16188_/A VGND VGND VPWR VPWR _16227_/A sky130_fd_sc_hd__buf_2
XANTENNA__22623__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15139_ _14138_/X _23649_/Q VGND VGND VPWR VPWR _15139_/X sky130_fd_sc_hd__or2_4
XFILLER_5_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19947_ _17961_/X _18726_/Y _17856_/X _19946_/Y VGND VGND VPWR VPWR _19947_/X sky130_fd_sc_hd__a211o_4
XANTENNA__14599__A _14151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19878_ _19678_/A _19876_/X _19877_/X _16919_/Y _19531_/A VGND VGND VPWR VPWR _19878_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_60_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18829_ _16374_/X _18827_/X _24409_/Q _18828_/X VGND VGND VPWR VPWR _18829_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21840_ _21555_/A VGND VGND VPWR VPWR _21840_/X sky130_fd_sc_hd__buf_2
XANTENNA__13008__A _12915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19555__A1 _20342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21225__A _21795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21771_ _21558_/X _21769_/X _13767_/B _21766_/X VGND VGND VPWR VPWR _23624_/D sky130_fd_sc_hd__o22a_4
XFILLER_64_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12847__A _12443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20165__A2 IRQ[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23510_ _23539_/CLK _21984_/X VGND VGND VPWR VPWR _12213_/B sky130_fd_sc_hd__dfxtp_4
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11751__A _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20722_ _20722_/A VGND VGND VPWR VPWR _21265_/A sky130_fd_sc_hd__buf_2
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15223__A _14215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19307__A1 _18864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19307__B2 _19306_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23441_ _23889_/CLK _23441_/D VGND VGND VPWR VPWR _13166_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20653_ _20424_/A VGND VGND VPWR VPWR _20653_/X sky130_fd_sc_hd__buf_2
XFILLER_56_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_100_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR _23354_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23372_ _23404_/CLK _22232_/X VGND VGND VPWR VPWR _15432_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21665__A2 _21662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20584_ _20630_/A _20584_/B VGND VGND VPWR VPWR _20584_/Y sky130_fd_sc_hd__nor2_4
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15877__B _15815_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18190__A1_N _18425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22056__A _22035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22323_ _13794_/B VGND VGND VPWR VPWR _23303_/D sky130_fd_sc_hd__buf_2
XFILLER_118_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22254_ _22269_/A VGND VGND VPWR VPWR _22262_/A sky130_fd_sc_hd__buf_2
XANTENNA__21417__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21205_ _20893_/X _21204_/X _14689_/B _21201_/X VGND VGND VPWR VPWR _23940_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15893__A _13529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22185_ _22122_/X _22179_/X _13970_/B _22183_/X VGND VGND VPWR VPWR _22185_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19491__B1 _18864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22090__A2 _22089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21136_ _20574_/X _21133_/X _23985_/Q _21130_/X VGND VGND VPWR VPWR _21136_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21067_ _21067_/A VGND VGND VPWR VPWR _21075_/A sky130_fd_sc_hd__buf_2
XFILLER_115_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14302__A _12260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20928__B2 _20453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20018_ _19994_/A VGND VGND VPWR VPWR _20018_/X sky130_fd_sc_hd__buf_2
XFILLER_74_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12840_ _11800_/X _12840_/B _12839_/X VGND VGND VPWR VPWR _12841_/C sky130_fd_sc_hd__or3_4
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19546__A1 _20317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14956__B _14889_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19546__B2 HRDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12771_ _12948_/A VGND VGND VPWR VPWR _12771_/X sky130_fd_sc_hd__buf_2
X_21969_ _22002_/A VGND VGND VPWR VPWR _21985_/A sky130_fd_sc_hd__inv_2
XFILLER_76_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12757__A _13129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16229__A _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11661__A _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21353__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _13998_/A VGND VGND VPWR VPWR _11723_/A sky130_fd_sc_hd__buf_2
X_14510_ _13895_/A VGND VGND VPWR VPWR _14536_/A sky130_fd_sc_hd__buf_2
XFILLER_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15497_/A _15490_/B VGND VGND VPWR VPWR _15491_/C sky130_fd_sc_hd__or2_4
X_23708_ _23867_/CLK _23708_/D VGND VGND VPWR VPWR _23708_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11652_/X VGND VGND VPWR VPWR _14073_/A sky130_fd_sc_hd__buf_2
X_14441_ _14464_/A _14441_/B _14441_/C VGND VGND VPWR VPWR _14441_/X sky130_fd_sc_hd__and3_4
X_23639_ _23316_/CLK _23639_/D VGND VGND VPWR VPWR _23639_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18444__A _18390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21105__B2 _21100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19849__A2 _19845_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14372_ _13847_/A VGND VGND VPWR VPWR _15601_/A sky130_fd_sc_hd__buf_2
X_17160_ _17160_/A VGND VGND VPWR VPWR _17160_/X sky130_fd_sc_hd__buf_2
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ _11584_/A VGND VGND VPWR VPWR _11585_/A sky130_fd_sc_hd__inv_2
XANTENNA__21656__A2 _21655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13323_ _13281_/X _13321_/X _13322_/X VGND VGND VPWR VPWR _13324_/C sky130_fd_sc_hd__and3_4
X_16111_ _16139_/A _23543_/Q VGND VGND VPWR VPWR _16111_/X sky130_fd_sc_hd__or2_4
XFILLER_7_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17091_ _17049_/B _17090_/X VGND VGND VPWR VPWR _17096_/C sky130_fd_sc_hd__nor2_4
XANTENNA__12492__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13254_ _13242_/A _13254_/B VGND VGND VPWR VPWR _13255_/C sky130_fd_sc_hd__or2_4
X_16042_ _16058_/A _16040_/X _16042_/C VGND VGND VPWR VPWR _16042_/X sky130_fd_sc_hd__and3_4
XFILLER_87_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22605__B2 _22604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12205_ _12496_/A VGND VGND VPWR VPWR _12553_/A sky130_fd_sc_hd__buf_2
XFILLER_108_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13185_ _12738_/A _23473_/Q VGND VGND VPWR VPWR _13185_/X sky130_fd_sc_hd__or2_4
XFILLER_83_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19801_ _19742_/A _19775_/Y VGND VGND VPWR VPWR _19801_/X sky130_fd_sc_hd__or2_4
XANTENNA__20092__A1 _20076_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12136_ _12167_/A _23933_/Q VGND VGND VPWR VPWR _12136_/X sky130_fd_sc_hd__or2_4
XANTENNA__20092__B2 _18649_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17993_ _18085_/A _18083_/A _17572_/X VGND VGND VPWR VPWR _17993_/X sky130_fd_sc_hd__o21a_4
X_19732_ _19784_/B _19643_/B _19637_/Y _19857_/C VGND VGND VPWR VPWR _19732_/X sky130_fd_sc_hd__and4_4
XFILLER_81_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11836__A _16677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12067_ _12088_/A _12064_/X _12067_/C VGND VGND VPWR VPWR _12073_/B sky130_fd_sc_hd__and3_4
X_16944_ _24132_/Q VGND VGND VPWR VPWR _17661_/A sky130_fd_sc_hd__inv_2
XANTENNA__15308__A _14748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14212__A _14367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19663_ _19663_/A VGND VGND VPWR VPWR _19663_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15027__B _23807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16875_ _13590_/X _16874_/X _13590_/X _16874_/X VGND VGND VPWR VPWR _16876_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19722__B _19689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21592__B2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18614_ _17336_/B VGND VGND VPWR VPWR _18614_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15826_ _12522_/A _15826_/B _15826_/C VGND VGND VPWR VPWR _15827_/C sky130_fd_sc_hd__and3_4
XFILLER_24_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19594_ _19593_/X VGND VGND VPWR VPWR _19624_/A sky130_fd_sc_hd__buf_2
XFILLER_59_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14866__B _14866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18545_ _18697_/A _17598_/Y VGND VGND VPWR VPWR _18545_/X sky130_fd_sc_hd__and2_4
XFILLER_98_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15757_ _15750_/A _15757_/B VGND VGND VPWR VPWR _15759_/B sky130_fd_sc_hd__or2_4
XFILLER_80_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12969_ _12981_/A _23411_/Q VGND VGND VPWR VPWR _12969_/X sky130_fd_sc_hd__or2_4
XFILLER_45_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16139__A _16139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21344__B2 _21301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22541__B1 _13291_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14708_ _15592_/A _14708_/B _14707_/X VGND VGND VPWR VPWR _14708_/X sky130_fd_sc_hd__and3_4
X_18476_ _18458_/X _18463_/Y _18357_/X _18475_/X VGND VGND VPWR VPWR _18476_/X sky130_fd_sc_hd__o22a_4
XFILLER_94_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21895__A2 _21894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15688_ _15688_/A _15688_/B _15687_/X VGND VGND VPWR VPWR _15688_/X sky130_fd_sc_hd__or3_4
XFILLER_21_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17427_ _14263_/X _17427_/B VGND VGND VPWR VPWR _17427_/X sky130_fd_sc_hd__or2_4
X_14639_ _12267_/X _14613_/X _14622_/X _14630_/X _14638_/X VGND VGND VPWR VPWR _14639_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_53_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17358_ _17356_/B VGND VGND VPWR VPWR _17432_/B sky130_fd_sc_hd__inv_2
XFILLER_105_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22844__A1 _17298_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21647__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15697__B _15697_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23624__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16309_ _16322_/A _16244_/B VGND VGND VPWR VPWR _16309_/X sky130_fd_sc_hd__or2_4
XANTENNA__13498__A _15884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17289_ _17543_/A VGND VGND VPWR VPWR _17290_/A sky130_fd_sc_hd__inv_2
XFILLER_101_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19028_ _19024_/X _19025_/Y _19026_/Y _19027_/X VGND VGND VPWR VPWR _19028_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22604__A _22583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20607__B1 _20606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19473__B1 HRDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23990_ _24084_/CLK _23990_/D VGND VGND VPWR VPWR _12248_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_69_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14122__A _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_25_0_HCLK clkbuf_7_25_0_HCLK/A VGND VGND VPWR VPWR _23104_/CLK sky130_fd_sc_hd__clkbuf_1
X_22941_ _22952_/A _22939_/Y _22941_/C VGND VGND VPWR VPWR _22941_/X sky130_fd_sc_hd__and3_4
XFILLER_112_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_88_0_HCLK clkbuf_6_44_0_HCLK/X VGND VGND VPWR VPWR _24059_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_56_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13961__A _13611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22872_ _22872_/A _22872_/B VGND VGND VPWR VPWR HWDATA[28] sky130_fd_sc_hd__nor2_4
XANTENNA__20791__C1 _20790_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21823_ _20591_/A VGND VGND VPWR VPWR _21823_/X sky130_fd_sc_hd__buf_2
XFILLER_71_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12577__A _12638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21335__A1 _21273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21335__B2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22532__B1 _12228_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21754_ _21529_/X _21748_/X _12836_/B _21752_/X VGND VGND VPWR VPWR _21754_/X sky130_fd_sc_hd__o22a_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20705_ _24395_/Q _20595_/B VGND VGND VPWR VPWR _20705_/Y sky130_fd_sc_hd__nand2_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24473_ _24473_/CLK _24473_/D HRESETn VGND VGND VPWR VPWR _19981_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15888__A _13522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21685_ _21684_/X VGND VGND VPWR VPWR _21690_/A sky130_fd_sc_hd__buf_2
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14792__A _12575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23424_ _23104_/CLK _22146_/X VGND VGND VPWR VPWR _14883_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20636_ _22112_/A VGND VGND VPWR VPWR _21543_/A sky130_fd_sc_hd__buf_2
XANTENNA__22835__A1 _17115_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23355_ _23293_/CLK _22261_/X VGND VGND VPWR VPWR _16749_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15400__B _15463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20567_ _18309_/X _20424_/X _20516_/X _20566_/Y VGND VGND VPWR VPWR _20568_/A sky130_fd_sc_hd__a211o_4
X_22306_ _15960_/B VGND VGND VPWR VPWR _23320_/D sky130_fd_sc_hd__buf_2
XFILLER_10_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23286_ _23473_/CLK _23286_/D VGND VGND VPWR VPWR _12241_/B sky130_fd_sc_hd__dfxtp_4
X_20498_ _20403_/X _20496_/X _19225_/A _20497_/X VGND VGND VPWR VPWR _20498_/X sky130_fd_sc_hd__o22a_4
XFILLER_106_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22599__B1 _14025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22237_ _22124_/X _22236_/X _23369_/Q _22233_/X VGND VGND VPWR VPWR _23369_/D sky130_fd_sc_hd__o22a_4
XFILLER_30_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22063__A2 _22059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16512__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22168_ _22093_/X _22165_/X _12298_/B _22162_/X VGND VGND VPWR VPWR _22168_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21810__A2 _21805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18019__A1 _18011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21119_ _21133_/A VGND VGND VPWR VPWR _21119_/X sky130_fd_sc_hd__buf_2
XFILLER_47_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11656__A _11656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14990_ _14990_/A _23487_/Q VGND VGND VPWR VPWR _14991_/C sky130_fd_sc_hd__or2_4
X_22099_ _22098_/X _22089_/X _12711_/B _22096_/X VGND VGND VPWR VPWR _23444_/D sky130_fd_sc_hd__o22a_4
XFILLER_47_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19767__A1 _19429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13941_ _12302_/A _13937_/X _13941_/C VGND VGND VPWR VPWR _13941_/X sky130_fd_sc_hd__or3_4
XFILLER_59_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20377__A2 _20754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16660_ _16599_/X _16660_/B _16659_/X VGND VGND VPWR VPWR _16660_/X sky130_fd_sc_hd__or3_4
XANTENNA__23064__B _23064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13872_ _13872_/A VGND VGND VPWR VPWR _13909_/A sky130_fd_sc_hd__buf_2
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15611_ _15611_/A _15611_/B _15611_/C VGND VGND VPWR VPWR _15612_/C sky130_fd_sc_hd__or3_4
X_12823_ _12799_/A _12823_/B VGND VGND VPWR VPWR _12825_/B sky130_fd_sc_hd__or2_4
X_16591_ _12025_/A _16591_/B _16590_/X VGND VGND VPWR VPWR _16592_/C sky130_fd_sc_hd__and3_4
XFILLER_90_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12487__A _13022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18330_ _18330_/A VGND VGND VPWR VPWR _18330_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15542_ _12533_/A _15538_/X _15541_/X VGND VGND VPWR VPWR _15542_/X sky130_fd_sc_hd__or3_4
X_12754_ _12947_/A VGND VGND VPWR VPWR _12754_/X sky130_fd_sc_hd__buf_2
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11803_/A _11705_/B VGND VGND VPWR VPWR _11705_/X sky130_fd_sc_hd__or2_4
X_18261_ _17672_/A _16980_/B _16981_/B VGND VGND VPWR VPWR _22992_/B sky130_fd_sc_hd__a21bo_4
XFILLER_43_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15798__A _12462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _15654_/A _12685_/B _12685_/C VGND VGND VPWR VPWR _12689_/B sky130_fd_sc_hd__and3_4
X_15473_ _15480_/A _15473_/B VGND VGND VPWR VPWR _15473_/X sky130_fd_sc_hd__or2_4
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17182_/Y _17155_/X _14263_/X _17186_/X VGND VGND VPWR VPWR _17212_/X sky130_fd_sc_hd__o22a_4
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ _19927_/A VGND VGND VPWR VPWR _16891_/A sky130_fd_sc_hd__inv_2
X_14424_ _14423_/X VGND VGND VPWR VPWR _14425_/A sky130_fd_sc_hd__buf_2
XFILLER_50_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18192_ _18191_/A _18190_/X _18048_/X VGND VGND VPWR VPWR _18192_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21629__A2 _21626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20209__A _20444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17143_ _14852_/Y VGND VGND VPWR VPWR _17143_/X sky130_fd_sc_hd__buf_2
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11567_ _24442_/Q IRQ[27] _11566_/X VGND VGND VPWR VPWR _11567_/X sky130_fd_sc_hd__a21o_4
X_14355_ _15614_/A _14275_/B VGND VGND VPWR VPWR _14355_/X sky130_fd_sc_hd__or2_4
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14207__A _14207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13111__A _13104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13306_ _13303_/X _13304_/X _13305_/X VGND VGND VPWR VPWR _13306_/X sky130_fd_sc_hd__and3_4
X_14286_ _15543_/A VGND VGND VPWR VPWR _15536_/A sky130_fd_sc_hd__buf_2
X_17074_ _17224_/A _17073_/X VGND VGND VPWR VPWR _18498_/A sky130_fd_sc_hd__or2_4
XFILLER_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13237_ _11664_/A _13237_/B _13237_/C VGND VGND VPWR VPWR _13237_/X sky130_fd_sc_hd__or3_4
X_16025_ _16025_/A VGND VGND VPWR VPWR _16050_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22054__A2 _22052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19455__B1 _20224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13168_ _12713_/A _13164_/X _13167_/X VGND VGND VPWR VPWR _13168_/X sky130_fd_sc_hd__or3_4
XANTENNA__21801__A2 _21793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16141__B _16226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12119_ _16072_/A VGND VGND VPWR VPWR _12153_/A sky130_fd_sc_hd__buf_2
XANTENNA__15038__A _14778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13099_ _13115_/A _23538_/Q VGND VGND VPWR VPWR _13100_/C sky130_fd_sc_hd__or2_4
X_17976_ _17911_/X _17831_/X _17807_/X _17827_/X VGND VGND VPWR VPWR _17976_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19715_ _19876_/B _19663_/A _19692_/X VGND VGND VPWR VPWR _19715_/Y sky130_fd_sc_hd__a21oi_4
X_16927_ _16927_/A VGND VGND VPWR VPWR _16927_/X sky130_fd_sc_hd__buf_2
XFILLER_22_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19646_ _19629_/A _19645_/A _19629_/B VGND VGND VPWR VPWR _19646_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16858_ _15386_/X _14855_/Y _16857_/Y _14855_/A VGND VGND VPWR VPWR _16858_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15809_ _12886_/A _15864_/B VGND VGND VPWR VPWR _15810_/C sky130_fd_sc_hd__or2_4
XFILLER_65_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19577_ _19639_/A VGND VGND VPWR VPWR _19722_/A sky130_fd_sc_hd__buf_2
XFILLER_94_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16789_ _16773_/A _23835_/Q VGND VGND VPWR VPWR _16790_/C sky130_fd_sc_hd__or2_4
XFILLER_59_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21317__B2 _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18528_ _18486_/X _18520_/Y _18521_/X _18523_/X _18527_/Y VGND VGND VPWR VPWR _18528_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24132__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21503__A _21515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18459_ _18459_/A _18350_/B VGND VGND VPWR VPWR _18459_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__17941__B1 _17874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21470_ _21470_/A VGND VGND VPWR VPWR _21470_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20421_ _20421_/A VGND VGND VPWR VPWR _20421_/X sky130_fd_sc_hd__buf_2
XANTENNA__18812__A _11599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23140_ _23433_/CLK _23140_/D VGND VGND VPWR VPWR _14674_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13021__A _12494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20352_ _20209_/X _20343_/Y _20350_/X _20351_/Y _20233_/X VGND VGND VPWR VPWR _20353_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23071_ _23487_/CLK _23071_/D VGND VGND VPWR VPWR _23071_/Q sky130_fd_sc_hd__dfxtp_4
X_20283_ _20421_/A VGND VGND VPWR VPWR _20283_/X sky130_fd_sc_hd__buf_2
XANTENNA__12860__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22022_ _22016_/Y _22021_/X _21789_/X _22021_/X VGND VGND VPWR VPWR _22022_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19997__A1 _18169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19749__A1 _19554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23973_ _23973_/CLK _21153_/X VGND VGND VPWR VPWR _14447_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14787__A _13872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22924_ _22924_/A VGND VGND VPWR VPWR _22924_/X sky130_fd_sc_hd__buf_2
XFILLER_112_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22855_ _22855_/A VGND VGND VPWR VPWR _22855_/X sky130_fd_sc_hd__buf_2
XANTENNA__21308__A1 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21308__B2 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21806_ _21804_/X _21805_/X _23608_/Q _21800_/X VGND VGND VPWR VPWR _23608_/D sky130_fd_sc_hd__o22a_4
X_22786_ _17109_/Y _22782_/X VGND VGND VPWR VPWR HWDATA[3] sky130_fd_sc_hd__nor2_4
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12100__A _16541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21737_ _21752_/A VGND VGND VPWR VPWR _21737_/X sky130_fd_sc_hd__buf_2
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19921__B2 _20939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15411__A _15411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12470_ _12868_/A _24021_/Q VGND VGND VPWR VPWR _12479_/B sky130_fd_sc_hd__or2_4
XANTENNA__22808__A1 _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21668_ _21553_/X _21662_/X _23690_/Q _21666_/X VGND VGND VPWR VPWR _21668_/X sky130_fd_sc_hd__o22a_4
X_24456_ _24203_/CLK _24456_/D HRESETn VGND VGND VPWR VPWR _24456_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16226__B _16226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20619_ _20802_/A VGND VGND VPWR VPWR _20619_/X sky130_fd_sc_hd__buf_2
X_23407_ _23311_/CLK _22178_/X VGND VGND VPWR VPWR _13554_/B sky130_fd_sc_hd__dfxtp_4
X_24387_ _24425_/CLK _18859_/X HRESETn VGND VGND VPWR VPWR _24387_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22284__A2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21599_ _21519_/X _21598_/X _23736_/Q _21595_/X VGND VGND VPWR VPWR _23736_/D sky130_fd_sc_hd__o22a_4
X_14140_ _14318_/A _23817_/Q VGND VGND VPWR VPWR _14141_/C sky130_fd_sc_hd__or2_4
X_23338_ _24011_/CLK _22285_/X VGND VGND VPWR VPWR _23338_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14071_ _14071_/A _14062_/X _14070_/X VGND VGND VPWR VPWR _14072_/C sky130_fd_sc_hd__and3_4
XANTENNA__13866__A _11670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23269_ _23365_/CLK _22374_/X VGND VGND VPWR VPWR _14511_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12770__A _12753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16242__A _16147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13022_ _13022_/A _13089_/B VGND VGND VPWR VPWR _13024_/B sky130_fd_sc_hd__or2_4
XFILLER_112_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17999__B1 _17998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17830_ _17826_/X _17188_/X _17804_/A _17205_/X VGND VGND VPWR VPWR _17830_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18660__A1 _18424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20699__A HRDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17761_ _17755_/X _17756_/Y _17669_/X _17760_/X VGND VGND VPWR VPWR _17761_/X sky130_fd_sc_hd__or4_4
X_14973_ _15072_/A _14912_/B VGND VGND VPWR VPWR _14975_/B sky130_fd_sc_hd__or2_4
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14697__A _15114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19500_ _19483_/X VGND VGND VPWR VPWR _19500_/X sky130_fd_sc_hd__buf_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21547__B2 _21539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16712_ _12036_/X _16689_/X _16696_/X _16703_/X _16711_/X VGND VGND VPWR VPWR _16712_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17073__A _18728_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13924_ _15047_/A VGND VGND VPWR VPWR _14172_/A sky130_fd_sc_hd__buf_2
X_17692_ _17692_/A VGND VGND VPWR VPWR _17692_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_71_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR _24330_/CLK sky130_fd_sc_hd__clkbuf_1
X_19431_ _19433_/A VGND VGND VPWR VPWR _19431_/X sky130_fd_sc_hd__buf_2
X_16643_ _16640_/X _16641_/X _16643_/C VGND VGND VPWR VPWR _16643_/X sky130_fd_sc_hd__and3_4
XFILLER_47_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13855_ _13710_/A VGND VGND VPWR VPWR _14499_/A sky130_fd_sc_hd__buf_2
XFILLER_95_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12806_ _12822_/A _12806_/B _12806_/C VGND VGND VPWR VPWR _12807_/C sky130_fd_sc_hd__and3_4
X_19362_ _19306_/Y _16992_/Y _24140_/Q _16992_/A VGND VGND VPWR VPWR _23056_/B sky130_fd_sc_hd__o22a_4
X_16574_ _16567_/A _16657_/B VGND VGND VPWR VPWR _16576_/B sky130_fd_sc_hd__or2_4
XANTENNA__12010__A _16536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13786_ _12450_/A _13784_/X _13785_/X VGND VGND VPWR VPWR _13786_/X sky130_fd_sc_hd__and3_4
X_18313_ _18291_/X _18312_/X _24465_/Q _18291_/X VGND VGND VPWR VPWR _18313_/X sky130_fd_sc_hd__a2bb2o_4
X_15525_ _15552_/A _23339_/Q VGND VGND VPWR VPWR _15525_/X sky130_fd_sc_hd__or2_4
XANTENNA__21323__A _21316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19912__B2 _20400_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12737_ _12737_/A _12735_/X _12737_/C VGND VGND VPWR VPWR _12737_/X sky130_fd_sc_hd__and3_4
X_19293_ _19207_/B VGND VGND VPWR VPWR _19293_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18244_ _18244_/A _18241_/Y _18244_/C _18243_/X VGND VGND VPWR VPWR _18245_/A sky130_fd_sc_hd__or4_4
XANTENNA__15321__A _11638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15456_ _15495_/A _15454_/X _15455_/X VGND VGND VPWR VPWR _15456_/X sky130_fd_sc_hd__and3_4
X_12668_ _12622_/X _12668_/B VGND VGND VPWR VPWR _12669_/C sky130_fd_sc_hd__or2_4
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _14379_/A _14328_/B VGND VGND VPWR VPWR _14407_/X sky130_fd_sc_hd__or2_4
XANTENNA__15040__B _23071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11619_ _11618_/X VGND VGND VPWR VPWR _11619_/X sky130_fd_sc_hd__buf_2
X_18175_ _18172_/Y _18174_/X _18172_/Y _18174_/X VGND VGND VPWR VPWR _19378_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22275__A2 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15387_ _15387_/A _15387_/B VGND VGND VPWR VPWR _15387_/X sky130_fd_sc_hd__and2_4
X_12599_ _12599_/A VGND VGND VPWR VPWR _12617_/A sky130_fd_sc_hd__buf_2
XFILLER_117_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17126_ _11634_/A _17036_/A _24165_/Q _15784_/A _17125_/Y VGND VGND VPWR VPWR _17126_/X
+ sky130_fd_sc_hd__a32o_4
X_14338_ _13686_/A VGND VGND VPWR VPWR _15589_/A sky130_fd_sc_hd__buf_2
XFILLER_102_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22154__A _22169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17057_ _17057_/A VGND VGND VPWR VPWR _17224_/A sky130_fd_sc_hd__inv_2
X_14269_ _12238_/X _14269_/B VGND VGND VPWR VPWR _14270_/C sky130_fd_sc_hd__or2_4
XFILLER_83_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16008_ _16007_/X VGND VGND VPWR VPWR _16008_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20105__C _19027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17959_ _17779_/X _17959_/B _17959_/C _17959_/D VGND VGND VPWR VPWR _17960_/A sky130_fd_sc_hd__or4_4
XFILLER_111_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23812__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18079__A _17871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24384__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20970_ _20970_/A VGND VGND VPWR VPWR _20970_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14400__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19629_ _19629_/A _19629_/B VGND VGND VPWR VPWR _19629_/X sky130_fd_sc_hd__and2_4
XFILLER_54_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22640_ _22633_/A VGND VGND VPWR VPWR _22640_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13016__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22571_ _22600_/A VGND VGND VPWR VPWR _22586_/A sky130_fd_sc_hd__buf_2
XFILLER_35_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12855__A _12458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21710__B2 _21709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21522_ _20442_/A VGND VGND VPWR VPWR _21522_/X sky130_fd_sc_hd__buf_2
X_24310_ _24301_/CLK _19156_/X HRESETn VGND VGND VPWR VPWR _24310_/Q sky130_fd_sc_hd__dfrtp_4
X_24241_ _24241_/CLK _19331_/X HRESETn VGND VGND VPWR VPWR _24241_/Q sky130_fd_sc_hd__dfrtp_4
X_21453_ _21452_/X VGND VGND VPWR VPWR _21453_/X sky130_fd_sc_hd__buf_2
XANTENNA__22266__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18542__A _18392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20404_ _18813_/X VGND VGND VPWR VPWR _20405_/A sky130_fd_sc_hd__buf_2
X_24172_ _24299_/CLK _19799_/Y HRESETn VGND VGND VPWR VPWR _17069_/A sky130_fd_sc_hd__dfrtp_4
X_21384_ _21270_/X _21383_/X _23849_/Q _21380_/X VGND VGND VPWR VPWR _23849_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17142__A1 _15381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23123_ _24082_/CLK _23123_/D VGND VGND VPWR VPWR _12965_/B sky130_fd_sc_hd__dfxtp_4
X_20335_ _20209_/X _20318_/Y _20333_/X _20334_/Y _20233_/X VGND VGND VPWR VPWR _20335_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13686__A _13686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18890__A1 _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22999__A _18256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23054_ _19925_/X _16937_/X _23026_/X _23053_/X VGND VGND VPWR VPWR _23055_/A sky130_fd_sc_hd__a211o_4
XFILLER_118_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20266_ _20525_/A VGND VGND VPWR VPWR _20518_/A sky130_fd_sc_hd__inv_2
XFILLER_116_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22005_ _21845_/X _22002_/X _23495_/Q _21999_/X VGND VGND VPWR VPWR _23495_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21777__B2 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24339__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20197_ _22017_/A _20197_/B _21212_/B VGND VGND VPWR VPWR _21866_/D sky130_fd_sc_hd__or3_4
XFILLER_76_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23492__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20312__A _20484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22726__B1 _23064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15406__A _13794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11934__A _11933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11970_ _11962_/X VGND VGND VPWR VPWR _11971_/A sky130_fd_sc_hd__buf_2
X_23956_ _24021_/CLK _21182_/X VGND VGND VPWR VPWR _23956_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_58_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22907_ _22899_/X _22907_/B VGND VGND VPWR VPWR _22911_/B sky130_fd_sc_hd__or2_4
XFILLER_5_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23887_ _23859_/CLK _21325_/X VGND VGND VPWR VPWR _23887_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13640_ _13659_/A _13723_/B VGND VGND VPWR VPWR _13640_/X sky130_fd_sc_hd__or2_4
X_22838_ _17109_/Y _22826_/X _22827_/X VGND VGND VPWR VPWR _22838_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22884__D _19888_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18158__B1 _18082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _12771_/X _13571_/B _13570_/X VGND VGND VPWR VPWR _13572_/C sky130_fd_sc_hd__or3_4
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22769_ _22741_/Y _22768_/A VGND VGND VPWR VPWR _22773_/B sky130_fd_sc_hd__or2_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12765__A _13097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21701__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15310_ _14172_/A _15309_/X VGND VGND VPWR VPWR _15310_/X sky130_fd_sc_hd__and2_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A _12519_/X _12522_/C VGND VGND VPWR VPWR _12528_/B sky130_fd_sc_hd__and3_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16290_ _15934_/X _16368_/B VGND VGND VPWR VPWR _16290_/X sky130_fd_sc_hd__or2_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20982__A _21291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15241_ _15234_/A _15241_/B VGND VGND VPWR VPWR _15241_/X sky130_fd_sc_hd__or2_4
X_12453_ _12850_/A VGND VGND VPWR VPWR _12462_/A sky130_fd_sc_hd__buf_2
X_24439_ _24277_/CLK _24439_/D HRESETn VGND VGND VPWR VPWR _20427_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12384_ _12958_/A VGND VGND VPWR VPWR _12384_/X sky130_fd_sc_hd__buf_2
X_15172_ _14725_/A _15243_/B VGND VGND VPWR VPWR _15172_/X sky130_fd_sc_hd__or2_4
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14123_ _14998_/A _14123_/B _14122_/X VGND VGND VPWR VPWR _14123_/X sky130_fd_sc_hd__and3_4
XFILLER_67_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19980_ _19979_/X VGND VGND VPWR VPWR _19980_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18881__A1 _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18931_ _18931_/A _20268_/A VGND VGND VPWR VPWR _18931_/X sky130_fd_sc_hd__and2_4
XFILLER_119_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14054_ _14037_/A _14050_/X _14054_/C VGND VGND VPWR VPWR _14055_/C sky130_fd_sc_hd__or3_4
XFILLER_79_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21768__B2 _21766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13005_ _12879_/A _13005_/B VGND VGND VPWR VPWR _13005_/X sky130_fd_sc_hd__or2_4
X_18862_ _15121_/X _18834_/A _24384_/Q _18835_/A VGND VGND VPWR VPWR _24384_/D sky130_fd_sc_hd__o22a_4
XFILLER_84_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12005__A _11966_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17813_ _17825_/A VGND VGND VPWR VPWR _17813_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18793_ _17191_/X _18788_/X _24428_/Q _18789_/X VGND VGND VPWR VPWR _18793_/X sky130_fd_sc_hd__o22a_4
XFILLER_43_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17744_ _17744_/A _17730_/X _17744_/C VGND VGND VPWR VPWR _17745_/C sky130_fd_sc_hd__and3_4
XANTENNA__15316__A _13708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14956_ _12582_/A _14889_/B VGND VGND VPWR VPWR _14956_/X sky130_fd_sc_hd__or2_4
XFILLER_43_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23985__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14220__A _14345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13907_ _13700_/A _13907_/B _13907_/C VGND VGND VPWR VPWR _13907_/X sky130_fd_sc_hd__and3_4
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17675_ _17677_/A _17675_/B VGND VGND VPWR VPWR _17684_/B sky130_fd_sc_hd__or2_4
XFILLER_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14887_ _13987_/A _14862_/X _14870_/X _14878_/X _14886_/X VGND VGND VPWR VPWR _14887_/X
+ sky130_fd_sc_hd__a32o_4
X_19414_ _19414_/A VGND VGND VPWR VPWR _22978_/A sky130_fd_sc_hd__buf_2
XFILLER_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21940__B2 _21935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16626_ _16610_/A _23580_/Q VGND VGND VPWR VPWR _16627_/C sky130_fd_sc_hd__or2_4
X_13838_ _13690_/A VGND VGND VPWR VPWR _13896_/A sky130_fd_sc_hd__buf_2
XFILLER_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23215__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19345_ _19343_/X _18551_/X _19343_/X _20792_/A VGND VGND VPWR VPWR _19345_/X sky130_fd_sc_hd__a2bb2o_4
X_16557_ _12025_/A _16557_/B _16557_/C VGND VGND VPWR VPWR _16561_/B sky130_fd_sc_hd__and3_4
Xclkbuf_7_1_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR _24203_/CLK sky130_fd_sc_hd__clkbuf_1
X_13769_ _13731_/A _13769_/B _13769_/C VGND VGND VPWR VPWR _13769_/X sky130_fd_sc_hd__or3_4
XANTENNA__12675__A _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22496__A2 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16147__A _16147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15051__A _15050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15508_ _13735_/A _23468_/Q VGND VGND VPWR VPWR _15508_/X sky130_fd_sc_hd__or2_4
X_19276_ _19215_/A _19215_/B _19275_/Y VGND VGND VPWR VPWR _24266_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21988__A _21988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16488_ _16363_/X _16484_/X _16488_/C VGND VGND VPWR VPWR _16488_/X sky130_fd_sc_hd__or3_4
XANTENNA__20892__A _20892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12394__B _12287_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18227_ _18198_/X _18223_/X _18224_/X _18226_/X VGND VGND VPWR VPWR _18227_/X sky130_fd_sc_hd__o22a_4
X_15439_ _15436_/A _15511_/B VGND VGND VPWR VPWR _15441_/B sky130_fd_sc_hd__or2_4
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15383__B1 _15185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22248__A2 _22243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18362__A _18244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18158_ _17989_/X _17471_/X _18152_/X _18082_/X _18157_/Y VGND VGND VPWR VPWR _18158_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_117_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17109_ _15312_/X VGND VGND VPWR VPWR _17109_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18089_ _17762_/X _17660_/X _17653_/X VGND VGND VPWR VPWR _18089_/X sky130_fd_sc_hd__o21a_4
XFILLER_102_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20120_ _11567_/X VGND VGND VPWR VPWR _20120_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20051_ _20042_/X _18459_/A _20048_/X _20050_/X VGND VGND VPWR VPWR _20051_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18624__A1 _17779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13953__B _14025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23810_ _23812_/CLK _23810_/D VGND VGND VPWR VPWR _15290_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14130__A _11879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22184__B2 _22183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20953_ _24225_/Q VGND VGND VPWR VPWR _20953_/Y sky130_fd_sc_hd__inv_2
X_23741_ _23931_/CLK _23741_/D VGND VGND VPWR VPWR _23741_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20884_ _20733_/X _20883_/X _11509_/A _20686_/X VGND VGND VPWR VPWR _20884_/X sky130_fd_sc_hd__o22a_4
X_23672_ _23316_/CLK _23672_/D VGND VGND VPWR VPWR _23672_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22059__A _22052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22623_ _22390_/X _22622_/X _12159_/B _22619_/X VGND VGND VPWR VPWR _23133_/D sky130_fd_sc_hd__o22a_4
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22487__A2 _22486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12585__A _12585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22554_ _22533_/A VGND VGND VPWR VPWR _22554_/X sky130_fd_sc_hd__buf_2
XANTENNA__21898__A _21884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20498__B2 _20497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21505_ _21498_/Y _21503_/X _21504_/X _21503_/X VGND VGND VPWR VPWR _23774_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15896__A _13500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22485_ _22413_/X _22479_/X _23220_/Q _22483_/X VGND VGND VPWR VPWR _23220_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22239__A2 _22236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18272__A _18392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21436_ _21275_/X _21433_/X _13815_/B _21430_/X VGND VGND VPWR VPWR _21436_/X sky130_fd_sc_hd__o22a_4
X_24224_ _24250_/CLK _24224_/D HRESETn VGND VGND VPWR VPWR _24224_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23858__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21998__B2 _21992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16504__B _16427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24155_ _24162_/CLK _19906_/X HRESETn VGND VGND VPWR VPWR _24155_/Q sky130_fd_sc_hd__dfrtp_4
X_21367_ _21241_/X _21362_/X _12661_/B _21366_/X VGND VGND VPWR VPWR _21367_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18863__A1 _15119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14305__A _15533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18863__B2 _18835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20318_ _20229_/X _20317_/X _20213_/X VGND VGND VPWR VPWR _20318_/Y sky130_fd_sc_hd__o21ai_4
X_23106_ _23812_/CLK _23106_/D VGND VGND VPWR VPWR _15289_/B sky130_fd_sc_hd__dfxtp_4
X_24086_ _24084_/CLK _20465_/X VGND VGND VPWR VPWR _12316_/B sky130_fd_sc_hd__dfxtp_4
X_21298_ _21348_/A _21784_/B _21784_/C _21634_/D VGND VGND VPWR VPWR _21299_/A sky130_fd_sc_hd__or4_4
XANTENNA__22522__A _22536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23037_ _22968_/A _17891_/B _17952_/X VGND VGND VPWR VPWR _23037_/X sky130_fd_sc_hd__or3_4
X_20249_ _20301_/A VGND VGND VPWR VPWR _20468_/A sky130_fd_sc_hd__inv_2
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18615__A1 _17792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14959__B _14892_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20042__A _19994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20973__A2 _20972_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14810_ _14810_/A VGND VGND VPWR VPWR _14811_/A sky130_fd_sc_hd__buf_2
XANTENNA__15136__A _11954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11664__A _11664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15790_ _12458_/A _15786_/X _15790_/C VGND VGND VPWR VPWR _15790_/X sky130_fd_sc_hd__or3_4
XANTENNA__14040__A _11798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22175__B2 _22169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23238__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14741_ _13603_/A _14741_/B _14740_/X VGND VGND VPWR VPWR _14741_/X sky130_fd_sc_hd__and3_4
XFILLER_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11953_ _14906_/A VGND VGND VPWR VPWR _11954_/A sky130_fd_sc_hd__buf_2
X_23939_ _23270_/CLK _21206_/X VGND VGND VPWR VPWR _14820_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20186__B1 _19313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14975__A _14195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21922__B2 _21921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17460_ _12338_/Y _17014_/X _17022_/X _17459_/Y VGND VGND VPWR VPWR _17461_/B sky130_fd_sc_hd__o22a_4
X_14672_ _14672_/A _23556_/Q VGND VGND VPWR VPWR _14673_/C sky130_fd_sc_hd__or2_4
X_11884_ _13427_/A VGND VGND VPWR VPWR _11884_/X sky130_fd_sc_hd__buf_2
X_16411_ _11980_/X _16411_/B VGND VGND VPWR VPWR _16411_/X sky130_fd_sc_hd__and2_4
X_13623_ _13623_/A _23272_/Q VGND VGND VPWR VPWR _13624_/C sky130_fd_sc_hd__or2_4
XFILLER_38_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17391_ _17391_/A VGND VGND VPWR VPWR _17422_/A sky130_fd_sc_hd__buf_2
XANTENNA__22478__A2 _22472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12495__A _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19130_ _24309_/Q _19129_/X VGND VGND VPWR VPWR _19157_/A sky130_fd_sc_hd__and2_4
X_16342_ _16366_/A _16340_/X _16341_/X VGND VGND VPWR VPWR _16342_/X sky130_fd_sc_hd__and3_4
XFILLER_41_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20489__B2 _20488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13554_ _13554_/A _13554_/B VGND VGND VPWR VPWR _13555_/C sky130_fd_sc_hd__or2_4
XFILLER_105_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21150__A2 _21147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12505_ _13029_/A _12505_/B VGND VGND VPWR VPWR _12506_/C sky130_fd_sc_hd__or2_4
X_19061_ _24328_/Q _11513_/B _19054_/Y VGND VGND VPWR VPWR _19061_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_51_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16273_ _16252_/X _16273_/B VGND VGND VPWR VPWR _16273_/X sky130_fd_sc_hd__or2_4
X_13485_ _12905_/A _13485_/B VGND VGND VPWR VPWR _13485_/X sky130_fd_sc_hd__or2_4
XFILLER_51_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18012_ _16942_/Y VGND VGND VPWR VPWR _18012_/X sky130_fd_sc_hd__buf_2
X_15224_ _14201_/A _15220_/X _15224_/C VGND VGND VPWR VPWR _15224_/X sky130_fd_sc_hd__or3_4
X_12436_ _11610_/A VGND VGND VPWR VPWR _15013_/A sky130_fd_sc_hd__buf_2
XFILLER_51_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17106__B2 _17105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21989__A1 _21816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12942__B _23923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21989__B2 _21985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15155_ _14083_/A _23873_/Q VGND VGND VPWR VPWR _15157_/B sky130_fd_sc_hd__or2_4
XANTENNA__18854__A1 _14425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12367_ _12367_/A VGND VGND VPWR VPWR _15882_/A sky130_fd_sc_hd__buf_2
XFILLER_114_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14215__A _14215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14106_ _14997_/A VGND VGND VPWR VPWR _14318_/A sky130_fd_sc_hd__buf_2
XANTENNA__20661__A1 _20518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20661__B2 _20525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12298_ _15667_/A _12298_/B VGND VGND VPWR VPWR _12298_/X sky130_fd_sc_hd__or2_4
X_15086_ _14039_/A _15086_/B _15086_/C VGND VGND VPWR VPWR _15086_/X sky130_fd_sc_hd__or3_4
X_19963_ _17772_/X _19961_/X _19962_/Y _19957_/X VGND VGND VPWR VPWR _19963_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22432__A _20696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14037_ _14037_/A _14033_/X _14036_/X VGND VGND VPWR VPWR _14038_/C sky130_fd_sc_hd__or3_4
X_18914_ _14564_/X _18912_/X _19079_/A _18913_/X VGND VGND VPWR VPWR _24357_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22402__A2 _22392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19894_ _19933_/A _19893_/X VGND VGND VPWR VPWR _19894_/X sky130_fd_sc_hd__or2_4
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20413__A1 _18087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13773__B _13772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21048__A _21027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18845_ _15911_/X _18841_/X _24397_/Q _18842_/X VGND VGND VPWR VPWR _18845_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24322__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18776_ _16374_/X _18774_/X _20379_/A _18775_/X VGND VGND VPWR VPWR _24441_/D sky130_fd_sc_hd__o22a_4
XFILLER_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15988_ _16096_/A _23480_/Q VGND VGND VPWR VPWR _15988_/X sky130_fd_sc_hd__or2_4
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17727_ _17726_/X _17300_/X VGND VGND VPWR VPWR _17744_/A sky130_fd_sc_hd__or2_4
XFILLER_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14939_ _11645_/A VGND VGND VPWR VPWR _15072_/A sky130_fd_sc_hd__buf_2
XFILLER_110_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24163__CLK _24162_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18357__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21913__B2 _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_41_0_HCLK clkbuf_6_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_82_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17658_ _17658_/A VGND VGND VPWR VPWR _17658_/Y sky130_fd_sc_hd__inv_2
X_16609_ _11780_/X VGND VGND VPWR VPWR _16610_/A sky130_fd_sc_hd__buf_2
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17589_ _17499_/X _17589_/B VGND VGND VPWR VPWR _17589_/X sky130_fd_sc_hd__and2_4
XANTENNA__21214__C _21162_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19328_ _19328_/A VGND VGND VPWR VPWR _19328_/X sky130_fd_sc_hd__buf_2
XFILLER_52_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21141__A2 _21140_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22607__A _22600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19259_ _19223_/X VGND VGND VPWR VPWR _19259_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13013__B _23986_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16605__A _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22270_ _22095_/X _22265_/X _12580_/B _22269_/X VGND VGND VPWR VPWR _22270_/X sky130_fd_sc_hd__o22a_4
X_21221_ _21791_/A VGND VGND VPWR VPWR _21221_/X sky130_fd_sc_hd__buf_2
XANTENNA__11749__A _11803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18845__A1 _15911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19916__A _19909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14125__A _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22641__A2 _22636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16856__B1 _16840_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21152_ _20838_/X _21147_/X _14379_/B _21151_/X VGND VGND VPWR VPWR _23974_/D sky130_fd_sc_hd__o22a_4
X_20103_ _11570_/X _20134_/A VGND VGND VPWR VPWR _20103_/X sky130_fd_sc_hd__or2_4
XFILLER_67_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21083_ _20537_/X _21082_/X _24019_/Q _21079_/X VGND VGND VPWR VPWR _21083_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16340__A _16185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14779__B _14779_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20034_ _24462_/Q VGND VGND VPWR VPWR _20034_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21601__B1 _12224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12893__A1 _13491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_123_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR _23311_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_101_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17820__A2 _17816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21985_ _21985_/A VGND VGND VPWR VPWR _21985_/X sky130_fd_sc_hd__buf_2
XFILLER_113_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18267__A _18267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21904__B2 _21898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17171__A _14073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23724_ _23404_/CLK _21615_/X VGND VGND VPWR VPWR _15459_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _22456_/A VGND VGND VPWR VPWR _21287_/A sky130_fd_sc_hd__buf_2
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _20913_/A _20866_/X VGND VGND VPWR VPWR _20867_/X sky130_fd_sc_hd__or2_4
X_23655_ _23368_/CLK _21722_/X VGND VGND VPWR VPWR _13791_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15403__B _15403_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13204__A _12794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22606_ _22449_/X _22600_/X _14518_/B _22604_/X VGND VGND VPWR VPWR _22606_/X sky130_fd_sc_hd__o22a_4
XFILLER_41_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21668__B1 _23690_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20798_ _20750_/X _20797_/X _24072_/Q _20724_/X VGND VGND VPWR VPWR _24072_/D sky130_fd_sc_hd__o22a_4
X_23586_ _23522_/CLK _23586_/D VGND VGND VPWR VPWR _15285_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22517__A _22521_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22537_ _22415_/X _22536_/X _12857_/B _22533_/X VGND VGND VPWR VPWR _23187_/D sky130_fd_sc_hd__o22a_4
XFILLER_52_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20340__B1 _24092_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16515__A _16444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13270_ _13270_/A VGND VGND VPWR VPWR _13270_/X sky130_fd_sc_hd__buf_2
X_22468_ _22483_/A VGND VGND VPWR VPWR _22476_/A sky130_fd_sc_hd__buf_2
X_12221_ _12496_/A VGND VGND VPWR VPWR _12221_/X sky130_fd_sc_hd__buf_2
X_24207_ _24208_/CLK _24207_/D HRESETn VGND VGND VPWR VPWR _24207_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11659__A _11658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21419_ _21419_/A VGND VGND VPWR VPWR _21419_/X sky130_fd_sc_hd__buf_2
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18836__A1 _17181_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19826__A _19829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22399_ _22386_/X VGND VGND VPWR VPWR _22399_/X sky130_fd_sc_hd__buf_2
XANTENNA__22632__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12152_ _12152_/A _23901_/Q VGND VGND VPWR VPWR _12152_/X sky130_fd_sc_hd__or2_4
XANTENNA__24416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24138_ _24229_/CLK _19969_/Y HRESETn VGND VGND VPWR VPWR _17002_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_2_2_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13874__A _13862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12083_ _12083_/A _23901_/Q VGND VGND VPWR VPWR _12085_/B sky130_fd_sc_hd__or2_4
X_16960_ _16960_/A VGND VGND VPWR VPWR _18558_/A sky130_fd_sc_hd__inv_2
X_24069_ _23365_/CLK _20871_/X VGND VGND VPWR VPWR _14477_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_77_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21199__A2 _21197_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14689__B _14689_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15911_ _15907_/X VGND VGND VPWR VPWR _15911_/X sky130_fd_sc_hd__buf_2
X_16891_ _16891_/A _16890_/X VGND VGND VPWR VPWR _16891_/Y sky130_fd_sc_hd__nand2_4
XFILLER_81_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24186__CLK _24223_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18630_ _18630_/A VGND VGND VPWR VPWR _18630_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15842_ _12922_/A _15842_/B VGND VGND VPWR VPWR _15842_/X sky130_fd_sc_hd__and2_4
XFILLER_92_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22148__B2 _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18561_ _17792_/A _17621_/D _17966_/X _17338_/X VGND VGND VPWR VPWR _18561_/X sky130_fd_sc_hd__o22a_4
XFILLER_40_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15773_ _12795_/A _15700_/B VGND VGND VPWR VPWR _15773_/X sky130_fd_sc_hd__or2_4
X_12985_ _12947_/A _12983_/X _12984_/X VGND VGND VPWR VPWR _12985_/X sky130_fd_sc_hd__and3_4
XANTENNA__22699__A2 _22693_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17512_ _17512_/A VGND VGND VPWR VPWR _18307_/A sky130_fd_sc_hd__inv_2
X_14724_ _14722_/Y _14724_/B VGND VGND VPWR VPWR _14724_/X sky130_fd_sc_hd__or2_4
Xclkbuf_5_28_0_HCLK clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_11936_ _16130_/A VGND VGND VPWR VPWR _11936_/X sky130_fd_sc_hd__buf_2
X_18492_ _17422_/D _18491_/X _17427_/X VGND VGND VPWR VPWR _18492_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_72_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21371__A2 _21369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17443_ _17439_/Y _17014_/A _17022_/A _17667_/B VGND VGND VPWR VPWR _17524_/B sky130_fd_sc_hd__o22a_4
X_14655_ _14673_/A _14652_/X _14655_/C VGND VGND VPWR VPWR _14655_/X sky130_fd_sc_hd__and3_4
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11867_ _13968_/A VGND VGND VPWR VPWR _13654_/A sky130_fd_sc_hd__buf_2
XANTENNA__18905__A _18898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13606_ _13606_/A VGND VGND VPWR VPWR _15399_/A sky130_fd_sc_hd__buf_2
X_17374_ _11631_/A _17364_/A _17365_/A VGND VGND VPWR VPWR _17374_/X sky130_fd_sc_hd__o21a_4
X_14586_ _14727_/A _14584_/X _14586_/C VGND VGND VPWR VPWR _14586_/X sky130_fd_sc_hd__and3_4
XFILLER_92_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11798_ _11798_/A VGND VGND VPWR VPWR _11799_/A sky130_fd_sc_hd__buf_2
XANTENNA__22427__A _22112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19113_ _19113_/A _19112_/X VGND VGND VPWR VPWR _19113_/X sky130_fd_sc_hd__and2_4
X_16325_ _11700_/X VGND VGND VPWR VPWR _16364_/A sky130_fd_sc_hd__buf_2
XFILLER_53_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13537_ _13557_/A _13528_/X _13537_/C VGND VGND VPWR VPWR _13538_/C sky130_fd_sc_hd__and3_4
X_19044_ _24363_/Q VGND VGND VPWR VPWR _19044_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20882__A1 _20681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16256_ _16286_/A _16256_/B VGND VGND VPWR VPWR _16256_/X sky130_fd_sc_hd__or2_4
X_13468_ _13483_/A _13464_/X _13468_/C VGND VGND VPWR VPWR _13468_/X sky130_fd_sc_hd__or3_4
X_15207_ _14201_/A _15207_/B _15207_/C VGND VGND VPWR VPWR _15207_/X sky130_fd_sc_hd__or3_4
X_12419_ _12419_/A _12316_/B VGND VGND VPWR VPWR _12420_/C sky130_fd_sc_hd__or2_4
X_16187_ _11713_/X VGND VGND VPWR VPWR _16188_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22623__A2 _22622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13399_ _13399_/A _13399_/B _13398_/X VGND VGND VPWR VPWR _13400_/C sky130_fd_sc_hd__and3_4
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15138_ _14136_/A _15134_/X _15137_/X VGND VGND VPWR VPWR _15138_/X sky130_fd_sc_hd__or3_4
XFILLER_86_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16302__A2 _11619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22162__A _22162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15069_ _15069_/A _23903_/Q VGND VGND VPWR VPWR _15069_/X sky130_fd_sc_hd__or2_4
X_19946_ _17968_/X _18733_/X VGND VGND VPWR VPWR _19946_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16160__A _16159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19877_ _19877_/A _19877_/B VGND VGND VPWR VPWR _19877_/X sky130_fd_sc_hd__or2_4
XFILLER_25_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18828_ _18835_/A VGND VGND VPWR VPWR _18828_/X sky130_fd_sc_hd__buf_2
XFILLER_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15813__A1 _12682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21506__A _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13008__B _24018_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18759_ _18759_/A _16916_/B _17083_/A _11591_/C VGND VGND VPWR VPWR _18762_/A sky130_fd_sc_hd__or4_4
XFILLER_97_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21770_ _21555_/X _21769_/X _23625_/Q _21766_/X VGND VGND VPWR VPWR _21770_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17422__C _17422_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20721_ _24203_/Q _20614_/X _20720_/X VGND VGND VPWR VPWR _20722_/A sky130_fd_sc_hd__o21a_4
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20570__B1 _20569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18815__A _18762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13024__A _12465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20652_ _20619_/X _20651_/X VGND VGND VPWR VPWR _20652_/X sky130_fd_sc_hd__or2_4
X_23440_ _23920_/CLK _23440_/D VGND VGND VPWR VPWR _13312_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22337__A _22344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23371_ _23688_/CLK _23371_/D VGND VGND VPWR VPWR _23371_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13959__A _13959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20583_ _20493_/X _20582_/X _24304_/Q _20500_/X VGND VGND VPWR VPWR _20584_/B sky130_fd_sc_hd__o22a_4
XFILLER_20_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16335__A _16365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12863__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_48_0_HCLK clkbuf_6_24_0_HCLK/X VGND VGND VPWR VPWR _23978_/CLK sky130_fd_sc_hd__clkbuf_1
X_22322_ _23304_/Q VGND VGND VPWR VPWR _22322_/X sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_5_19_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22253_ _22286_/A VGND VGND VPWR VPWR _22269_/A sky130_fd_sc_hd__inv_2
XFILLER_69_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21204_ _21168_/A VGND VGND VPWR VPWR _21204_/X sky130_fd_sc_hd__buf_2
XFILLER_69_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22184_ _22119_/X _22179_/X _23403_/Q _22183_/X VGND VGND VPWR VPWR _23403_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22072__A _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21135_ _20553_/X _21133_/X _23986_/Q _21130_/X VGND VGND VPWR VPWR _21135_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22378__B2 _22372_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21066_ _21058_/Y _21065_/X _20277_/X _21065_/X VGND VGND VPWR VPWR _21066_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20389__B1 _20288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14302__B _14302_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20017_ _20017_/A VGND VGND VPWR VPWR _24128_/D sky130_fd_sc_hd__inv_2
XFILLER_58_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21050__B2 _21048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12103__A _12098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21416__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20320__A _20447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15414__A _13641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21889__B1 _13085_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12770_ _12753_/X _12770_/B _12769_/X VGND VGND VPWR VPWR _12787_/B sky130_fd_sc_hd__or3_4
XFILLER_15_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21968_ _21967_/X VGND VGND VPWR VPWR _22002_/A sky130_fd_sc_hd__buf_2
XFILLER_55_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _13708_/A VGND VGND VPWR VPWR _13998_/A sky130_fd_sc_hd__buf_2
X_23707_ _23707_/CLK _23707_/D VGND VGND VPWR VPWR _23707_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ _20875_/A _20358_/B VGND VGND VPWR VPWR _20919_/X sky130_fd_sc_hd__or2_4
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ _21835_/X _21894_/X _23563_/Q _21898_/X VGND VGND VPWR VPWR _23563_/D sky130_fd_sc_hd__o22a_4
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14463_/A _14506_/B VGND VGND VPWR VPWR _14441_/C sky130_fd_sc_hd__or2_4
XFILLER_70_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _15611_/A _12421_/A _12965_/A _11652_/D VGND VGND VPWR VPWR _11652_/X sky130_fd_sc_hd__or4_4
X_23638_ _23920_/CLK _23638_/D VGND VGND VPWR VPWR _12424_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_42_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18506__B1 _18497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21105__A2 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21151__A _21130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _14371_/A VGND VGND VPWR VPWR _15631_/A sky130_fd_sc_hd__buf_2
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11583_ _17024_/C _17030_/B VGND VGND VPWR VPWR _11634_/B sky130_fd_sc_hd__or2_4
X_23569_ _24082_/CLK _21890_/X VGND VGND VPWR VPWR _23569_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16110_ _16107_/A _22307_/A VGND VGND VPWR VPWR _16112_/B sky130_fd_sc_hd__or2_4
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _13301_/A _24048_/Q VGND VGND VPWR VPWR _13322_/X sky130_fd_sc_hd__or2_4
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17090_ _18101_/A VGND VGND VPWR VPWR _17090_/X sky130_fd_sc_hd__buf_2
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16041_ _16069_/A _23544_/Q VGND VGND VPWR VPWR _16042_/C sky130_fd_sc_hd__or2_4
X_13253_ _13260_/A _13193_/B VGND VGND VPWR VPWR _13253_/X sky130_fd_sc_hd__or2_4
XANTENNA__18809__A1 _15121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19556__A _19877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22605__A2 _22600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18809__B2 _18782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12204_ _15432_/A VGND VGND VPWR VPWR _12496_/A sky130_fd_sc_hd__buf_2
XFILLER_89_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_5_0_HCLK clkbuf_6_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13184_ _15695_/A _13180_/X _13183_/X VGND VGND VPWR VPWR _13184_/X sky130_fd_sc_hd__or3_4
X_19800_ _19454_/A _19800_/B VGND VGND VPWR VPWR _19800_/X sky130_fd_sc_hd__or2_4
XANTENNA__20092__A2 _20091_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12135_ _11675_/X _12127_/X _12134_/X VGND VGND VPWR VPWR _12135_/X sky130_fd_sc_hd__and3_4
XANTENNA__17076__A _18418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17992_ _17532_/Y _17568_/Y _17571_/Y VGND VGND VPWR VPWR _18083_/A sky130_fd_sc_hd__o21a_4
XANTENNA__23576__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22369__B2 _22365_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16943_ _16943_/A VGND VGND VPWR VPWR _16985_/A sky130_fd_sc_hd__inv_2
X_19731_ _19857_/C _19726_/X _19730_/X VGND VGND VPWR VPWR _19731_/X sky130_fd_sc_hd__a21bo_4
X_12066_ _12065_/X _23997_/Q VGND VGND VPWR VPWR _12067_/C sky130_fd_sc_hd__or2_4
XFILLER_77_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16874_ _16824_/D _13593_/B _13578_/A VGND VGND VPWR VPWR _16874_/X sky130_fd_sc_hd__o21a_4
X_19662_ _19662_/A VGND VGND VPWR VPWR _19663_/A sky130_fd_sc_hd__buf_2
XANTENNA__12013__A _12020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15825_ _12520_/X _15825_/B VGND VGND VPWR VPWR _15826_/C sky130_fd_sc_hd__or2_4
X_18613_ _17724_/X _18612_/Y _16966_/A _18611_/X VGND VGND VPWR VPWR _18613_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21326__A _21319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19593_ _19428_/A _19441_/A VGND VGND VPWR VPWR _19593_/X sky130_fd_sc_hd__or2_4
XFILLER_65_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12948__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11852__A _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15756_ _13109_/A _15754_/X _15755_/X VGND VGND VPWR VPWR _15760_/B sky130_fd_sc_hd__and3_4
X_18544_ _18499_/X _17395_/X _18500_/X VGND VGND VPWR VPWR _18544_/X sky130_fd_sc_hd__a21o_4
X_12968_ _12980_/A _23379_/Q VGND VGND VPWR VPWR _12970_/B sky130_fd_sc_hd__or2_4
XFILLER_59_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21344__A2 _21340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22541__B2 _22540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12667__B _12667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14707_ _14714_/A _14635_/B VGND VGND VPWR VPWR _14707_/X sky130_fd_sc_hd__or2_4
XANTENNA__11571__B IRQ[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11919_ _11983_/A VGND VGND VPWR VPWR _11993_/A sky130_fd_sc_hd__buf_2
X_18475_ _18464_/X _18469_/Y _18471_/X _18473_/X _18474_/Y VGND VGND VPWR VPWR _18475_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15043__B _23679_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15687_ _15687_/A _15687_/B _15687_/C VGND VGND VPWR VPWR _15687_/X sky130_fd_sc_hd__and3_4
X_12899_ _12870_/A _12899_/B _12899_/C VGND VGND VPWR VPWR _12900_/C sky130_fd_sc_hd__and3_4
X_17426_ _17422_/B _17424_/X _17425_/X VGND VGND VPWR VPWR _17426_/X sky130_fd_sc_hd__o21a_4
X_14638_ _14172_/A _14637_/X VGND VGND VPWR VPWR _14638_/X sky130_fd_sc_hd__and2_4
XANTENNA__22157__A _22153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14882__B _14882_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21061__A _21112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17357_ _17356_/X VGND VGND VPWR VPWR _17361_/A sky130_fd_sc_hd__inv_2
XFILLER_105_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14569_ _14138_/X _14569_/B VGND VGND VPWR VPWR _14569_/X sky130_fd_sc_hd__or2_4
XANTENNA__12683__A _12553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16308_ _11700_/X VGND VGND VPWR VPWR _16322_/A sky130_fd_sc_hd__buf_2
X_17288_ _17283_/Y _17012_/A _17018_/X _17287_/X VGND VGND VPWR VPWR _17313_/B sky130_fd_sc_hd__o22a_4
X_19027_ _19027_/A VGND VGND VPWR VPWR _19027_/X sky130_fd_sc_hd__buf_2
X_16239_ _16081_/X _16239_/B VGND VGND VPWR VPWR _16239_/X sky130_fd_sc_hd__or2_4
XANTENNA__18370__A _17874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19929_ _19996_/A VGND VGND VPWR VPWR _19929_/X sky130_fd_sc_hd__buf_2
XFILLER_116_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15218__B _23873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13019__A _13019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21032__B2 _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22940_ _18528_/X _22945_/B VGND VGND VPWR VPWR _22941_/C sky130_fd_sc_hd__or2_4
XFILLER_56_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22871_ _17272_/Y _22863_/X _22853_/X _22870_/X VGND VGND VPWR VPWR _22872_/B sky130_fd_sc_hd__o22a_4
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20140__A IRQ[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12858__A _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21822_ _21821_/X _21817_/X _13174_/B _21812_/X VGND VGND VPWR VPWR _23601_/D sky130_fd_sc_hd__o22a_4
XFILLER_37_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21335__A2 _21333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_11_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21753_ _21526_/X _21748_/X _12668_/B _21752_/X VGND VGND VPWR VPWR _23637_/D sky130_fd_sc_hd__o22a_4
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18545__A _18697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20704_ _20468_/A VGND VGND VPWR VPWR _20704_/X sky130_fd_sc_hd__buf_2
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24472_ _24241_/CLK _24472_/D HRESETn VGND VGND VPWR VPWR _19986_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21684_ _21684_/A _21784_/B _21684_/C _21784_/D VGND VGND VPWR VPWR _21684_/X sky130_fd_sc_hd__or4_4
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23423_ _23487_/CLK _22148_/X VGND VGND VPWR VPWR _23423_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13689__A _14207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21099__B2 _21093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22296__B1 _15255_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20635_ _24206_/Q _20614_/X _20634_/Y VGND VGND VPWR VPWR _22112_/A sky130_fd_sc_hd__o21a_4
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20566_ _20603_/A _20566_/B VGND VGND VPWR VPWR _20566_/Y sky130_fd_sc_hd__nor2_4
X_23354_ _23354_/CLK _23354_/D VGND VGND VPWR VPWR _16383_/B sky130_fd_sc_hd__dfxtp_4
X_22305_ _16259_/B VGND VGND VPWR VPWR _22305_/X sky130_fd_sc_hd__buf_2
X_20497_ _20497_/A VGND VGND VPWR VPWR _20497_/X sky130_fd_sc_hd__buf_2
X_23285_ _23987_/CLK _22352_/X VGND VGND VPWR VPWR _12607_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22599__B2 _22597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22236_ _22207_/A VGND VGND VPWR VPWR _22236_/X sky130_fd_sc_hd__buf_2
XFILLER_69_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20315__A _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11937__A _11936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22167_ _22091_/X _22165_/X _16135_/B _22162_/X VGND VGND VPWR VPWR _23415_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15409__A _15432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14313__A _11911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21118_ _21118_/A VGND VGND VPWR VPWR _21133_/A sky130_fd_sc_hd__buf_2
XFILLER_43_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22098_ _22413_/A VGND VGND VPWR VPWR _22098_/X sky130_fd_sc_hd__buf_2
XANTENNA__23012__A2 _16945_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13940_ _13968_/A _13940_/B _13940_/C VGND VGND VPWR VPWR _13941_/C sky130_fd_sc_hd__and3_4
X_21049_ _20838_/X _21044_/X _14305_/B _21048_/X VGND VGND VPWR VPWR _24038_/D sky130_fd_sc_hd__o22a_4
XFILLER_115_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13871_ _13871_/A VGND VGND VPWR VPWR _13872_/A sky130_fd_sc_hd__buf_2
XFILLER_75_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23064__C _23064_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15610_ _14499_/A _15610_/B _15610_/C VGND VGND VPWR VPWR _15611_/C sky130_fd_sc_hd__and3_4
XFILLER_90_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11672__A _13133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12822_ _12822_/A _12822_/B _12821_/X VGND VGND VPWR VPWR _12840_/B sky130_fd_sc_hd__and3_4
X_16590_ _11903_/A _23868_/Q VGND VGND VPWR VPWR _16590_/X sky130_fd_sc_hd__or2_4
XFILLER_90_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22523__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15541_ _14464_/A _15541_/B _15541_/C VGND VGND VPWR VPWR _15541_/X sky130_fd_sc_hd__and3_4
X_12753_ _12955_/A VGND VGND VPWR VPWR _12753_/X sky130_fd_sc_hd__buf_2
XFILLER_91_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _16071_/A VGND VGND VPWR VPWR _11803_/A sky130_fd_sc_hd__buf_2
X_18260_ _18228_/X _18259_/X _20010_/A _18228_/X VGND VGND VPWR VPWR _24467_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _12638_/A _15470_/X _15471_/X VGND VGND VPWR VPWR _15472_/X sky130_fd_sc_hd__and3_4
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _13046_/A _23508_/Q VGND VGND VPWR VPWR _12685_/C sky130_fd_sc_hd__or2_4
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17141_/X _17209_/X _17154_/X _17210_/X VGND VGND VPWR VPWR _17211_/X sky130_fd_sc_hd__o22a_4
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _13918_/A _14423_/B _14422_/X VGND VGND VPWR VPWR _14423_/X sky130_fd_sc_hd__and3_4
XFILLER_54_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13599__A _14782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _17069_/A _11579_/X VGND VGND VPWR VPWR _19927_/A sky130_fd_sc_hd__or2_4
X_18191_ _18191_/A _18190_/X VGND VGND VPWR VPWR _18191_/X sky130_fd_sc_hd__or2_4
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17142_ _15381_/X _17161_/A _16814_/B _17157_/A VGND VGND VPWR VPWR _17142_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14354_ _14359_/A VGND VGND VPWR VPWR _15614_/A sky130_fd_sc_hd__buf_2
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _20379_/A IRQ[26] VGND VGND VPWR VPWR _11566_/X sky130_fd_sc_hd__and2_4
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13305_ _13428_/A _23536_/Q VGND VGND VPWR VPWR _13305_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_31_0_HCLK clkbuf_7_30_0_HCLK/A VGND VGND VPWR VPWR _23391_/CLK sky130_fd_sc_hd__clkbuf_1
X_17073_ _18728_/B _17073_/B VGND VGND VPWR VPWR _17073_/X sky130_fd_sc_hd__or2_4
XFILLER_116_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14285_ _15534_/A _14283_/X _14284_/X VGND VGND VPWR VPWR _14285_/X sky130_fd_sc_hd__and3_4
XANTENNA__16703__A _12096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_94_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR _23485_/CLK sky130_fd_sc_hd__clkbuf_1
X_16024_ _16037_/A _24024_/Q VGND VGND VPWR VPWR _16027_/B sky130_fd_sc_hd__or2_4
XFILLER_100_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13236_ _15484_/A _13227_/X _13236_/C VGND VGND VPWR VPWR _13237_/C sky130_fd_sc_hd__and3_4
XFILLER_6_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19455__A1 _24157_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11847__A _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21262__B2 _21254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13167_ _12435_/A _13165_/X _13166_/X VGND VGND VPWR VPWR _13167_/X sky130_fd_sc_hd__and3_4
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14223__A _14039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12118_ _12152_/A _12118_/B VGND VGND VPWR VPWR _12118_/X sky130_fd_sc_hd__or2_4
XFILLER_112_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11566__B IRQ[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13098_ _13098_/A _23314_/Q VGND VGND VPWR VPWR _13100_/B sky130_fd_sc_hd__or2_4
X_17975_ _17975_/A VGND VGND VPWR VPWR _17975_/X sky130_fd_sc_hd__buf_2
XFILLER_61_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22440__A _22384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17218__B1 _14988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_HCLK clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19714_ _19744_/A _19643_/A _19600_/B _19784_/B _19759_/B VGND VGND VPWR VPWR _19714_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_84_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21014__B2 _21013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22211__B1 _16791_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12049_ _12044_/X _12049_/B _12049_/C VGND VGND VPWR VPWR _12050_/C sky130_fd_sc_hd__and3_4
X_16926_ _16925_/Y VGND VGND VPWR VPWR _16927_/A sky130_fd_sc_hd__buf_2
XFILLER_65_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19645_ _19645_/A VGND VGND VPWR VPWR _19857_/C sky130_fd_sc_hd__buf_2
X_16857_ _15386_/X VGND VGND VPWR VPWR _16857_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15054__A _14046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15808_ _12879_/A _15863_/B VGND VGND VPWR VPWR _15810_/B sky130_fd_sc_hd__or2_4
XFILLER_81_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16788_ _16772_/A _16788_/B VGND VGND VPWR VPWR _16788_/X sky130_fd_sc_hd__or2_4
X_19576_ _19538_/A VGND VGND VPWR VPWR _19639_/A sky130_fd_sc_hd__inv_2
XFILLER_59_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21317__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12397__B _24054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15739_ _15751_/A _15667_/B VGND VGND VPWR VPWR _15739_/X sky130_fd_sc_hd__or2_4
X_18527_ _18527_/A VGND VGND VPWR VPWR _18527_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15989__A _15997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18194__B2 _18193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18458_ _18171_/A VGND VGND VPWR VPWR _18458_/X sky130_fd_sc_hd__buf_2
XFILLER_72_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17941__A1 _18327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17409_ _17409_/A _17408_/Y VGND VGND VPWR VPWR _17621_/A sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_3_5_0_HCLK_A clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18389_ _18266_/A _17370_/X VGND VGND VPWR VPWR _18389_/X sky130_fd_sc_hd__and2_4
XANTENNA__15501__B _23084_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20420_ _20396_/X _20419_/X _24088_/Q _20374_/X VGND VGND VPWR VPWR _24088_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20828__A1 _20622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18812__B _18866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24101__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20351_ _24251_/Q VGND VGND VPWR VPWR _20351_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16613__A _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23070_ _17052_/A VGND VGND VPWR VPWR HSIZE[1] sky130_fd_sc_hd__buf_2
X_20282_ _20282_/A VGND VGND VPWR VPWR _20282_/X sky130_fd_sc_hd__buf_2
XANTENNA__20135__A _24432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22021_ _22020_/X VGND VGND VPWR VPWR _22021_/X sky130_fd_sc_hd__buf_2
XFILLER_66_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16332__B _23993_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19997__A2 _19985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19924__A _20190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14133__A _14315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17209__B1 _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17444__A _12992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23972_ _23363_/CLK _23972_/D VGND VGND VPWR VPWR _14680_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22923_ _19201_/X _22920_/X _22923_/C VGND VGND VPWR VPWR HADDR[7] sky130_fd_sc_hd__and3_4
XFILLER_84_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12588__A _12655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22854_ _19893_/X VGND VGND VPWR VPWR _22854_/X sky130_fd_sc_hd__buf_2
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21308__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22505__B2 _22504_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21805_ _21817_/A VGND VGND VPWR VPWR _21805_/X sky130_fd_sc_hd__buf_2
XANTENNA__15899__A _15892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22785_ _17115_/Y _22782_/X VGND VGND VPWR VPWR HWDATA[2] sky130_fd_sc_hd__nor2_4
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21736_ _21740_/A VGND VGND VPWR VPWR _21752_/A sky130_fd_sc_hd__inv_2
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16507__B _16430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24455_ _24202_/CLK _24455_/D HRESETn VGND VGND VPWR VPWR _24455_/Q sky130_fd_sc_hd__dfrtp_4
X_21667_ _21550_/X _21662_/X _23691_/Q _21666_/X VGND VGND VPWR VPWR _23691_/D sky130_fd_sc_hd__o22a_4
XFILLER_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14308__A _15552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23406_ _23922_/CLK _22180_/X VGND VGND VPWR VPWR _15758_/B sky130_fd_sc_hd__dfxtp_4
X_20618_ _16891_/A _20618_/B VGND VGND VPWR VPWR _20802_/A sky130_fd_sc_hd__and2_4
X_24386_ _24425_/CLK _24386_/D HRESETn VGND VGND VPWR VPWR _24386_/Q sky130_fd_sc_hd__dfrtp_4
X_21598_ _21605_/A VGND VGND VPWR VPWR _21598_/X sky130_fd_sc_hd__buf_2
XFILLER_32_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21492__A1 _21282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23337_ _23561_/CLK _23337_/D VGND VGND VPWR VPWR _23337_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_18_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_18_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_20549_ _20444_/X _20540_/Y _20547_/X _20548_/Y _20459_/X VGND VGND VPWR VPWR _20550_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21492__B2 _21488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14070_ _14847_/A _14070_/B _14069_/X VGND VGND VPWR VPWR _14070_/X sky130_fd_sc_hd__or3_4
XFILLER_49_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23268_ _23522_/CLK _23268_/D VGND VGND VPWR VPWR _14667_/B sky130_fd_sc_hd__dfxtp_4
X_13021_ _12494_/A _13021_/B _13021_/C VGND VGND VPWR VPWR _13021_/X sky130_fd_sc_hd__and3_4
XANTENNA__11667__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22219_ _22219_/A VGND VGND VPWR VPWR _22219_/X sky130_fd_sc_hd__buf_2
XFILLER_45_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23199_ _23889_/CLK _22513_/X VGND VGND VPWR VPWR _23199_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14043__A _14815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19553__B HRDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14978__A _15074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13882__A _13910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14972_ _11642_/A _14970_/X _14972_/C VGND VGND VPWR VPWR _14976_/B sky130_fd_sc_hd__and3_4
X_17760_ _17677_/X _17678_/X _17758_/X _17759_/X VGND VGND VPWR VPWR _17760_/X sky130_fd_sc_hd__or4_4
XANTENNA__21547__A2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13923_ _13837_/X _13920_/X _13922_/Y VGND VGND VPWR VPWR _16840_/B sky130_fd_sc_hd__a21o_4
X_16711_ _11982_/X _16711_/B VGND VGND VPWR VPWR _16711_/X sky130_fd_sc_hd__and2_4
XFILLER_75_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17691_ _17662_/X _17687_/Y _17755_/B _17690_/Y VGND VGND VPWR VPWR _17692_/A sky130_fd_sc_hd__a211o_4
XFILLER_48_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12498__A _12497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16642_ _16670_/A _23548_/Q VGND VGND VPWR VPWR _16643_/C sky130_fd_sc_hd__or2_4
X_19430_ _16997_/X _19430_/B VGND VGND VPWR VPWR _19433_/A sky130_fd_sc_hd__or2_4
X_13854_ _13884_/A _13846_/X _13854_/C VGND VGND VPWR VPWR _13854_/X sky130_fd_sc_hd__or3_4
XFILLER_35_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12805_ _12753_/X _12805_/B _12805_/C VGND VGND VPWR VPWR _12806_/C sky130_fd_sc_hd__or3_4
X_16573_ _16569_/A _16573_/B _16573_/C VGND VGND VPWR VPWR _16577_/B sky130_fd_sc_hd__and3_4
X_19361_ _17000_/A _18013_/B _18174_/C VGND VGND VPWR VPWR _19361_/X sky130_fd_sc_hd__o21a_4
X_13785_ _13608_/A _23751_/Q VGND VGND VPWR VPWR _13785_/X sky130_fd_sc_hd__or2_4
X_15524_ _12320_/A _15522_/X _15523_/X VGND VGND VPWR VPWR _15524_/X sky130_fd_sc_hd__and3_4
X_18312_ _18198_/X _18310_/X _18224_/X _18311_/X VGND VGND VPWR VPWR _18312_/X sky130_fd_sc_hd__o22a_4
XFILLER_43_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12736_ _15693_/A _24084_/Q VGND VGND VPWR VPWR _12737_/C sky130_fd_sc_hd__or2_4
X_19292_ _24258_/Q _19207_/B _19291_/Y VGND VGND VPWR VPWR _19292_/X sky130_fd_sc_hd__o21a_4
XFILLER_91_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17923__B2 _17922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12945__B _12945_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18243_ _18297_/A _17447_/A VGND VGND VPWR VPWR _18243_/X sky130_fd_sc_hd__and2_4
X_15455_ _15487_/A _15455_/B VGND VGND VPWR VPWR _15455_/X sky130_fd_sc_hd__or2_4
X_12667_ _12660_/A _12667_/B VGND VGND VPWR VPWR _12667_/X sky130_fd_sc_hd__or2_4
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18913__A _18877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ _15598_/A _14327_/B VGND VGND VPWR VPWR _14406_/X sky130_fd_sc_hd__or2_4
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ _11618_/A VGND VGND VPWR VPWR _11618_/X sky130_fd_sc_hd__buf_2
X_18174_ _24130_/Q _18174_/B _18174_/C _18174_/D VGND VGND VPWR VPWR _18174_/X sky130_fd_sc_hd__and4_4
X_15386_ _15124_/X _15385_/X _15384_/A _15382_/X VGND VGND VPWR VPWR _15386_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19676__A1 _16997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12598_ _12598_/A VGND VGND VPWR VPWR _12599_/A sky130_fd_sc_hd__buf_2
XANTENNA__19676__B2 HRDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22435__A _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17125_ _17105_/B VGND VGND VPWR VPWR _17125_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14337_ _11669_/A VGND VGND VPWR VPWR _15643_/A sky130_fd_sc_hd__buf_2
X_11549_ _20706_/A IRQ[12] VGND VGND VPWR VPWR _11549_/X sky130_fd_sc_hd__and2_4
XFILLER_32_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21483__B2 _21481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16433__A _16121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17056_ _17083_/B _17051_/X _17054_/X _20206_/A _17561_/B VGND VGND VPWR VPWR _17057_/A
+ sky130_fd_sc_hd__a32o_4
X_14268_ _12233_/X _14268_/B VGND VGND VPWR VPWR _14268_/X sky130_fd_sc_hd__or2_4
XFILLER_48_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16007_ _11843_/X _11619_/X _15973_/X _11597_/X _16006_/X VGND VGND VPWR VPWR _16007_/X
+ sky130_fd_sc_hd__a32o_4
X_13219_ _11671_/A _13219_/B _13219_/C VGND VGND VPWR VPWR _13237_/B sky130_fd_sc_hd__and3_4
XANTENNA__23144__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14199_ _14205_/A _23273_/Q VGND VGND VPWR VPWR _14200_/C sky130_fd_sc_hd__or2_4
XFILLER_63_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13792__A _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17958_ _18066_/A _17540_/A VGND VGND VPWR VPWR _17959_/D sky130_fd_sc_hd__and2_4
XANTENNA__22735__A1 SYSTICKCLKDIV[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16909_ _16910_/A _16909_/B VGND VGND VPWR VPWR _17088_/A sky130_fd_sc_hd__or2_4
X_17889_ _17889_/A VGND VGND VPWR VPWR _18342_/A sky130_fd_sc_hd__buf_2
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19628_ _19556_/Y _19621_/A VGND VGND VPWR VPWR _19628_/X sky130_fd_sc_hd__and2_4
XFILLER_96_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21514__A _21799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13016__B _23538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19559_ _19559_/A VGND VGND VPWR VPWR _19766_/A sky130_fd_sc_hd__buf_2
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17711__B _17393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19364__B1 _19306_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22570_ _22564_/Y _22569_/X _22388_/X _22569_/X VGND VGND VPWR VPWR _22570_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21710__A2 _21705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21521_ _21519_/X _21520_/X _23768_/Q _21515_/X VGND VGND VPWR VPWR _23768_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13032__A _13032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24240_ _24239_/CLK _24240_/D HRESETn VGND VGND VPWR VPWR _24240_/Q sky130_fd_sc_hd__dfrtp_4
X_21452_ _21467_/A VGND VGND VPWR VPWR _21452_/X sky130_fd_sc_hd__buf_2
X_20403_ _20403_/A VGND VGND VPWR VPWR _20403_/X sky130_fd_sc_hd__buf_2
X_21383_ _21383_/A VGND VGND VPWR VPWR _21383_/X sky130_fd_sc_hd__buf_2
X_24171_ _24293_/CLK _24171_/D HRESETn VGND VGND VPWR VPWR _17052_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17439__A _12924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12871__A _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16343__A _16364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23122_ _23122_/CLK _22638_/X VGND VGND VPWR VPWR _13111_/B sky130_fd_sc_hd__dfxtp_4
X_20334_ _24252_/Q VGND VGND VPWR VPWR _20334_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20265_ _20517_/A VGND VGND VPWR VPWR _20493_/A sky130_fd_sc_hd__buf_2
X_23053_ _23048_/A _23053_/B _23053_/C VGND VGND VPWR VPWR _23053_/X sky130_fd_sc_hd__and3_4
XANTENNA__21226__B2 _21218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21777__A2 _21776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22004_ _21843_/X _22002_/X _13698_/B _21999_/X VGND VGND VPWR VPWR _22004_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20196_ _20196_/A _20196_/B _20195_/X VGND VGND VPWR VPWR _21212_/B sky130_fd_sc_hd__or3_4
XANTENNA__14798__A _13862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22726__A1 _19909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23955_ _23827_/CLK _23955_/D VGND VGND VPWR VPWR _23955_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_9_0_HCLK clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22906_ _22906_/A VGND VGND VPWR VPWR HADDR[4] sky130_fd_sc_hd__inv_2
XFILLER_45_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23886_ _23922_/CLK _23886_/D VGND VGND VPWR VPWR _15747_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12111__A _11966_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22837_ _22837_/A VGND VGND VPWR VPWR HWDATA[18] sky130_fd_sc_hd__inv_2
XFILLER_60_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18158__A1 _17989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15422__A _13651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13570_ _12754_/X _13568_/X _13570_/C VGND VGND VPWR VPWR _13570_/X sky130_fd_sc_hd__and3_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22768_ _22768_/A _22767_/Y _22768_/C VGND VGND VPWR VPWR _24101_/D sky130_fd_sc_hd__and3_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23061__D _19933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21701__A2 _21698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12521_ _12520_/X _12640_/B VGND VGND VPWR VPWR _12522_/C sky130_fd_sc_hd__or2_4
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21719_ _21690_/A VGND VGND VPWR VPWR _21719_/X sky130_fd_sc_hd__buf_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19829__A _19829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22699_ _20748_/A _22693_/X _23082_/Q _22697_/X VGND VGND VPWR VPWR _23082_/D sky130_fd_sc_hd__o22a_4
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14038__A _14055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _14186_/A _15240_/B VGND VGND VPWR VPWR _15242_/B sky130_fd_sc_hd__or2_4
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12452_ _12887_/A VGND VGND VPWR VPWR _12522_/A sky130_fd_sc_hd__buf_2
X_24438_ _24277_/CLK _24438_/D HRESETn VGND VGND VPWR VPWR _24438_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22255__A _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15171_ _14117_/A _15169_/X _15170_/X VGND VGND VPWR VPWR _15171_/X sky130_fd_sc_hd__and3_4
XANTENNA__21465__B2 _21460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22662__B1 _14962_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12383_ _12383_/A VGND VGND VPWR VPWR _12958_/A sky130_fd_sc_hd__buf_2
X_24369_ _23358_/CLK _24369_/D HRESETn VGND VGND VPWR VPWR _19010_/A sky130_fd_sc_hd__dfstp_4
X_14122_ _14990_/A _23561_/Q VGND VGND VPWR VPWR _14122_/X sky130_fd_sc_hd__or2_4
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14053_ _14065_/A _14053_/B _14052_/X VGND VGND VPWR VPWR _14054_/C sky130_fd_sc_hd__and3_4
X_18930_ _18930_/A VGND VGND VPWR VPWR _18931_/A sky130_fd_sc_hd__inv_2
XANTENNA__22414__B1 _12758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13004_ _13004_/A _13000_/X _13004_/C VGND VGND VPWR VPWR _13004_/X sky130_fd_sc_hd__or3_4
XFILLER_97_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21768__A2 _21762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18861_ _15249_/X _18855_/X _24385_/Q _18856_/X VGND VGND VPWR VPWR _18861_/X sky130_fd_sc_hd__o22a_4
X_17812_ _17812_/A VGND VGND VPWR VPWR _17812_/X sky130_fd_sc_hd__buf_2
X_18792_ _15911_/X _18788_/X _20656_/A _18789_/X VGND VGND VPWR VPWR _24429_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22717__B2 _23064_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14955_ _11646_/A _23872_/Q VGND VGND VPWR VPWR _14955_/X sky130_fd_sc_hd__or2_4
X_17743_ _17743_/A _17743_/B _17742_/X VGND VGND VPWR VPWR _17744_/C sky130_fd_sc_hd__or3_4
XFILLER_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13906_ _13910_/A _13906_/B VGND VGND VPWR VPWR _13907_/C sky130_fd_sc_hd__or2_4
X_14886_ _13957_/A _14885_/X VGND VGND VPWR VPWR _14886_/X sky130_fd_sc_hd__and2_4
X_17674_ _17674_/A _17506_/X VGND VGND VPWR VPWR _17675_/B sky130_fd_sc_hd__or2_4
XANTENNA__21940__A2 _21938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19413_ _18653_/X _24191_/Q _19377_/X _17736_/A VGND VGND VPWR VPWR _24191_/D sky130_fd_sc_hd__o22a_4
X_13837_ _13594_/X _13595_/X _13806_/X _11595_/A _13836_/X VGND VGND VPWR VPWR _13837_/X
+ sky130_fd_sc_hd__a32o_4
X_16625_ _16617_/A _23932_/Q VGND VGND VPWR VPWR _16627_/B sky130_fd_sc_hd__or2_4
XFILLER_90_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18149__A1 _18274_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12956__A _13118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11860__A _13004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16556_ _12024_/A _23580_/Q VGND VGND VPWR VPWR _16557_/C sky130_fd_sc_hd__or2_4
X_19344_ _19340_/X _18530_/X _19343_/X _24233_/Q VGND VGND VPWR VPWR _24233_/D sky130_fd_sc_hd__a2bb2o_4
X_13768_ _15491_/A _13766_/X _13768_/C VGND VGND VPWR VPWR _13769_/C sky130_fd_sc_hd__and3_4
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12719_ _12286_/X _23956_/Q VGND VGND VPWR VPWR _12720_/C sky130_fd_sc_hd__or2_4
X_15507_ _12626_/A _15503_/X _15507_/C VGND VGND VPWR VPWR _15515_/B sky130_fd_sc_hd__or3_4
X_16487_ _16499_/A _16487_/B _16487_/C VGND VGND VPWR VPWR _16488_/C sky130_fd_sc_hd__and3_4
X_19275_ _19216_/B VGND VGND VPWR VPWR _19275_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13699_ _13699_/A _13696_/X _13699_/C VGND VGND VPWR VPWR _13699_/X sky130_fd_sc_hd__and3_4
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15438_ _13670_/A _15438_/B _15437_/X VGND VGND VPWR VPWR _15442_/B sky130_fd_sc_hd__and3_4
X_18226_ _17665_/X _18225_/X _17665_/X _18225_/X VGND VGND VPWR VPWR _18226_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22165__A _22172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24345__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13787__A _13651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15369_ _13992_/A _15365_/X _15369_/C VGND VGND VPWR VPWR _15369_/X sky130_fd_sc_hd__or3_4
X_18157_ _18191_/A _18156_/X _17527_/Y VGND VGND VPWR VPWR _18157_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_102_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17259__A _17259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12691__A _12691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24092__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17108_ _17201_/A VGND VGND VPWR VPWR _17860_/A sky130_fd_sc_hd__inv_2
X_18088_ _17950_/X _18061_/Y _18022_/X _18087_/X VGND VGND VPWR VPWR _18088_/X sky130_fd_sc_hd__o22a_4
X_17039_ _17039_/A VGND VGND VPWR VPWR _17039_/X sky130_fd_sc_hd__buf_2
XANTENNA__21208__B2 _21165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22405__B1 _23256_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20050_ _18478_/X _20033_/X _20049_/Y _20044_/X VGND VGND VPWR VPWR _20050_/X sky130_fd_sc_hd__o22a_4
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22708__B2 _22704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20719__B1 _20718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15226__B _23809_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22184__A2 _22179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18818__A _18834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23740_ _23931_/CLK _23740_/D VGND VGND VPWR VPWR _23740_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20952_ _18700_/X _20332_/A _20640_/X _20951_/Y VGND VGND VPWR VPWR _20952_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21392__B1 _14780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ _24084_/CLK _21700_/X VGND VGND VPWR VPWR _23671_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _20403_/A _20882_/X _19209_/A _20736_/X VGND VGND VPWR VPWR _20883_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12866__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16338__A _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11770__A _12822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22622_ _22636_/A VGND VGND VPWR VPWR _22622_/X sky130_fd_sc_hd__buf_2
XANTENNA__15242__A _15203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16057__B _23416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22553_ _22444_/X _22550_/X _13784_/B _22547_/X VGND VGND VPWR VPWR _23175_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22892__B1 _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19649__A HRDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21504_ _21789_/A VGND VGND VPWR VPWR _21504_/X sky130_fd_sc_hd__buf_2
XFILLER_22_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22484_ _22410_/X _22479_/X _12667_/B _22483_/X VGND VGND VPWR VPWR _23221_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12188__A1 _12116_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22075__A _20314_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24223_ _24223_/CLK _24223_/D HRESETn VGND VGND VPWR VPWR _20997_/A sky130_fd_sc_hd__dfrtp_4
X_21435_ _21273_/X _21433_/X _13662_/B _21430_/X VGND VGND VPWR VPWR _21435_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22644__B1 _15689_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21998__A2 _21995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24154_ _24293_/CLK _19907_/X HRESETn VGND VGND VPWR VPWR _24154_/Q sky130_fd_sc_hd__dfrtp_4
X_21366_ _21373_/A VGND VGND VPWR VPWR _21366_/X sky130_fd_sc_hd__buf_2
XANTENNA__18863__A2 _18834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14305__B _14305_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23105_ _23145_/CLK _23105_/D VGND VGND VPWR VPWR _15225_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20317_ _18759_/A _20317_/B VGND VGND VPWR VPWR _20317_/X sky130_fd_sc_hd__and2_4
XANTENNA__19384__A _19317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24085_ _24021_/CLK _20489_/X VGND VGND VPWR VPWR _24085_/Q sky130_fd_sc_hd__dfxtp_4
X_21297_ _21297_/A VGND VGND VPWR VPWR _21784_/C sky130_fd_sc_hd__buf_2
XANTENNA__16801__A _16616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23036_ _23036_/A VGND VGND VPWR VPWR HADDR[26] sky130_fd_sc_hd__inv_2
XFILLER_81_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21419__A _21419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20248_ _20248_/A _19926_/X VGND VGND VPWR VPWR _20301_/A sky130_fd_sc_hd__or2_4
XFILLER_7_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15417__A _13645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11945__A _11994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20179_ _19884_/X _18701_/X _20178_/X VGND VGND VPWR VPWR _20179_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_118_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14321__A _11911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_HCLK_A clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18379__B2 _18378_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18728__A _18728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22175__A2 _22172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14740_ _12883_/A _14811_/B VGND VGND VPWR VPWR _14740_/X sky130_fd_sc_hd__or2_4
XANTENNA__24275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11952_ _14880_/A VGND VGND VPWR VPWR _14906_/A sky130_fd_sc_hd__buf_2
X_23938_ _24066_/CLK _23938_/D VGND VGND VPWR VPWR _15283_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20186__A1 _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21154__A _21118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14671_ _14679_/A _23908_/Q VGND VGND VPWR VPWR _14671_/X sky130_fd_sc_hd__or2_4
X_11883_ _15784_/A VGND VGND VPWR VPWR _13427_/A sky130_fd_sc_hd__buf_2
X_23869_ _23867_/CLK _21356_/X VGND VGND VPWR VPWR _23869_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16248__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12776__A _12421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16410_ _11933_/X _16406_/X _16409_/X VGND VGND VPWR VPWR _16411_/B sky130_fd_sc_hd__or3_4
X_13622_ _13622_/A _24008_/Q VGND VGND VPWR VPWR _13624_/B sky130_fd_sc_hd__or2_4
XFILLER_73_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15152__A _14119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17390_ _17387_/X _17390_/B VGND VGND VPWR VPWR _17391_/A sky130_fd_sc_hd__and2_4
XANTENNA__21135__B1 _23986_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16341_ _16188_/A _16273_/B VGND VGND VPWR VPWR _16341_/X sky130_fd_sc_hd__or2_4
X_13553_ _12981_/A VGND VGND VPWR VPWR _13554_/A sky130_fd_sc_hd__buf_2
XFILLER_73_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14991__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12504_ _12518_/A _12614_/B VGND VGND VPWR VPWR _12506_/B sky130_fd_sc_hd__or2_4
X_19060_ _18935_/X VGND VGND VPWR VPWR _19060_/X sky130_fd_sc_hd__buf_2
X_16272_ _16243_/X _16272_/B VGND VGND VPWR VPWR _16272_/X sky130_fd_sc_hd__or2_4
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13484_ _12904_/A _13484_/B VGND VGND VPWR VPWR _13486_/B sky130_fd_sc_hd__or2_4
XFILLER_9_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15223_ _14215_/A _15221_/X _15222_/X VGND VGND VPWR VPWR _15224_/C sky130_fd_sc_hd__and3_4
X_18011_ _18174_/C VGND VGND VPWR VPWR _18011_/X sky130_fd_sc_hd__buf_2
XANTENNA__21438__A1 _21277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12435_ _12435_/A VGND VGND VPWR VPWR _15823_/A sky130_fd_sc_hd__buf_2
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21438__B2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17106__A2 _17032_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21989__A2 _21988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20217__B HRDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15154_ _11847_/A _15131_/X _15138_/X _15145_/X _15153_/X VGND VGND VPWR VPWR _15154_/X
+ sky130_fd_sc_hd__a32o_4
X_12366_ _11740_/A VGND VGND VPWR VPWR _12367_/A sky130_fd_sc_hd__buf_2
X_14105_ _15011_/A VGND VGND VPWR VPWR _14997_/A sky130_fd_sc_hd__buf_2
X_15085_ _14055_/A _15077_/X _15084_/X VGND VGND VPWR VPWR _15086_/C sky130_fd_sc_hd__and3_4
X_19962_ _24477_/Q VGND VGND VPWR VPWR _19962_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12297_ _15685_/A _12297_/B VGND VGND VPWR VPWR _12297_/X sky130_fd_sc_hd__or2_4
XFILLER_107_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12016__A _16541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16711__A _11982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14036_ _14065_/A _14036_/B _14036_/C VGND VGND VPWR VPWR _14036_/X sky130_fd_sc_hd__and3_4
X_18913_ _18877_/A VGND VGND VPWR VPWR _18913_/X sky130_fd_sc_hd__buf_2
X_19893_ _18752_/X VGND VGND VPWR VPWR _19893_/X sky130_fd_sc_hd__buf_2
XFILLER_49_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16430__B _16430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18844_ _15780_/B _18841_/X _24398_/Q _18842_/X VGND VGND VPWR VPWR _18844_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21610__B2 _21609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14231__A _14252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18775_ _18782_/A VGND VGND VPWR VPWR _18775_/X sky130_fd_sc_hd__buf_2
XFILLER_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15987_ _16095_/A _15987_/B _15987_/C VGND VGND VPWR VPWR _15987_/X sky130_fd_sc_hd__or3_4
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22166__A2 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17726_ _17726_/A VGND VGND VPWR VPWR _17726_/X sky130_fd_sc_hd__buf_2
XANTENNA__17542__A _16302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14938_ _13998_/A _14938_/B _14938_/C VGND VGND VPWR VPWR _14938_/X sky130_fd_sc_hd__and3_4
XANTENNA__21913__A2 _21908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21064__A _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17657_ _17651_/X _18003_/A VGND VGND VPWR VPWR _17765_/C sky130_fd_sc_hd__nor2_4
X_14869_ _13982_/A _14869_/B _14868_/X VGND VGND VPWR VPWR _14869_/X sky130_fd_sc_hd__and3_4
XFILLER_90_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12686__A _12284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18790__A1 _13575_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23332__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16608_ _16617_/A _16608_/B VGND VGND VPWR VPWR _16608_/X sky130_fd_sc_hd__or2_4
XANTENNA__24458__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21999__A _21985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17588_ _17508_/X _17587_/X _17501_/X _17510_/X VGND VGND VPWR VPWR _17589_/B sky130_fd_sc_hd__a211o_4
XFILLER_95_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19327_ _19325_/X _18226_/X _19325_/X _24244_/Q VGND VGND VPWR VPWR _19327_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15997__A _15997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16539_ _12024_/A VGND VGND VPWR VPWR _16565_/A sky130_fd_sc_hd__buf_2
XANTENNA__21677__B2 _21673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19258_ _24275_/Q _19223_/X _19257_/Y VGND VGND VPWR VPWR _19258_/X sky130_fd_sc_hd__o21a_4
XFILLER_108_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23482__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18209_ _18209_/A VGND VGND VPWR VPWR _18209_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21429__B2 _21423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19189_ _19115_/B VGND VGND VPWR VPWR _19189_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13310__A _12255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21220_ _21211_/Y _21218_/X _21219_/X _21218_/X VGND VGND VPWR VPWR _21220_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21151_ _21130_/A VGND VGND VPWR VPWR _21151_/X sky130_fd_sc_hd__buf_2
XANTENNA__16621__A _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20102_ _11569_/X _20090_/D VGND VGND VPWR VPWR _20134_/A sky130_fd_sc_hd__or2_4
X_21082_ _21075_/A VGND VGND VPWR VPWR _21082_/X sky130_fd_sc_hd__buf_2
XANTENNA__21239__A _20464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16340__B _16272_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20033_ _19985_/A VGND VGND VPWR VPWR _20033_/X sky130_fd_sc_hd__buf_2
XANTENNA__11765__A _14020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15237__A _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21601__B2 _21595_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19558__B1 HRDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17452__A _17181_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21984_ _21809_/X _21981_/X _12213_/B _21978_/X VGND VGND VPWR VPWR _21984_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21904__A2 _21901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23723_ _24011_/CLK _23723_/D VGND VGND VPWR VPWR _23723_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_76_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20935_ _24194_/Q _20873_/X _20934_/Y VGND VGND VPWR VPWR _22456_/A sky130_fd_sc_hd__o21a_4
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12596__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _23845_/CLK _23654_/D VGND VGND VPWR VPWR _14283_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _24229_/Q _20639_/X _20865_/X VGND VGND VPWR VPWR _20866_/X sky130_fd_sc_hd__o21a_4
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22605_ _22446_/X _22600_/X _14373_/B _22604_/X VGND VGND VPWR VPWR _23142_/D sky130_fd_sc_hd__o22a_4
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21702__A _21702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21668__B2 _21666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23585_ _23391_/CLK _23585_/D VGND VGND VPWR VPWR _23585_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20797_ _21843_/A VGND VGND VPWR VPWR _20797_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15700__A _12739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22536_ _22536_/A VGND VGND VPWR VPWR _22536_/X sky130_fd_sc_hd__buf_2
XANTENNA__16515__B _16514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20891__A2 _20873_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22467_ _22471_/A VGND VGND VPWR VPWR _22483_/A sky130_fd_sc_hd__inv_2
XFILLER_13_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12220_ _13054_/A VGND VGND VPWR VPWR _12688_/A sky130_fd_sc_hd__buf_2
X_24206_ _24208_/CLK _19393_/X HRESETn VGND VGND VPWR VPWR _24206_/Q sky130_fd_sc_hd__dfrtp_4
X_21418_ _21244_/X _21412_/X _23828_/Q _21416_/X VGND VGND VPWR VPWR _23828_/D sky130_fd_sc_hd__o22a_4
X_22398_ _20372_/A VGND VGND VPWR VPWR _22398_/X sky130_fd_sc_hd__buf_2
XANTENNA__22533__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12151_ _16045_/A _12135_/X _12150_/X VGND VGND VPWR VPWR _12183_/B sky130_fd_sc_hd__or3_4
X_24137_ _24473_/CLK _24137_/D HRESETn VGND VGND VPWR VPWR _16939_/A sky130_fd_sc_hd__dfrtp_4
X_21349_ _21348_/X VGND VGND VPWR VPWR _21383_/A sky130_fd_sc_hd__buf_2
XANTENNA__16531__A _16536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18049__B1 _18048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12082_ _12036_/X _12050_/X _12061_/X _12073_/X _12081_/X VGND VGND VPWR VPWR _12082_/X
+ sky130_fd_sc_hd__a32o_4
X_24068_ _23363_/CLK _24068_/D VGND VGND VPWR VPWR _24068_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23042__B1 _17944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11675__A _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15910_ _15844_/X VGND VGND VPWR VPWR _15910_/Y sky130_fd_sc_hd__inv_2
X_23019_ _23014_/X _17661_/A _22997_/X _23018_/X VGND VGND VPWR VPWR _23020_/A sky130_fd_sc_hd__a211o_4
XANTENNA__15147__A _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16890_ _16821_/X _16890_/B VGND VGND VPWR VPWR _16890_/X sky130_fd_sc_hd__and2_4
X_15841_ _13041_/A _15837_/X _15841_/C VGND VGND VPWR VPWR _15842_/B sky130_fd_sc_hd__or3_4
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18458__A _18171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14986__A _11652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22148__A2 _22101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13890__A _13890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18560_ _22927_/B _18559_/Y _16998_/A _18558_/X VGND VGND VPWR VPWR _18560_/X sky130_fd_sc_hd__o22a_4
X_12984_ _12622_/X _12912_/B VGND VGND VPWR VPWR _12984_/X sky130_fd_sc_hd__or2_4
X_15772_ _12792_/A _15699_/B VGND VGND VPWR VPWR _15772_/X sky130_fd_sc_hd__or2_4
XANTENNA__21356__B1 _23869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17511_ _18297_/B _17510_/X VGND VGND VPWR VPWR _17512_/A sky130_fd_sc_hd__or2_4
XANTENNA__18221__B1 _18160_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11935_ _16121_/A VGND VGND VPWR VPWR _16130_/A sky130_fd_sc_hd__buf_2
X_14723_ _14640_/X _14723_/B VGND VGND VPWR VPWR _14724_/B sky130_fd_sc_hd__and2_4
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18491_ _17422_/B _18538_/A _17425_/X VGND VGND VPWR VPWR _18491_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18772__A1 _17277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14654_ _14672_/A _14654_/B VGND VGND VPWR VPWR _14655_/C sky130_fd_sc_hd__or2_4
X_17442_ _17442_/A VGND VGND VPWR VPWR _17667_/B sky130_fd_sc_hd__inv_2
X_11866_ _13955_/A VGND VGND VPWR VPWR _13968_/A sky130_fd_sc_hd__buf_2
XANTENNA__21108__B1 _14866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13605_ _13959_/A VGND VGND VPWR VPWR _13606_/A sky130_fd_sc_hd__buf_2
XANTENNA__21612__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14585_ _14152_/A _14667_/B VGND VGND VPWR VPWR _14586_/C sky130_fd_sc_hd__or2_4
X_17373_ _17372_/X VGND VGND VPWR VPWR _18405_/A sky130_fd_sc_hd__inv_2
XFILLER_57_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22856__B1 _17383_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11797_ _11797_/A VGND VGND VPWR VPWR _11798_/A sky130_fd_sc_hd__buf_2
XFILLER_57_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16706__A _12025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19112_ _19112_/A _19112_/B VGND VGND VPWR VPWR _19112_/X sky130_fd_sc_hd__and2_4
X_13536_ _13494_/X _13536_/B _13536_/C VGND VGND VPWR VPWR _13537_/C sky130_fd_sc_hd__or3_4
X_16324_ _16366_/A _16322_/X _16324_/C VGND VGND VPWR VPWR _16330_/B sky130_fd_sc_hd__and3_4
XFILLER_43_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13349__B1 _11596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16255_ _15980_/A _16250_/X _16254_/X VGND VGND VPWR VPWR _16255_/X sky130_fd_sc_hd__or3_4
X_19043_ _19041_/Y _19042_/Y _11517_/B VGND VGND VPWR VPWR _19043_/X sky130_fd_sc_hd__o21a_4
X_13467_ _13467_/A _13467_/B _13467_/C VGND VGND VPWR VPWR _13468_/C sky130_fd_sc_hd__and3_4
X_15206_ _14246_/A _15204_/X _15206_/C VGND VGND VPWR VPWR _15207_/C sky130_fd_sc_hd__and3_4
XANTENNA__13130__A _13130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12418_ _12418_/A _12312_/B VGND VGND VPWR VPWR _12420_/B sky130_fd_sc_hd__or2_4
X_16186_ _16219_/A _16186_/B VGND VGND VPWR VPWR _16186_/X sky130_fd_sc_hd__or2_4
XANTENNA__11569__B IRQ[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13398_ _13397_/X _24048_/Q VGND VGND VPWR VPWR _13398_/X sky130_fd_sc_hd__or2_4
XANTENNA__20095__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15137_ _14098_/A _15135_/X _15136_/X VGND VGND VPWR VPWR _15137_/X sky130_fd_sc_hd__and3_4
X_12349_ _12412_/A VGND VGND VPWR VPWR _12350_/A sky130_fd_sc_hd__buf_2
XANTENNA__17537__A _17144_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16441__A _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15068_ _14071_/A _15068_/B _15068_/C VGND VGND VPWR VPWR _15086_/B sky130_fd_sc_hd__and3_4
X_19945_ _19945_/A VGND VGND VPWR VPWR _19945_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21059__A _21007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14019_ _14071_/A _14019_/B _14019_/C VGND VGND VPWR VPWR _14019_/X sky130_fd_sc_hd__and3_4
XFILLER_64_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19876_ _19793_/A _19876_/B VGND VGND VPWR VPWR _19876_/X sky130_fd_sc_hd__or2_4
XFILLER_64_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24126__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18827_ _18834_/A VGND VGND VPWR VPWR _18827_/X sky130_fd_sc_hd__buf_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18758_ _18757_/X VGND VGND VPWR VPWR _18759_/A sky130_fd_sc_hd__buf_2
XFILLER_55_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17709_ _17708_/X VGND VGND VPWR VPWR _17749_/B sky130_fd_sc_hd__inv_2
XFILLER_64_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23848__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18689_ _24450_/Q VGND VGND VPWR VPWR _18689_/Y sky130_fd_sc_hd__inv_2
X_20720_ _20534_/A _20719_/X VGND VGND VPWR VPWR _20720_/X sky130_fd_sc_hd__or2_4
XANTENNA__13305__A _13428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22618__A _22633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18815__B _18814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21522__A _20442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20651_ _20642_/X _20647_/X _20650_/X VGND VGND VPWR VPWR _20651_/X sky130_fd_sc_hd__and3_4
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16616__A _16616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23370_ _23978_/CLK _22235_/X VGND VGND VPWR VPWR _13969_/B sky130_fd_sc_hd__dfxtp_4
X_20582_ _20494_/X _20581_/X _24336_/Q _20453_/X VGND VGND VPWR VPWR _20582_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20138__A IRQ[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22321_ _14217_/B VGND VGND VPWR VPWR _23305_/D sky130_fd_sc_hd__buf_2
XFILLER_20_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14136__A _14136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13040__A _13017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22252_ _22251_/X VGND VGND VPWR VPWR _22286_/A sky130_fd_sc_hd__buf_2
XFILLER_118_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21203_ _20870_/X _21197_/X _14533_/B _21201_/X VGND VGND VPWR VPWR _23941_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13975__A _12217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22183_ _22169_/A VGND VGND VPWR VPWR _22183_/X sky130_fd_sc_hd__buf_2
XANTENNA__21822__B2 _21812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16351__A _16365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21134_ _20537_/X _21133_/X _23987_/Q _21130_/X VGND VGND VPWR VPWR _21134_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22378__A2 _22375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19779__B1 _19592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23378__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21065_ _21072_/A VGND VGND VPWR VPWR _21065_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20016_ _19994_/X _17672_/A _20000_/X _20015_/X VGND VGND VPWR VPWR _20017_/A sky130_fd_sc_hd__o22a_4
XFILLER_8_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21050__A2 _21044_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12103__B _23645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17182__A _17181_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21338__B1 _14301_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15414__B _15471_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21967_ _21684_/A _21634_/B _21684_/C _21008_/A VGND VGND VPWR VPWR _21967_/X sky130_fd_sc_hd__or4_4
XANTENNA__21889__B2 _21884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18754__A1 _17736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _13688_/A VGND VGND VPWR VPWR _13708_/A sky130_fd_sc_hd__inv_2
X_23706_ _23706_/CLK _21646_/X VGND VGND VPWR VPWR _16437_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ _20844_/A _20539_/B VGND VGND VPWR VPWR _20918_/X sky130_fd_sc_hd__or2_4
XFILLER_70_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ _21884_/A VGND VGND VPWR VPWR _21898_/X sky130_fd_sc_hd__buf_2
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11651_/A _13991_/A VGND VGND VPWR VPWR _11652_/D sky130_fd_sc_hd__or2_4
X_23637_ _24021_/CLK _23637_/D VGND VGND VPWR VPWR _12668_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ _20644_/A _20849_/B VGND VGND VPWR VPWR _20849_/X sky130_fd_sc_hd__and2_4
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16526__A _12022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15430__A _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _15616_/A _14368_/X _14370_/C VGND VGND VPWR VPWR _14377_/B sky130_fd_sc_hd__and3_4
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ _16919_/A VGND VGND VPWR VPWR _17024_/C sky130_fd_sc_hd__buf_2
X_23568_ _24047_/CLK _21892_/X VGND VGND VPWR VPWR _23568_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20048__A _20000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _13286_/X _23600_/Q VGND VGND VPWR VPWR _13321_/X sky130_fd_sc_hd__or2_4
XFILLER_70_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22519_ _22518_/X VGND VGND VPWR VPWR _22519_/X sky130_fd_sc_hd__buf_2
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19837__A _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23499_ _23915_/CLK _22000_/X VGND VGND VPWR VPWR _23499_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14046__A _14046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16040_ _16064_/A _15960_/B VGND VGND VPWR VPWR _16040_/X sky130_fd_sc_hd__or2_4
XFILLER_109_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13252_ _15484_/A _13252_/B _13252_/C VGND VGND VPWR VPWR _13268_/B sky130_fd_sc_hd__and3_4
XFILLER_108_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18809__A2 _18781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24153__CLK _24162_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12203_ _12203_/A VGND VGND VPWR VPWR _15432_/A sky130_fd_sc_hd__buf_2
X_13183_ _12737_/A _13181_/X _13182_/X VGND VGND VPWR VPWR _13183_/X sky130_fd_sc_hd__and3_4
XANTENNA__21813__B2 _21812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12134_ _11746_/X _12130_/X _12134_/C VGND VGND VPWR VPWR _12134_/X sky130_fd_sc_hd__or3_4
X_17991_ _18024_/B _17990_/X VGND VGND VPWR VPWR _17991_/X sky130_fd_sc_hd__or2_4
XFILLER_96_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22369__A2 _22368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19730_ _19730_/A _19818_/A _19861_/A _19730_/D VGND VGND VPWR VPWR _19730_/X sky130_fd_sc_hd__or4_4
XFILLER_46_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12065_ _11994_/A VGND VGND VPWR VPWR _12065_/X sky130_fd_sc_hd__buf_2
X_16942_ _17652_/A VGND VGND VPWR VPWR _16942_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19661_ _19661_/A _19661_/B VGND VGND VPWR VPWR _19662_/A sky130_fd_sc_hd__or2_4
X_16873_ _16850_/A _16850_/B VGND VGND VPWR VPWR _16876_/C sky130_fd_sc_hd__nand2_4
XFILLER_65_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20511__A _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18612_ _18611_/X VGND VGND VPWR VPWR _18612_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17092__A _17057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15824_ _12518_/X _15824_/B VGND VGND VPWR VPWR _15826_/B sky130_fd_sc_hd__or2_4
X_19592_ _19592_/A _19582_/Y VGND VGND VPWR VPWR _19592_/X sky130_fd_sc_hd__and2_4
XANTENNA__13806__A1 _13682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12948__B _12948_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18543_ _17794_/X _18186_/Y _17856_/X _18542_/X VGND VGND VPWR VPWR _18543_/X sky130_fd_sc_hd__a211o_4
XFILLER_79_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_54_0_HCLK clkbuf_7_54_0_HCLK/A VGND VGND VPWR VPWR _23404_/CLK sky130_fd_sc_hd__clkbuf_1
X_12967_ _12967_/A _12965_/X _12967_/C VGND VGND VPWR VPWR _12967_/X sky130_fd_sc_hd__and3_4
X_15755_ _15725_/A _15690_/B VGND VGND VPWR VPWR _15755_/X sky130_fd_sc_hd__or2_4
XFILLER_80_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22541__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11918_ _11886_/X VGND VGND VPWR VPWR _11983_/A sky130_fd_sc_hd__buf_2
X_14706_ _14341_/A _14706_/B VGND VGND VPWR VPWR _14708_/B sky130_fd_sc_hd__or2_4
X_18474_ _17382_/A _18473_/B _18048_/A VGND VGND VPWR VPWR _18474_/Y sky130_fd_sc_hd__a21oi_4
X_12898_ _12520_/X _24051_/Q VGND VGND VPWR VPWR _12899_/C sky130_fd_sc_hd__or2_4
X_15686_ _12722_/A _15686_/B VGND VGND VPWR VPWR _15687_/C sky130_fd_sc_hd__or2_4
X_17425_ _17179_/Y _17396_/Y VGND VGND VPWR VPWR _17425_/X sky130_fd_sc_hd__or2_4
XFILLER_33_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11849_ _13056_/A VGND VGND VPWR VPWR _11850_/A sky130_fd_sc_hd__buf_2
X_14637_ _14782_/A _14633_/X _14637_/C VGND VGND VPWR VPWR _14637_/X sky130_fd_sc_hd__or3_4
XFILLER_92_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12964__A _12964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16436__A _11872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14568_ _14567_/X VGND VGND VPWR VPWR _14568_/Y sky130_fd_sc_hd__inv_2
X_17356_ _17192_/Y _17356_/B VGND VGND VPWR VPWR _17356_/X sky130_fd_sc_hd__or2_4
XANTENNA__20304__A1 _20293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21061__B _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12683__B _12758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16307_ _12830_/A VGND VGND VPWR VPWR _16366_/A sky130_fd_sc_hd__buf_2
XFILLER_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13519_ _12596_/A VGND VGND VPWR VPWR _13522_/A sky130_fd_sc_hd__buf_2
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19747__A HRDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14499_ _14499_/A VGND VGND VPWR VPWR _14556_/A sky130_fd_sc_hd__buf_2
X_17287_ _17287_/A _17413_/B VGND VGND VPWR VPWR _17287_/X sky130_fd_sc_hd__or2_4
XFILLER_70_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19026_ _24366_/Q VGND VGND VPWR VPWR _19026_/Y sky130_fd_sc_hd__inv_2
X_16238_ _16155_/X _16235_/X _16237_/Y VGND VGND VPWR VPWR _16239_/B sky130_fd_sc_hd__a21o_4
XANTENNA__22057__B2 _22056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13795__A _13630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20607__A2 _20421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17267__A _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16169_ _13388_/A VGND VGND VPWR VPWR _16203_/A sky130_fd_sc_hd__buf_2
XFILLER_66_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24307__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19928_ _19927_/X VGND VGND VPWR VPWR _19996_/A sky130_fd_sc_hd__buf_2
XFILLER_69_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19482__A _19598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12204__A _15432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21032__A2 _21030_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21517__A _21802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19859_ _19534_/X _19622_/A _19854_/X _19858_/X VGND VGND VPWR VPWR _19859_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20421__A _20421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15515__A _11671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22870_ _22854_/X _22810_/X _17339_/Y _22855_/X VGND VGND VPWR VPWR _22870_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20791__A1 _18548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21821_ _20574_/A VGND VGND VPWR VPWR _21821_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15234__B _15177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22532__A2 _22529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13035__A _12915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21752_ _21752_/A VGND VGND VPWR VPWR _21752_/X sky130_fd_sc_hd__buf_2
XFILLER_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20543__B2 _20497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20703_ _20467_/A VGND VGND VPWR VPWR _20715_/A sky130_fd_sc_hd__buf_2
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24471_ _24241_/CLK _24471_/D HRESETn VGND VGND VPWR VPWR _19990_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21683_ _21683_/A VGND VGND VPWR VPWR _21683_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16346__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23422_ _23326_/CLK _22156_/X VGND VGND VPWR VPWR _11814_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15250__A _15249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20634_ _20634_/A _20634_/B VGND VGND VPWR VPWR _20634_/Y sky130_fd_sc_hd__nand2_4
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21099__A2 _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22296__B2 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23353_ _23354_/CLK _23353_/D VGND VGND VPWR VPWR _16244_/B sky130_fd_sc_hd__dfxtp_4
X_20565_ _20517_/X _20564_/X _24305_/Q _20527_/X VGND VGND VPWR VPWR _20566_/B sky130_fd_sc_hd__o22a_4
X_22304_ _22304_/A VGND VGND VPWR VPWR _23322_/D sky130_fd_sc_hd__buf_2
XFILLER_109_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22048__B2 _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23284_ _23157_/CLK _23284_/D VGND VGND VPWR VPWR _12784_/B sky130_fd_sc_hd__dfxtp_4
X_20496_ _20448_/X _20495_/X _24372_/Q _20407_/X VGND VGND VPWR VPWR _20496_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22083__A _20372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22599__A2 _22593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22235_ _22122_/X _22229_/X _13969_/B _22233_/X VGND VGND VPWR VPWR _22235_/X sky130_fd_sc_hd__o22a_4
X_22166_ _22088_/X _22165_/X _23416_/Q _22162_/X VGND VGND VPWR VPWR _23416_/D sky130_fd_sc_hd__o22a_4
X_21117_ _21110_/Y _21116_/X _20277_/X _21116_/X VGND VGND VPWR VPWR _23998_/D sky130_fd_sc_hd__a2bb2o_4
X_22097_ _22095_/X _22089_/X _12623_/B _22096_/X VGND VGND VPWR VPWR _23445_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21559__B1 _13713_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21048_ _21027_/A VGND VGND VPWR VPWR _21048_/X sky130_fd_sc_hd__buf_2
XFILLER_82_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22220__B2 _22219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15425__A _15429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11953__A _14906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13870_ _14178_/A VGND VGND VPWR VPWR _13871_/A sky130_fd_sc_hd__buf_2
XFILLER_41_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23064__D _23062_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12768__B _12768_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12821_ _12753_/X _12821_/B _12821_/C VGND VGND VPWR VPWR _12821_/X sky130_fd_sc_hd__or3_4
X_22999_ _18256_/X _23004_/B VGND VGND VPWR VPWR _23000_/C sky130_fd_sc_hd__or2_4
XFILLER_43_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14461__A1 _13056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22523__A2 _22522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20985__B _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12752_ _12751_/X VGND VGND VPWR VPWR _12752_/Y sky130_fd_sc_hd__inv_2
X_15540_ _14432_/A _23531_/Q VGND VGND VPWR VPWR _15541_/C sky130_fd_sc_hd__or2_4
XFILLER_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22258__A _22272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _16023_/A VGND VGND VPWR VPWR _16071_/A sky130_fd_sc_hd__buf_2
XFILLER_76_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _12585_/A _15471_/B VGND VGND VPWR VPWR _15471_/X sky130_fd_sc_hd__or2_4
X_12683_ _12553_/A _12758_/B VGND VGND VPWR VPWR _12685_/B sky130_fd_sc_hd__or2_4
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14040_/X _14422_/B _14422_/C VGND VGND VPWR VPWR _14422_/X sky130_fd_sc_hd__or3_4
X_17210_ _16235_/X _17131_/X _14429_/B _17186_/X VGND VGND VPWR VPWR _17210_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15160__A _14098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11634_/A _11634_/B _17009_/A _17285_/A VGND VGND VPWR VPWR _11634_/X sky130_fd_sc_hd__or4_4
XANTENNA__18174__C _18174_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18190_ _18425_/A _18156_/X _18189_/X _18151_/X VGND VGND VPWR VPWR _18190_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22287__B2 _22283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14353_ _14345_/A VGND VGND VPWR VPWR _15592_/A sky130_fd_sc_hd__buf_2
X_17141_ _17130_/A VGND VGND VPWR VPWR _17141_/X sky130_fd_sc_hd__buf_2
XFILLER_89_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _24440_/Q IRQ[25] _11564_/X VGND VGND VPWR VPWR _11565_/X sky130_fd_sc_hd__a21o_4
XFILLER_106_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13304_ _13300_/A _13304_/B VGND VGND VPWR VPWR _13304_/X sky130_fd_sc_hd__or2_4
XFILLER_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23543__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17072_ _17072_/A _18750_/A _17082_/B VGND VGND VPWR VPWR _17073_/B sky130_fd_sc_hd__or3_4
XANTENNA__22039__A1 _21816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14284_ _15533_/A _14379_/B VGND VGND VPWR VPWR _14284_/X sky130_fd_sc_hd__or2_4
XANTENNA__22039__B2 _22035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13235_ _13211_/A _13235_/B _13235_/C VGND VGND VPWR VPWR _13236_/C sky130_fd_sc_hd__or3_4
X_16023_ _16023_/A VGND VGND VPWR VPWR _16037_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14504__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24400__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13166_ _12315_/A _13166_/B VGND VGND VPWR VPWR _13166_/X sky130_fd_sc_hd__or2_4
XANTENNA__18663__B1 _17634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21262__A2 _21259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15319__B _15256_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12117_ _16071_/A VGND VGND VPWR VPWR _12152_/A sky130_fd_sc_hd__buf_2
XFILLER_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13097_ _13097_/A VGND VGND VPWR VPWR _13100_/A sky130_fd_sc_hd__buf_2
X_17974_ _17921_/X _17971_/Y _17800_/X _17973_/Y VGND VGND VPWR VPWR _17974_/X sky130_fd_sc_hd__o22a_4
XFILLER_97_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12024__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17218__A1 _17007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19713_ _20490_/B _19551_/X _19712_/X _19616_/X VGND VGND VPWR VPWR _19713_/X sky130_fd_sc_hd__a211o_4
X_12048_ _16698_/A _23741_/Q VGND VGND VPWR VPWR _12049_/C sky130_fd_sc_hd__or2_4
X_16925_ _16924_/X VGND VGND VPWR VPWR _16925_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21337__A _21316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22211__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12959__A _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20241__A _20447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19644_ _19640_/X _19806_/C _19481_/A VGND VGND VPWR VPWR _19644_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__24049__CLK _23155_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15335__A _14000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16856_ _16840_/C _16840_/B _16840_/C _16840_/B VGND VGND VPWR VPWR _16870_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18430__A3 _18426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15807_ _11912_/A _15807_/B _15806_/X VGND VGND VPWR VPWR _15807_/X sky130_fd_sc_hd__and3_4
XFILLER_53_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19575_ _19629_/A _19706_/A _19629_/B VGND VGND VPWR VPWR _19575_/X sky130_fd_sc_hd__o21a_4
X_16787_ _11834_/A _16783_/X _16787_/C VGND VGND VPWR VPWR _16787_/X sky130_fd_sc_hd__or3_4
XFILLER_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13999_ _11645_/A VGND VGND VPWR VPWR _14000_/A sky130_fd_sc_hd__buf_2
XFILLER_81_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20895__B _20895_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18526_ _17418_/X _18524_/X _18063_/A _18525_/X VGND VGND VPWR VPWR _18527_/A sky130_fd_sc_hd__a211o_4
XFILLER_46_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15738_ _12794_/A VGND VGND VPWR VPWR _15751_/A sky130_fd_sc_hd__buf_2
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21072__A _21072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19391__B2 _24207_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18457_ _18435_/X _18456_/X _20043_/A _18435_/X VGND VGND VPWR VPWR _18457_/X sky130_fd_sc_hd__a2bb2o_4
X_15669_ _12735_/A _15669_/B VGND VGND VPWR VPWR _15669_/X sky130_fd_sc_hd__or2_4
XFILLER_21_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12694__A _12240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17941__A2 _17577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17408_ _17407_/X VGND VGND VPWR VPWR _17408_/Y sky130_fd_sc_hd__inv_2
X_18388_ _18265_/A _17371_/X VGND VGND VPWR VPWR _18390_/C sky130_fd_sc_hd__nor2_4
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22278__B2 _22276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21800__A _21787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17339_ _15582_/X VGND VGND VPWR VPWR _17339_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18381__A _18381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20350_ _17944_/X _20238_/X _20319_/X _20349_/Y VGND VGND VPWR VPWR _20350_/X sky130_fd_sc_hd__a211o_4
XANTENNA__18812__C _18812_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19009_ _19007_/Y _19008_/Y _11522_/X VGND VGND VPWR VPWR _19009_/X sky130_fd_sc_hd__o21a_4
X_20281_ _20399_/A VGND VGND VPWR VPWR _20282_/A sky130_fd_sc_hd__buf_2
X_22020_ _22035_/A VGND VGND VPWR VPWR _22020_/X sky130_fd_sc_hd__buf_2
XANTENNA__18654__B1 _17742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24141__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22450__B2 _22447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17209__A1 _17156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18406__B1 _18160_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21247__A _21247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23971_ _23270_/CLK _23971_/D VGND VGND VPWR VPWR _14811_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_9_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12869__A _12477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22922_ _18593_/X _22908_/Y _22924_/A _22921_/X VGND VGND VPWR VPWR _22923_/C sky130_fd_sc_hd__a211o_4
XFILLER_60_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19940__A _18062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15245__A _14246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12588__B _12572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22853_ _19887_/X VGND VGND VPWR VPWR _22853_/X sky130_fd_sc_hd__buf_2
XFILLER_71_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18556__A _24190_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22505__A2 _22500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21804_ _21804_/A VGND VGND VPWR VPWR _21804_/X sky130_fd_sc_hd__buf_2
X_22784_ _15120_/Y _22782_/X VGND VGND VPWR VPWR HWDATA[1] sky130_fd_sc_hd__nor2_4
XANTENNA__15899__B _15829_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21735_ _21734_/X VGND VGND VPWR VPWR _21740_/A sky130_fd_sc_hd__buf_2
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16076__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23566__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24454_ _24202_/CLK _24454_/D HRESETn VGND VGND VPWR VPWR _20079_/A sky130_fd_sc_hd__dfrtp_4
X_21666_ _21659_/A VGND VGND VPWR VPWR _21666_/X sky130_fd_sc_hd__buf_2
XFILLER_71_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23405_ _23314_/CLK _22181_/X VGND VGND VPWR VPWR _15825_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14308__B _14308_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20617_ _20616_/X VGND VGND VPWR VPWR _20617_/X sky130_fd_sc_hd__buf_2
XFILLER_36_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24385_ _24425_/CLK _18861_/X HRESETn VGND VGND VPWR VPWR _24385_/Q sky130_fd_sc_hd__dfrtp_4
X_21597_ _21517_/X _21591_/X _16245_/B _21595_/X VGND VGND VPWR VPWR _21597_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18291__A _18129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23336_ _23336_/CLK _22288_/X VGND VGND VPWR VPWR _13702_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20548_ _24242_/Q VGND VGND VPWR VPWR _20548_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21492__A2 _21491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11948__A _16113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23267_ _23907_/CLK _23267_/D VGND VGND VPWR VPWR _14798_/B sky130_fd_sc_hd__dfxtp_4
X_20479_ _20603_/A _20479_/B VGND VGND VPWR VPWR _20479_/Y sky130_fd_sc_hd__nor2_4
XFILLER_84_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13020_ _13020_/A _13085_/B VGND VGND VPWR VPWR _13021_/C sky130_fd_sc_hd__or2_4
X_22218_ _22093_/X _22215_/X _12297_/B _22212_/X VGND VGND VPWR VPWR _22218_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15139__B _23649_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23198_ _23326_/CLK _22520_/X VGND VGND VPWR VPWR _11749_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22441__B2 _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22149_ _11814_/B VGND VGND VPWR VPWR _22149_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14978__B _14903_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14971_ _14937_/A _23776_/Q VGND VGND VPWR VPWR _14972_/C sky130_fd_sc_hd__or2_4
XFILLER_43_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16710_ _11936_/X _16710_/B _16709_/X VGND VGND VPWR VPWR _16711_/B sky130_fd_sc_hd__or3_4
XANTENNA__11683__A _13415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13922_ _13922_/A VGND VGND VPWR VPWR _13922_/Y sky130_fd_sc_hd__inv_2
X_17690_ _17690_/A VGND VGND VPWR VPWR _17690_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16641_ _16630_/X _16550_/B VGND VGND VPWR VPWR _16641_/X sky130_fd_sc_hd__or2_4
X_13853_ _13911_/A _13848_/X _13852_/X VGND VGND VPWR VPWR _13854_/C sky130_fd_sc_hd__and3_4
XANTENNA__14994__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17370__A _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12804_ _12769_/A _12804_/B _12804_/C VGND VGND VPWR VPWR _12805_/C sky130_fd_sc_hd__and3_4
X_19360_ _19355_/X _18754_/Y _19359_/X _20997_/A VGND VGND VPWR VPWR _24223_/D sky130_fd_sc_hd__a2bb2o_4
X_16572_ _16565_/A _23836_/Q VGND VGND VPWR VPWR _16573_/C sky130_fd_sc_hd__or2_4
XANTENNA__20507__A1 _24212_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13784_ _15399_/A _13784_/B VGND VGND VPWR VPWR _13784_/X sky130_fd_sc_hd__or2_4
XFILLER_56_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18311_ _17678_/X _18286_/X _17678_/X _18286_/X VGND VGND VPWR VPWR _18311_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15523_ _12238_/X _23499_/Q VGND VGND VPWR VPWR _15523_/X sky130_fd_sc_hd__or2_4
X_12735_ _12735_/A _12735_/B VGND VGND VPWR VPWR _12735_/X sky130_fd_sc_hd__or2_4
X_19291_ _19208_/B VGND VGND VPWR VPWR _19291_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15602__B _23435_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17923__A2 _17919_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18242_ _18242_/A _17446_/X VGND VGND VPWR VPWR _18244_/C sky130_fd_sc_hd__nor2_4
X_12666_ _12970_/A _12664_/X _12666_/C VGND VGND VPWR VPWR _12670_/B sky130_fd_sc_hd__and3_4
X_15454_ _15486_/A _15454_/B VGND VGND VPWR VPWR _15454_/X sky130_fd_sc_hd__or2_4
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22716__A _22932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _13595_/A VGND VGND VPWR VPWR _11618_/A sky130_fd_sc_hd__buf_2
X_14405_ _15628_/A _14397_/X _14404_/X VGND VGND VPWR VPWR _14422_/B sky130_fd_sc_hd__and3_4
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18173_ _16981_/X VGND VGND VPWR VPWR _18174_/B sky130_fd_sc_hd__inv_2
XANTENNA__19297__A _20190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _14177_/A VGND VGND VPWR VPWR _12598_/A sky130_fd_sc_hd__buf_2
X_15385_ _15185_/X _15251_/X _15382_/X _15384_/Y VGND VGND VPWR VPWR _15385_/X sky130_fd_sc_hd__a211o_4
XANTENNA__19676__A2 _19674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ _17160_/A VGND VGND VPWR VPWR _17220_/A sky130_fd_sc_hd__inv_2
XFILLER_106_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11548_ _11539_/X _11540_/X _11542_/X _20071_/B VGND VGND VPWR VPWR _11548_/X sky130_fd_sc_hd__or4_4
X_14336_ _13594_/X _13595_/X _14300_/X _11595_/A _14335_/X VGND VGND VPWR VPWR _14336_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21483__A2 _21477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22680__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11858__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14267_ _14077_/X _14267_/B VGND VGND VPWR VPWR _14267_/X sky130_fd_sc_hd__or2_4
X_17055_ _11584_/A VGND VGND VPWR VPWR _20206_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13218_ _12367_/A _13214_/X _13218_/C VGND VGND VPWR VPWR _13219_/C sky130_fd_sc_hd__or3_4
X_16006_ _11982_/A _15980_/X _15987_/X _15995_/X _16005_/X VGND VGND VPWR VPWR _16006_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_28_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14198_ _14204_/A _24009_/Q VGND VGND VPWR VPWR _14200_/B sky130_fd_sc_hd__or2_4
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22451__A _20892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13149_ _15667_/A _13149_/B VGND VGND VPWR VPWR _13149_/X sky130_fd_sc_hd__or2_4
XFILLER_44_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17545__A _17544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22983__A2 _17681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20994__A1 _20493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14888__B _23872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21067__A _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17957_ _18265_/A _17957_/B VGND VGND VPWR VPWR _17959_/C sky130_fd_sc_hd__nor2_4
XFILLER_39_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12689__A _12556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16908_ _17052_/A VGND VGND VPWR VPWR _16910_/A sky130_fd_sc_hd__inv_2
X_17888_ _18129_/A VGND VGND VPWR VPWR _17888_/X sky130_fd_sc_hd__buf_2
XFILLER_22_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20746__A1 _24202_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24368__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19627_ _19637_/A _19626_/X VGND VGND VPWR VPWR _19627_/Y sky130_fd_sc_hd__nor2_4
X_16839_ _15914_/D _16838_/X _15914_/D _16838_/X VGND VGND VPWR VPWR _16839_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19558_ _19422_/X _19557_/X HRDATA[9] _19438_/X VGND VGND VPWR VPWR _19559_/A sky130_fd_sc_hd__o22a_4
XFILLER_59_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22499__B2 _22497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_24_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_24_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18509_ _17748_/X _17710_/X _17708_/X VGND VGND VPWR VPWR _18509_/X sky130_fd_sc_hd__o21a_4
XFILLER_62_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19489_ _19536_/A _19481_/X _19537_/A VGND VGND VPWR VPWR _19489_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21171__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21520_ _21532_/A VGND VGND VPWR VPWR _21520_/X sky130_fd_sc_hd__buf_2
XANTENNA__13313__A _12740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22626__A _22626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21451_ _21455_/A VGND VGND VPWR VPWR _21467_/A sky130_fd_sc_hd__inv_2
XFILLER_33_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24393__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16624__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20402_ _20468_/A VGND VGND VPWR VPWR _20403_/A sky130_fd_sc_hd__buf_2
XANTENNA__17678__A1 _17674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24170_ _24293_/CLK _19816_/X HRESETn VGND VGND VPWR VPWR _16893_/A sky130_fd_sc_hd__dfrtp_4
X_21382_ _21268_/X _21376_/X _23850_/Q _21380_/X VGND VGND VPWR VPWR _23850_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20146__A IRQ[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23121_ _23217_/CLK _23121_/D VGND VGND VPWR VPWR _13178_/B sky130_fd_sc_hd__dfxtp_4
X_20333_ _17880_/X _20238_/X _20319_/X _20332_/Y VGND VGND VPWR VPWR _20333_/X sky130_fd_sc_hd__a211o_4
XANTENNA__11768__A _15484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23052_ _17636_/X _23038_/B VGND VGND VPWR VPWR _23053_/C sky130_fd_sc_hd__or2_4
XFILLER_66_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20264_ _20242_/X VGND VGND VPWR VPWR _20517_/A sky130_fd_sc_hd__inv_2
XANTENNA__22361__A _22354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22003_ _21840_/X _22002_/X _23497_/Q _21999_/X VGND VGND VPWR VPWR _22003_/X sky130_fd_sc_hd__o22a_4
XFILLER_1_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20195_ _16929_/X _17025_/A _17072_/A _20195_/D VGND VGND VPWR VPWR _20195_/X sky130_fd_sc_hd__and4_4
XFILLER_9_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12599__A _12599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_106_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR _23314_/CLK sky130_fd_sc_hd__clkbuf_1
X_23954_ _23986_/CLK _23954_/D VGND VGND VPWR VPWR _23954_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20737__A1 _20622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21934__B1 _12263_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22905_ _22886_/X _18607_/X _22887_/X _22904_/X VGND VGND VPWR VPWR _22906_/A sky130_fd_sc_hd__a211o_4
XANTENNA__21705__A _21705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23885_ _23698_/CLK _23885_/D VGND VGND VPWR VPWR _23885_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22836_ _17504_/Y _22825_/X _22831_/X _22835_/X VGND VGND VPWR VPWR _22837_/A sky130_fd_sc_hd__a211o_4
XANTENNA__15703__A _12742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22767_ _22744_/Y _22765_/B VGND VGND VPWR VPWR _22767_/Y sky130_fd_sc_hd__nand2_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _13029_/A VGND VGND VPWR VPWR _12520_/X sky130_fd_sc_hd__buf_2
XANTENNA__13223__A _12383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21718_ _21553_/X _21712_/X _23658_/Q _21716_/X VGND VGND VPWR VPWR _21718_/X sky130_fd_sc_hd__o22a_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22698_ _21265_/A _22693_/X _15573_/B _22697_/X VGND VGND VPWR VPWR _23083_/D sky130_fd_sc_hd__o22a_4
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22536__A _22536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12451_ _12494_/A VGND VGND VPWR VPWR _12887_/A sky130_fd_sc_hd__buf_2
X_21649_ _21519_/X _21648_/X _23704_/Q _21645_/X VGND VGND VPWR VPWR _23704_/D sky130_fd_sc_hd__o22a_4
X_24437_ _24277_/CLK _18780_/X HRESETn VGND VGND VPWR VPWR _20470_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_51_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16534__A _11936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15170_ _14152_/A _15241_/B VGND VGND VPWR VPWR _15170_/X sky130_fd_sc_hd__or2_4
X_12382_ _12398_/A _12382_/B _12382_/C VGND VGND VPWR VPWR _12389_/B sky130_fd_sc_hd__and3_4
X_24368_ _23358_/CLK _24368_/D HRESETn VGND VGND VPWR VPWR _24368_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21465__A2 _21463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20122__C1 _18940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24173__D _19792_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22662__B2 _22626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12781__B _24020_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14121_ _14121_/A _23913_/Q VGND VGND VPWR VPWR _14123_/B sky130_fd_sc_hd__or2_4
XANTENNA__16253__B _16253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23319_ _23316_/CLK _23319_/D VGND VGND VPWR VPWR _22307_/A sky130_fd_sc_hd__dfxtp_4
X_24299_ _24299_/CLK _24299_/D HRESETn VGND VGND VPWR VPWR _19120_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_84_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14052_ _14035_/A _13970_/B VGND VGND VPWR VPWR _14052_/X sky130_fd_sc_hd__or2_4
XANTENNA__22414__A1 _22413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22414__B2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14989__A _14121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13003_ _12887_/A _13003_/B _13002_/X VGND VGND VPWR VPWR _13004_/C sky130_fd_sc_hd__and3_4
X_18860_ _15379_/X _18855_/X _24386_/Q _18856_/X VGND VGND VPWR VPWR _24386_/D sky130_fd_sc_hd__o22a_4
X_17811_ _17811_/A VGND VGND VPWR VPWR _17812_/A sky130_fd_sc_hd__buf_2
XFILLER_67_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18791_ _15780_/B _18788_/X _24430_/Q _18789_/X VGND VGND VPWR VPWR _18791_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17742_ _17734_/A _17111_/X _17734_/X _17741_/X VGND VGND VPWR VPWR _17742_/X sky130_fd_sc_hd__o22a_4
X_14954_ _11661_/A _14954_/B _14953_/X VGND VGND VPWR VPWR _14986_/B sky130_fd_sc_hd__or3_4
XFILLER_3_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12302__A _12302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13905_ _13909_/A _13831_/B VGND VGND VPWR VPWR _13907_/B sky130_fd_sc_hd__or2_4
XFILLER_1_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17673_ _17673_/A VGND VGND VPWR VPWR _17674_/A sky130_fd_sc_hd__buf_2
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14885_ _12301_/A _14885_/B _14884_/X VGND VGND VPWR VPWR _14885_/X sky130_fd_sc_hd__or3_4
XANTENNA__16709__A _11875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19412_ _19411_/X _18710_/X _19411_/X _24192_/Q VGND VGND VPWR VPWR _24192_/D sky130_fd_sc_hd__a2bb2o_4
X_16624_ _11772_/X VGND VGND VPWR VPWR _16624_/X sky130_fd_sc_hd__buf_2
XANTENNA__15613__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13836_ _12269_/A _13813_/X _13820_/X _13827_/X _13835_/X VGND VGND VPWR VPWR _13836_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19346__B2 _24231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19343_ _19336_/A VGND VGND VPWR VPWR _19343_/X sky130_fd_sc_hd__buf_2
X_16555_ _12022_/A _23932_/Q VGND VGND VPWR VPWR _16557_/B sky130_fd_sc_hd__or2_4
XFILLER_56_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15332__B _15273_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13767_ _12652_/A _13767_/B VGND VGND VPWR VPWR _13768_/C sky130_fd_sc_hd__or2_4
XANTENNA__21153__B2 _21151_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15506_ _13097_/A _15504_/X _15506_/C VGND VGND VPWR VPWR _15507_/C sky130_fd_sc_hd__and3_4
XANTENNA__13133__A _13133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12718_ _12284_/X _23892_/Q VGND VGND VPWR VPWR _12720_/B sky130_fd_sc_hd__or2_4
X_19274_ _19216_/A _19216_/B _19273_/Y VGND VGND VPWR VPWR _19274_/X sky130_fd_sc_hd__o21a_4
X_16486_ _16473_/X _16417_/B VGND VGND VPWR VPWR _16487_/C sky130_fd_sc_hd__or2_4
X_13698_ _13697_/X _13698_/B VGND VGND VPWR VPWR _13699_/C sky130_fd_sc_hd__or2_4
XANTENNA__22446__A _22446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18225_ _17668_/Y _18165_/X _17667_/X VGND VGND VPWR VPWR _18225_/X sky130_fd_sc_hd__o21a_4
X_15437_ _13636_/A _15437_/B VGND VGND VPWR VPWR _15437_/X sky130_fd_sc_hd__or2_4
X_12649_ _12951_/A _12647_/X _12648_/X VGND VGND VPWR VPWR _12649_/X sky130_fd_sc_hd__and3_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12972__A _13118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16444__A _16443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22102__B1 _23443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18156_ _17456_/Y _18155_/X _17525_/X VGND VGND VPWR VPWR _18156_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15368_ _14009_/A _15368_/B _15368_/C VGND VGND VPWR VPWR _15369_/C sky130_fd_sc_hd__and3_4
XANTENNA__22653__B2 _22647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12691__B _12774_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17107_ _14786_/Y _17010_/X _17018_/X _17106_/X VGND VGND VPWR VPWR _17201_/A sky130_fd_sc_hd__o22a_4
X_14319_ _15574_/A VGND VGND VPWR VPWR _14432_/A sky130_fd_sc_hd__buf_2
X_18087_ _18062_/X _18068_/Y _18080_/X _18085_/X _18086_/Y VGND VGND VPWR VPWR _18087_/X
+ sky130_fd_sc_hd__a32o_4
X_15299_ _14758_/A _15299_/B VGND VGND VPWR VPWR _15299_/X sky130_fd_sc_hd__or2_4
X_17038_ _17037_/Y VGND VGND VPWR VPWR _17039_/A sky130_fd_sc_hd__buf_2
XANTENNA__21208__A2 _21204_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18989_ _18971_/X _18986_/X _18988_/X _18982_/A VGND VGND VPWR VPWR _24341_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15843__B1 _15834_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22708__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13308__A _15685_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12212__A _12211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20719__A1 _24235_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20951_ _20825_/X _20950_/X VGND VGND VPWR VPWR _20951_/Y sky130_fd_sc_hd__nor2_4
XFILLER_113_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21392__B2 _21387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15523__A _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23670_ _23920_/CLK _23670_/D VGND VGND VPWR VPWR _12246_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20882_ _20681_/X _20881_/X _19083_/A _18870_/X VGND VGND VPWR VPWR _20882_/X sky130_fd_sc_hd__o22a_4
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22621_ _22621_/A VGND VGND VPWR VPWR _22636_/A sky130_fd_sc_hd__buf_2
XFILLER_81_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22341__B1 _12132_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18834__A _18834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13043__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22552_ _22442_/X _22550_/X _13712_/B _22547_/X VGND VGND VPWR VPWR _23176_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21503_ _21515_/A VGND VGND VPWR VPWR _21503_/X sky130_fd_sc_hd__buf_2
XFILLER_10_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13978__A _12196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22483_ _22483_/A VGND VGND VPWR VPWR _22483_/X sky130_fd_sc_hd__buf_2
XANTENNA__12882__A _13960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16354__A _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24222_ _24216_/CLK _19365_/X HRESETn VGND VGND VPWR VPWR _24222_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12188__A2 _12184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21434_ _21270_/X _21433_/X _23817_/Q _21430_/X VGND VGND VPWR VPWR _23817_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22644__B2 _22640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24153_ _24162_/CLK _24153_/D HRESETn VGND VGND VPWR VPWR _24153_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21365_ _21239_/X _21362_/X _12332_/B _21359_/X VGND VGND VPWR VPWR _21365_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19665__A _19800_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23104_ _23104_/CLK _22662_/X VGND VGND VPWR VPWR _14962_/B sky130_fd_sc_hd__dfxtp_4
X_20316_ _20280_/X _20315_/X _24093_/Q _20203_/X VGND VGND VPWR VPWR _20316_/X sky130_fd_sc_hd__o22a_4
X_24084_ _24084_/CLK _24084_/D VGND VGND VPWR VPWR _24084_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21296_ _21296_/A VGND VGND VPWR VPWR _21784_/B sky130_fd_sc_hd__buf_2
XANTENNA__22091__A _20441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20898__A1_N _19734_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23035_ _23014_/X _17646_/A _23026_/X _23034_/X VGND VGND VPWR VPWR _23036_/A sky130_fd_sc_hd__a211o_4
XFILLER_46_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20247_ _20453_/A VGND VGND VPWR VPWR _20247_/X sky130_fd_sc_hd__buf_2
XFILLER_81_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14602__A _15030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21080__B1 _24021_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20178_ _19313_/A _20177_/X VGND VGND VPWR VPWR _20178_/X sky130_fd_sc_hd__or2_4
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13218__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12122__A _16071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18728__B _18728_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11951_ _11890_/A VGND VGND VPWR VPWR _14880_/A sky130_fd_sc_hd__buf_2
X_23937_ _23145_/CLK _23937_/D VGND VGND VPWR VPWR _15156_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_79_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20186__A2 _17737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16529__A _16541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22580__B1 _15967_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24351__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15433__A _12211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11882_ _15706_/A VGND VGND VPWR VPWR _15784_/A sky130_fd_sc_hd__buf_2
X_14670_ _14071_/A _14656_/X _14669_/X VGND VGND VPWR VPWR _14670_/X sky130_fd_sc_hd__and3_4
X_23868_ _23867_/CLK _23868_/D VGND VGND VPWR VPWR _23868_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16248__B _16248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13621_ _15424_/A _13618_/X _13621_/C VGND VGND VPWR VPWR _13621_/X sky130_fd_sc_hd__and3_4
X_22819_ _15910_/Y _22814_/X _22795_/X _22818_/X VGND VGND VPWR VPWR _22820_/B sky130_fd_sc_hd__o22a_4
XANTENNA__14049__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23799_ _23632_/CLK _23799_/D VGND VGND VPWR VPWR _16217_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21135__B2 _21130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16340_ _16185_/A _16272_/B VGND VGND VPWR VPWR _16340_/X sky130_fd_sc_hd__or2_4
XANTENNA__24244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13552_ _13551_/X _13552_/B VGND VGND VPWR VPWR _13555_/B sky130_fd_sc_hd__or2_4
XFILLER_105_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12503_ _12503_/A _12503_/B _12502_/X VGND VGND VPWR VPWR _12503_/X sky130_fd_sc_hd__or3_4
XANTENNA__13888__A _13895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13483_ _13483_/A _13483_/B _13483_/C VGND VGND VPWR VPWR _13483_/X sky130_fd_sc_hd__or3_4
X_16271_ _11852_/X _16247_/X _16255_/X _16262_/X _16270_/X VGND VGND VPWR VPWR _16271_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_41_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12792__A _12792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18010_ _17889_/A VGND VGND VPWR VPWR _18174_/C sky130_fd_sc_hd__buf_2
X_12434_ _12434_/A _12433_/Y VGND VGND VPWR VPWR _12434_/X sky130_fd_sc_hd__or2_4
X_15222_ _15234_/A _15159_/B VGND VGND VPWR VPWR _15222_/X sky130_fd_sc_hd__or2_4
XANTENNA__22635__A1 _22413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21438__A2 _21433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17079__B _17224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22635__B2 _22633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12365_ _15484_/A VGND VGND VPWR VPWR _13557_/A sky130_fd_sc_hd__buf_2
X_15153_ _14128_/A _15153_/B VGND VGND VPWR VPWR _15153_/X sky130_fd_sc_hd__and2_4
XFILLER_86_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14104_ _14315_/A _23657_/Q VGND VGND VPWR VPWR _14108_/B sky130_fd_sc_hd__or2_4
XFILLER_5_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15084_ _15108_/A _15080_/X _15084_/C VGND VGND VPWR VPWR _15084_/X sky130_fd_sc_hd__or3_4
X_19961_ _19985_/A VGND VGND VPWR VPWR _19961_/X sky130_fd_sc_hd__buf_2
X_12296_ _12742_/A VGND VGND VPWR VPWR _15685_/A sky130_fd_sc_hd__buf_2
X_14035_ _14035_/A _23530_/Q VGND VGND VPWR VPWR _14036_/C sky130_fd_sc_hd__or2_4
X_18912_ _18898_/A VGND VGND VPWR VPWR _18912_/X sky130_fd_sc_hd__buf_2
XFILLER_45_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19892_ _20849_/B VGND VGND VPWR VPWR _20875_/A sky130_fd_sc_hd__buf_2
XFILLER_80_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20949__A1 _20494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20949__B2 _20453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18843_ _13575_/X _18841_/X _20595_/A _18842_/X VGND VGND VPWR VPWR _24399_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21610__A2 _21605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15327__B _15262_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18774_ _18781_/A VGND VGND VPWR VPWR _18774_/X sky130_fd_sc_hd__buf_2
XANTENNA__12032__A _11837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15986_ _15986_/A _15986_/B _15986_/C VGND VGND VPWR VPWR _15987_/C sky130_fd_sc_hd__and3_4
X_17725_ _17724_/X _17290_/X _17720_/X VGND VGND VPWR VPWR _17745_/B sky130_fd_sc_hd__a21bo_4
XFILLER_76_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14937_ _14937_/A _23552_/Q VGND VGND VPWR VPWR _14938_/C sky130_fd_sc_hd__or2_4
XFILLER_97_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16439__A _13447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12967__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21374__B2 _21373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11871__A _13014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15343__A _12567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17656_ _17659_/A _17654_/Y _17658_/A VGND VGND VPWR VPWR _18003_/A sky130_fd_sc_hd__o21ai_4
X_14868_ _14867_/X _14868_/B VGND VGND VPWR VPWR _14868_/X sky130_fd_sc_hd__or2_4
XFILLER_63_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16158__B _16158_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19319__B2 _24250_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16607_ _11821_/A VGND VGND VPWR VPWR _16617_/A sky130_fd_sc_hd__buf_2
X_13819_ _13796_/A _13819_/B _13819_/C VGND VGND VPWR VPWR _13820_/C sky130_fd_sc_hd__and3_4
XFILLER_63_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17587_ _17481_/X _17489_/X _17493_/Y VGND VGND VPWR VPWR _17587_/X sky130_fd_sc_hd__a21o_4
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14799_ _14050_/A _14799_/B _14798_/X VGND VGND VPWR VPWR _14799_/X sky130_fd_sc_hd__and3_4
X_19326_ _19325_/X _18195_/X _19325_/X _24245_/Q VGND VGND VPWR VPWR _24245_/D sky130_fd_sc_hd__a2bb2o_4
X_16538_ _16538_/A _24028_/Q VGND VGND VPWR VPWR _16541_/B sky130_fd_sc_hd__or2_4
XANTENNA__21677__A2 _21676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22874__A1 _16596_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22176__A _22169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19257_ _19257_/A VGND VGND VPWR VPWR _19257_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13798__A _15413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16469_ _16194_/A _16467_/X _16468_/X VGND VGND VPWR VPWR _16470_/C sky130_fd_sc_hd__and3_4
X_18208_ _18267_/A _18205_/X _18208_/C _18207_/X VGND VGND VPWR VPWR _18209_/A sky130_fd_sc_hd__or4_4
XANTENNA__21429__A2 _21426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19188_ _24294_/Q _19115_/B _19187_/Y VGND VGND VPWR VPWR _24294_/D sky130_fd_sc_hd__o21a_4
XANTENNA__22904__A _22899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18139_ _18267_/A _18135_/X _18136_/Y _18139_/D VGND VGND VPWR VPWR _18140_/A sky130_fd_sc_hd__or4_4
XFILLER_117_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21150_ _20819_/X _21147_/X _13792_/B _21144_/X VGND VGND VPWR VPWR _23975_/D sky130_fd_sc_hd__o22a_4
XFILLER_117_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20101_ _20098_/X _20100_/Y _20089_/C VGND VGND VPWR VPWR _20101_/Y sky130_fd_sc_hd__o21ai_4
X_21081_ _20509_/X _21075_/X _24020_/Q _21079_/X VGND VGND VPWR VPWR _21081_/X sky130_fd_sc_hd__o22a_4
XFILLER_99_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15518__A _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14422__A _14040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20032_ _20031_/X VGND VGND VPWR VPWR _20032_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21601__A2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15237__B _15180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13038__A _13015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21983_ _21807_/X _21981_/X _23511_/Q _21978_/X VGND VGND VPWR VPWR _23511_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21365__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15253__A _11954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11781__A _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20934_ _20282_/A _20933_/X VGND VGND VPWR VPWR _20934_/Y sky130_fd_sc_hd__nand2_4
X_23722_ _24011_/CLK _23722_/D VGND VGND VPWR VPWR _23722_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18230__A1 _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _20616_/X _20853_/X _20757_/X _20864_/Y VGND VGND VPWR VPWR _20865_/X sky130_fd_sc_hd__a211o_4
X_23653_ _23973_/CLK _21725_/X VGND VGND VPWR VPWR _14523_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21117__B2 _21116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18564__A _18082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22604_ _22583_/A VGND VGND VPWR VPWR _22604_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23584_ _23584_/CLK _23584_/D VGND VGND VPWR VPWR _23584_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22865__A1 _17542_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21668__A2 _21662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20796_ _22127_/A VGND VGND VPWR VPWR _21843_/A sky130_fd_sc_hd__buf_2
XANTENNA__22086__A _20393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22535_ _22413_/X _22529_/X _12773_/B _22533_/X VGND VGND VPWR VPWR _23188_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20876__B1 HRDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15700__B _15700_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13501__A _12965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22466_ _22465_/X VGND VGND VPWR VPWR _22471_/A sky130_fd_sc_hd__buf_2
XFILLER_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21417_ _21241_/X _21412_/X _12648_/B _21416_/X VGND VGND VPWR VPWR _21417_/X sky130_fd_sc_hd__o22a_4
X_24205_ _24208_/CLK _19394_/X HRESETn VGND VGND VPWR VPWR _24205_/Q sky130_fd_sc_hd__dfrtp_4
X_22397_ _22396_/X _22392_/X _16744_/B _22387_/X VGND VGND VPWR VPWR _22397_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12117__A _16071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16812__A _16077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12150_ _11772_/X _12142_/X _12149_/X VGND VGND VPWR VPWR _12150_/X sky130_fd_sc_hd__and3_4
X_24136_ _24239_/CLK _19980_/Y HRESETn VGND VGND VPWR VPWR _17644_/A sky130_fd_sc_hd__dfrtp_4
X_21348_ _21348_/A _21348_/B _21348_/C _20199_/B VGND VGND VPWR VPWR _21348_/X sky130_fd_sc_hd__or4_4
XFILLER_68_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11956__A _15533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12081_ _11992_/X _12081_/B VGND VGND VPWR VPWR _12081_/X sky130_fd_sc_hd__and2_4
X_24067_ _23270_/CLK _24067_/D VGND VGND VPWR VPWR _14770_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15428__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21279_ _21277_/X _21271_/X _14292_/B _21278_/X VGND VGND VPWR VPWR _23910_/D sky130_fd_sc_hd__o22a_4
XFILLER_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23018_ _23018_/A _23018_/B _23018_/C VGND VGND VPWR VPWR _23018_/X sky130_fd_sc_hd__and3_4
XFILLER_104_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15147__B _23553_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15840_ _12920_/A _15838_/X _15839_/X VGND VGND VPWR VPWR _15841_/C sky130_fd_sc_hd__and3_4
XFILLER_49_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17643__A _17766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21165__A _21180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15771_ _12765_/X _15771_/B _15770_/X VGND VGND VPWR VPWR _15771_/X sky130_fd_sc_hd__and3_4
X_12983_ _12660_/A _12983_/B VGND VGND VPWR VPWR _12983_/X sky130_fd_sc_hd__or2_4
XANTENNA__12787__A _12787_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21356__A1 _21221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20159__A2 IRQ[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21356__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17510_ _13278_/X _17510_/B VGND VGND VPWR VPWR _17510_/X sky130_fd_sc_hd__and2_4
X_14722_ _15387_/A VGND VGND VPWR VPWR _14722_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24082__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11934_ _11933_/X VGND VGND VPWR VPWR _16121_/A sky130_fd_sc_hd__buf_2
X_18490_ _18399_/Y _17422_/A _17424_/X VGND VGND VPWR VPWR _18538_/A sky130_fd_sc_hd__o21a_4
XFILLER_40_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22156__A2_N _22155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17441_ _17037_/Y _17440_/X _17042_/A VGND VGND VPWR VPWR _17442_/A sky130_fd_sc_hd__o21a_4
X_14653_ _15190_/A VGND VGND VPWR VPWR _14672_/A sky130_fd_sc_hd__buf_2
X_11865_ _11606_/A VGND VGND VPWR VPWR _13955_/A sky130_fd_sc_hd__buf_2
XFILLER_96_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21108__B2 _21072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13604_ _11611_/A VGND VGND VPWR VPWR _13959_/A sky130_fd_sc_hd__buf_2
X_17372_ _17370_/X _17371_/X VGND VGND VPWR VPWR _17372_/X sky130_fd_sc_hd__or2_4
X_11796_ _11661_/A VGND VGND VPWR VPWR _11797_/A sky130_fd_sc_hd__inv_2
X_14584_ _14149_/A _24004_/Q VGND VGND VPWR VPWR _14584_/X sky130_fd_sc_hd__or2_4
X_19111_ _19111_/A _19197_/A VGND VGND VPWR VPWR _19112_/B sky130_fd_sc_hd__and2_4
X_16323_ _16323_/A _23577_/Q VGND VGND VPWR VPWR _16324_/C sky130_fd_sc_hd__or2_4
X_13535_ _13563_/A _13535_/B _13534_/X VGND VGND VPWR VPWR _13536_/C sky130_fd_sc_hd__and3_4
XFILLER_18_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20331__A2 _20329_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13349__A1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19042_ _11516_/B VGND VGND VPWR VPWR _19042_/Y sky130_fd_sc_hd__inv_2
X_16254_ _16147_/A _16251_/X _16253_/X VGND VGND VPWR VPWR _16254_/X sky130_fd_sc_hd__and3_4
X_13466_ _13450_/A _13466_/B VGND VGND VPWR VPWR _13467_/C sky130_fd_sc_hd__or2_4
XFILLER_16_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22608__B2 _22604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14226__B _23945_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15205_ _14252_/A _15150_/B VGND VGND VPWR VPWR _15206_/C sky130_fd_sc_hd__or2_4
X_12417_ _15889_/A _12411_/X _12416_/X VGND VGND VPWR VPWR _12417_/X sky130_fd_sc_hd__or3_4
X_16185_ _16185_/A VGND VGND VPWR VPWR _16219_/A sky130_fd_sc_hd__buf_2
X_13397_ _12829_/A VGND VGND VPWR VPWR _13397_/X sky130_fd_sc_hd__buf_2
XANTENNA__12027__A _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_14_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR _23107_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21292__B1 _14879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15136_ _11954_/A _15197_/B VGND VGND VPWR VPWR _15136_/X sky130_fd_sc_hd__or2_4
X_12348_ _15774_/A _12344_/X _12348_/C VGND VGND VPWR VPWR _12354_/B sky130_fd_sc_hd__and3_4
XFILLER_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_77_0_HCLK clkbuf_6_38_0_HCLK/X VGND VGND VPWR VPWR _23260_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12279_ _13026_/A _12278_/X VGND VGND VPWR VPWR _12279_/X sky130_fd_sc_hd__and2_4
X_15067_ _15115_/A _15062_/X _15066_/X VGND VGND VPWR VPWR _15068_/C sky130_fd_sc_hd__or3_4
X_19944_ _17779_/X _19944_/B _19944_/C _19944_/D VGND VGND VPWR VPWR _19945_/A sky130_fd_sc_hd__or4_4
XFILLER_9_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21059__B _22017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19788__A1 _19866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14018_ _14847_/A _14013_/X _14018_/C VGND VGND VPWR VPWR _14019_/C sky130_fd_sc_hd__or3_4
XFILLER_29_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15057__B _23711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19875_ _19585_/X _19874_/X _16929_/B _19549_/X VGND VGND VPWR VPWR _19875_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19752__B HRDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18826_ _16514_/X _18818_/X _24410_/Q _18821_/X VGND VGND VPWR VPWR _24410_/D sky130_fd_sc_hd__o22a_4
XFILLER_116_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21075__A _21075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18757_ _16916_/A VGND VGND VPWR VPWR _18757_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15969_ _15997_/A _15969_/B VGND VGND VPWR VPWR _15970_/C sky130_fd_sc_hd__or2_4
XFILLER_23_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12697__A _12198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22544__B1 _15659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17708_ _17708_/A _17413_/X VGND VGND VPWR VPWR _17708_/X sky130_fd_sc_hd__or2_4
XFILLER_97_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18688_ _16925_/Y _18683_/X _16925_/Y _18687_/X VGND VGND VPWR VPWR _18688_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17639_ _17639_/A VGND VGND VPWR VPWR _17639_/X sky130_fd_sc_hd__buf_2
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20570__A2 _20421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20650_ _20650_/A _20822_/B VGND VGND VPWR VPWR _20650_/X sky130_fd_sc_hd__or2_4
XFILLER_36_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22847__A1 _14493_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15801__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14785__B1 _11594_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19309_ _19305_/Y _19308_/A _19304_/X _19308_/Y VGND VGND VPWR VPWR _19309_/X sky130_fd_sc_hd__o22a_4
XFILLER_17_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20581_ _20403_/X _20580_/X _24272_/Q _20497_/X VGND VGND VPWR VPWR _20581_/X sky130_fd_sc_hd__o22a_4
X_22320_ _22320_/A VGND VGND VPWR VPWR _23306_/D sky130_fd_sc_hd__buf_2
XANTENNA__21303__A2_N _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22251_ _22068_/A _21634_/B _22383_/C _21634_/D VGND VGND VPWR VPWR _22251_/X sky130_fd_sc_hd__or4_4
XANTENNA__19476__B1 HRDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21202_ _20838_/X _21197_/X _14302_/B _21201_/X VGND VGND VPWR VPWR _21202_/X sky130_fd_sc_hd__o22a_4
X_22182_ _22117_/X _22179_/X _23404_/Q _22176_/X VGND VGND VPWR VPWR _22182_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21822__A2 _21817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16351__B _16283_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21133_ _21133_/A VGND VGND VPWR VPWR _21133_/X sky130_fd_sc_hd__buf_2
XFILLER_105_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15248__A _11798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19943__A _18066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14152__A _14152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19779__B2 _19789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21064_ _21079_/A VGND VGND VPWR VPWR _21072_/A sky130_fd_sc_hd__buf_2
XFILLER_8_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20015_ _18289_/X _20009_/X _20014_/Y _19996_/X VGND VGND VPWR VPWR _20015_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13991__A _13991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17463__A _17156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_28_0_HCLK_A clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21338__A1 _21277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16079__A _16008_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21338__B2 _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12400__A _12826_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21889__A2 _21887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21966_ _23518_/Q VGND VGND VPWR VPWR _21966_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18754__A2 _17126_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23705_ _23770_/CLK _21647_/X VGND VGND VPWR VPWR _16296_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _20872_/X _20916_/X _14770_/B _20839_/X VGND VGND VPWR VPWR _24067_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13215__B _24017_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _21833_/X _21894_/X _15471_/B _21891_/X VGND VGND VPWR VPWR _23564_/D sky130_fd_sc_hd__o22a_4
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16807__A _16800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _14175_/A VGND VGND VPWR VPWR _13991_/A sky130_fd_sc_hd__buf_2
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _20842_/X _20844_/X _20845_/X HRDATA[14] _20847_/X VGND VGND VPWR VPWR _20848_/X
+ sky130_fd_sc_hd__a32o_4
X_23636_ _23316_/CLK _21754_/X VGND VGND VPWR VPWR _12836_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22838__A1 _17109_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _11580_/Y VGND VGND VPWR VPWR _11634_/A sky130_fd_sc_hd__buf_2
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ _21555_/A VGND VGND VPWR VPWR _20779_/X sky130_fd_sc_hd__buf_2
X_23567_ _23827_/CLK _21893_/X VGND VGND VPWR VPWR _13521_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _13303_/X _13318_/X _13319_/X VGND VGND VPWR VPWR _13320_/X sky130_fd_sc_hd__and3_4
XANTENNA__16880__A2_N _16816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22518_ _22533_/A VGND VGND VPWR VPWR _22518_/X sky130_fd_sc_hd__buf_2
XFILLER_11_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23498_ _23819_/CLK _23498_/D VGND VGND VPWR VPWR _23498_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13251_ _13211_/A _13251_/B _13251_/C VGND VGND VPWR VPWR _13252_/C sky130_fd_sc_hd__or3_4
X_22449_ _22134_/A VGND VGND VPWR VPWR _22449_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12202_ _12202_/A VGND VGND VPWR VPWR _12203_/A sky130_fd_sc_hd__buf_2
X_13182_ _15697_/A _13249_/B VGND VGND VPWR VPWR _13182_/X sky130_fd_sc_hd__or2_4
XANTENNA__24181__D _24181_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21813__A2 _21805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12133_ _12169_/A _12131_/X _12133_/C VGND VGND VPWR VPWR _12134_/C sky130_fd_sc_hd__and3_4
XANTENNA__11686__A _12421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24119_ _24202_/CLK _20061_/Y HRESETn VGND VGND VPWR VPWR _16957_/A sky130_fd_sc_hd__dfrtp_4
X_17990_ _18081_/B _17583_/X _17581_/Y VGND VGND VPWR VPWR _17990_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23322__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24448__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18690__B2 _11629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21026__B1 _24054_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12064_ _12093_/A _23677_/Q VGND VGND VPWR VPWR _12064_/X sky130_fd_sc_hd__or2_4
X_16941_ _24135_/Q VGND VGND VPWR VPWR _17646_/A sky130_fd_sc_hd__inv_2
XFILLER_61_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14997__A _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21577__B2 _21515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19660_ _19719_/A _19718_/B VGND VGND VPWR VPWR _19661_/B sky130_fd_sc_hd__or2_4
XFILLER_78_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16872_ _16853_/X _16855_/X _16870_/X _16872_/D VGND VGND VPWR VPWR _16872_/X sky130_fd_sc_hd__and4_4
XFILLER_93_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18611_ _18607_/X _18610_/X _17726_/X VGND VGND VPWR VPWR _18611_/X sky130_fd_sc_hd__or3_4
X_15823_ _15823_/A _15821_/X _15823_/C VGND VGND VPWR VPWR _15823_/X sky130_fd_sc_hd__and3_4
XFILLER_77_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19591_ _19729_/B VGND VGND VPWR VPWR _19592_/A sky130_fd_sc_hd__buf_2
XANTENNA__15605__B _23659_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21329__B2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18542_ _18392_/A _18185_/Y VGND VGND VPWR VPWR _18542_/X sky130_fd_sc_hd__and2_4
X_15754_ _15724_/A _15689_/B VGND VGND VPWR VPWR _15754_/X sky130_fd_sc_hd__or2_4
X_12966_ _12959_/A _23827_/Q VGND VGND VPWR VPWR _12967_/C sky130_fd_sc_hd__or2_4
XANTENNA__12310__A _15552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22719__A _22967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14705_ _14664_/X _14703_/X _14704_/X VGND VGND VPWR VPWR _14705_/X sky130_fd_sc_hd__and3_4
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21623__A _21602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11917_ _11916_/X VGND VGND VPWR VPWR _11995_/A sky130_fd_sc_hd__buf_2
X_18473_ _17382_/A _18473_/B VGND VGND VPWR VPWR _18473_/X sky130_fd_sc_hd__or2_4
X_15685_ _15685_/A _15685_/B VGND VGND VPWR VPWR _15687_/B sky130_fd_sc_hd__or2_4
X_12897_ _12868_/A _23603_/Q VGND VGND VPWR VPWR _12899_/B sky130_fd_sc_hd__or2_4
X_17424_ _13920_/X _17424_/B VGND VGND VPWR VPWR _17424_/X sky130_fd_sc_hd__or2_4
X_14636_ _13611_/A _14634_/X _14636_/C VGND VGND VPWR VPWR _14637_/C sky130_fd_sc_hd__and3_4
XANTENNA__22829__A1 _17477_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11848_ _13682_/A VGND VGND VPWR VPWR _13056_/A sky130_fd_sc_hd__buf_2
XFILLER_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12964__B _12964_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17355_ _15453_/Y _17340_/X _17020_/A _17354_/X VGND VGND VPWR VPWR _17356_/B sky130_fd_sc_hd__o22a_4
X_14567_ _14493_/Y _14564_/X _14566_/X VGND VGND VPWR VPWR _14567_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21061__C _21162_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11779_ _11821_/A _11779_/B VGND VGND VPWR VPWR _11779_/X sky130_fd_sc_hd__or2_4
X_16306_ _16303_/X _16306_/B _16306_/C VGND VGND VPWR VPWR _16306_/X sky130_fd_sc_hd__and3_4
XFILLER_14_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13141__A _12240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13518_ _13572_/A _13506_/X _13518_/C VGND VGND VPWR VPWR _13538_/B sky130_fd_sc_hd__and3_4
X_17286_ _17286_/A VGND VGND VPWR VPWR _17413_/B sky130_fd_sc_hd__buf_2
X_14498_ _14494_/X _14495_/X _14497_/X VGND VGND VPWR VPWR _14498_/X sky130_fd_sc_hd__and3_4
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22454__A _20915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19025_ _11519_/A _11519_/B _19019_/Y VGND VGND VPWR VPWR _19025_/Y sky130_fd_sc_hd__a21oi_4
X_16237_ _16236_/X VGND VGND VPWR VPWR _16237_/Y sky130_fd_sc_hd__inv_2
X_13449_ _13448_/X _23311_/Q VGND VGND VPWR VPWR _13451_/B sky130_fd_sc_hd__or2_4
XANTENNA__22057__A2 _22052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12980__A _12980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20068__A1 _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16168_ _16198_/A _16161_/X _16168_/C VGND VGND VPWR VPWR _16168_/X sky130_fd_sc_hd__or3_4
XFILLER_66_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11596__A _11596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15119_ _15118_/X VGND VGND VPWR VPWR _15119_/X sky130_fd_sc_hd__buf_2
XANTENNA__15068__A _14071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16099_ _16127_/A _16175_/B VGND VGND VPWR VPWR _16104_/B sky130_fd_sc_hd__or2_4
XFILLER_102_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19927_ _19927_/A _11591_/C _18812_/C _19926_/X VGND VGND VPWR VPWR _19927_/X sky130_fd_sc_hd__or4_4
XFILLER_29_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17283__A _14336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_7_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR _24241_/CLK sky130_fd_sc_hd__clkbuf_1
X_19858_ _19667_/A _19856_/X _19445_/A _19857_/X VGND VGND VPWR VPWR _19858_/X sky130_fd_sc_hd__a211o_4
XANTENNA__18433__B2 _18432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14700__A _14673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18809_ _15121_/X _18781_/A _20966_/A _18782_/A VGND VGND VPWR VPWR _24416_/D sky130_fd_sc_hd__o22a_4
XFILLER_84_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19789_ _19622_/A _19789_/B VGND VGND VPWR VPWR _19789_/X sky130_fd_sc_hd__and2_4
XFILLER_37_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21820_ _21819_/X _21817_/X _23602_/Q _21812_/X VGND VGND VPWR VPWR _21820_/X sky130_fd_sc_hd__o22a_4
XFILLER_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12220__A _13054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22629__A _22636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21751_ _21524_/X _21748_/X _12424_/B _21745_/X VGND VGND VPWR VPWR _23638_/D sky130_fd_sc_hd__o22a_4
XFILLER_58_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16627__A _16616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20702_ _20802_/A _20701_/X VGND VGND VPWR VPWR _20702_/X sky130_fd_sc_hd__or2_4
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15531__A _12307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21682_ _21578_/X _21662_/A _23679_/Q _21637_/X VGND VGND VPWR VPWR _23679_/D sky130_fd_sc_hd__o22a_4
X_24470_ _23522_/CLK _24470_/D HRESETn VGND VGND VPWR VPWR _19995_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20633_ _20444_/X _20621_/Y _20631_/X _20632_/Y _20459_/X VGND VGND VPWR VPWR _20634_/B
+ sky130_fd_sc_hd__a32o_4
X_23421_ _23100_/CLK _23421_/D VGND VGND VPWR VPWR _23421_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22296__A2 _22293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13051__A _12465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23352_ _23383_/CLK _23352_/D VGND VGND VPWR VPWR _23352_/Q sky130_fd_sc_hd__dfxtp_4
X_20564_ _20518_/X _20563_/X _24337_/Q _20525_/X VGND VGND VPWR VPWR _20564_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22303_ _16775_/B VGND VGND VPWR VPWR _23323_/D sky130_fd_sc_hd__buf_2
XFILLER_109_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23283_ _23859_/CLK _22355_/X VGND VGND VPWR VPWR _23283_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22048__A2 _22045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20495_ _24404_/Q _20405_/X _24436_/Q _20449_/X VGND VGND VPWR VPWR _20495_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12890__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22234_ _22119_/X _22229_/X _23371_/Q _22233_/X VGND VGND VPWR VPWR _23371_/D sky130_fd_sc_hd__o22a_4
XFILLER_30_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18121__B1 _17259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22165_ _22172_/A VGND VGND VPWR VPWR _22165_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_60_0_HCLK clkbuf_6_30_0_HCLK/X VGND VGND VPWR VPWR _23342_/CLK sky130_fd_sc_hd__clkbuf_1
X_21116_ _21115_/X VGND VGND VPWR VPWR _21116_/X sky130_fd_sc_hd__buf_2
XFILLER_59_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22096_ _22108_/A VGND VGND VPWR VPWR _22096_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23495__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21559__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21047_ _20819_/X _21044_/X _24039_/Q _21041_/X VGND VGND VPWR VPWR _21047_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15706__A _15706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22220__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14610__A _14725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12820_ _12769_/A _12818_/X _12820_/C VGND VGND VPWR VPWR _12821_/C sky130_fd_sc_hd__and3_4
XFILLER_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13226__A _13243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12130__A _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22998_ _22998_/A _22998_/B VGND VGND VPWR VPWR _23000_/B sky130_fd_sc_hd__or2_4
XFILLER_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12751_ _12189_/X _12681_/X _12715_/X _12281_/X _12750_/X VGND VGND VPWR VPWR _12751_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ _21935_/A VGND VGND VPWR VPWR _21949_/X sky130_fd_sc_hd__buf_2
XFILLER_42_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16537__A _12011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21731__B2 _21687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11702_/A VGND VGND VPWR VPWR _16023_/A sky130_fd_sc_hd__buf_2
XANTENNA__15441__A _13631_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15477_/A _23916_/Q VGND VGND VPWR VPWR _15470_/X sky130_fd_sc_hd__or2_4
XANTENNA__24176__D _19760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _13056_/A VGND VGND VPWR VPWR _12682_/X sky130_fd_sc_hd__buf_2
XFILLER_54_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16256__B _16256_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _15643_/A _14421_/B _14421_/C VGND VGND VPWR VPWR _14422_/C sky130_fd_sc_hd__and3_4
XANTENNA__24120__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11633_/A VGND VGND VPWR VPWR _17285_/A sky130_fd_sc_hd__buf_2
X_23619_ _23270_/CLK _23619_/D VGND VGND VPWR VPWR _14773_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18174__D _18174_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22287__A2 _22286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17140_ _17130_/X _17134_/X _17815_/A _17139_/X VGND VGND VPWR VPWR _17140_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__21495__B1 _15177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14352_ _14367_/A VGND VGND VPWR VPWR _14397_/A sky130_fd_sc_hd__buf_2
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ _20427_/A IRQ[24] VGND VGND VPWR VPWR _11564_/X sky130_fd_sc_hd__and2_4
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _12255_/X VGND VGND VPWR VPWR _13303_/X sky130_fd_sc_hd__buf_2
XFILLER_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17071_ _17069_/A _17068_/Y _11632_/X _17070_/Y VGND VGND VPWR VPWR _17082_/B sky130_fd_sc_hd__a211o_4
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22039__A2 _22038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14283_ _14283_/A _14283_/B VGND VGND VPWR VPWR _14283_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24270__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16022_ _16039_/A VGND VGND VPWR VPWR _16063_/A sky130_fd_sc_hd__buf_2
X_13234_ _12350_/A _13234_/B _13233_/X VGND VGND VPWR VPWR _13235_/C sky130_fd_sc_hd__and3_4
XANTENNA__21798__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13165_ _12745_/A _13165_/B VGND VGND VPWR VPWR _13165_/X sky130_fd_sc_hd__or2_4
XANTENNA__19860__B1 _22017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12305__A _12713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12116_ _12115_/X VGND VGND VPWR VPWR _12116_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13096_ _13096_/A _13094_/X _13095_/X VGND VGND VPWR VPWR _13101_/B sky130_fd_sc_hd__and3_4
X_17973_ _17973_/A VGND VGND VPWR VPWR _17973_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12047_ _11921_/X VGND VGND VPWR VPWR _16698_/A sky130_fd_sc_hd__buf_2
X_16924_ _16923_/X VGND VGND VPWR VPWR _16924_/X sky130_fd_sc_hd__buf_2
X_19712_ _19712_/A HRDATA[5] VGND VGND VPWR VPWR _19712_/X sky130_fd_sc_hd__and2_4
XFILLER_61_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16855_ _13776_/X _16854_/X _13776_/X _16854_/X VGND VGND VPWR VPWR _16855_/X sky130_fd_sc_hd__a2bb2o_4
X_19643_ _19643_/A _19643_/B VGND VGND VPWR VPWR _19806_/C sky130_fd_sc_hd__and2_4
XFILLER_4_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15806_ _12852_/A _15861_/B VGND VGND VPWR VPWR _15806_/X sky130_fd_sc_hd__or2_4
XANTENNA__13136__A _13059_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19574_ _19481_/A _19659_/A _19573_/Y VGND VGND VPWR VPWR _19629_/B sky130_fd_sc_hd__o21a_4
X_16786_ _16757_/X _16784_/X _16786_/C VGND VGND VPWR VPWR _16787_/C sky130_fd_sc_hd__and3_4
XFILLER_92_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13998_ _13998_/A VGND VGND VPWR VPWR _14065_/A sky130_fd_sc_hd__buf_2
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23218__CLK _23155_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22449__A _22134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18525_ _18137_/A _18525_/B VGND VGND VPWR VPWR _18525_/X sky130_fd_sc_hd__and2_4
X_15737_ _15750_/A _15737_/B VGND VGND VPWR VPWR _15737_/X sky130_fd_sc_hd__or2_4
XANTENNA__19915__B2 _20844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12949_ _12949_/A _23667_/Q VGND VGND VPWR VPWR _12951_/B sky130_fd_sc_hd__or2_4
XFILLER_45_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12975__A _12951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16447__A _16447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21722__B2 _21716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18456_ _18340_/X _18454_/X _18377_/X _18455_/X VGND VGND VPWR VPWR _18456_/X sky130_fd_sc_hd__o22a_4
XFILLER_34_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15668_ _15687_/A _15668_/B _15667_/X VGND VGND VPWR VPWR _15668_/X sky130_fd_sc_hd__and3_4
XFILLER_59_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17407_ _14073_/X _17407_/B VGND VGND VPWR VPWR _17407_/X sky130_fd_sc_hd__or2_4
XFILLER_18_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14619_ _13927_/A VGND VGND VPWR VPWR _14756_/A sky130_fd_sc_hd__buf_2
XANTENNA__15070__B _23551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18387_ _18264_/A _18387_/B VGND VGND VPWR VPWR _18390_/B sky130_fd_sc_hd__and2_4
XANTENNA__19679__B1 _11599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22278__A2 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15599_ _14379_/A _23563_/Q VGND VGND VPWR VPWR _15599_/X sky130_fd_sc_hd__or2_4
XFILLER_119_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17338_ _14425_/A _17313_/B _17316_/Y _17337_/Y VGND VGND VPWR VPWR _17338_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17278__A _17277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17269_ _17785_/B VGND VGND VPWR VPWR _17270_/B sky130_fd_sc_hd__inv_2
XFILLER_119_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24328__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16901__A1 _16524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19008_ _19008_/A VGND VGND VPWR VPWR _19008_/Y sky130_fd_sc_hd__inv_2
X_20280_ _20511_/A VGND VGND VPWR VPWR _20280_/X sky130_fd_sc_hd__buf_2
XANTENNA__22450__A2 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_47_0_HCLK clkbuf_5_23_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23970_ _24066_/CLK _23970_/D VGND VGND VPWR VPWR _15267_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_99_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22921_ _23027_/A _22921_/B VGND VGND VPWR VPWR _22921_/X sky130_fd_sc_hd__and2_4
XFILLER_84_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24110__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13046__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21961__B2 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22852_ _22852_/A VGND VGND VPWR VPWR HWDATA[23] sky130_fd_sc_hd__inv_2
XANTENNA__18556__B _16996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_21803_ _21802_/X _21793_/X _23609_/Q _21800_/X VGND VGND VPWR VPWR _23609_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19906__B2 _20317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22783_ _15051_/X _22782_/X VGND VGND VPWR VPWR HWDATA[0] sky130_fd_sc_hd__nor2_4
XFILLER_25_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15261__A _11909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21713__B2 _21709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22910__B1 _22924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21734_ _20199_/A _21734_/B VGND VGND VPWR VPWR _21734_/X sky130_fd_sc_hd__or2_4
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24453_ _24199_/CLK _18628_/Y HRESETn VGND VGND VPWR VPWR _24453_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19668__A _19800_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21665_ _21548_/X _21662_/X _15504_/B _21659_/X VGND VGND VPWR VPWR _23692_/D sky130_fd_sc_hd__o22a_4
XFILLER_36_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24293__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23404_ _23404_/CLK _22182_/X VGND VGND VPWR VPWR _23404_/Q sky130_fd_sc_hd__dfxtp_4
X_20616_ _20290_/X VGND VGND VPWR VPWR _20616_/X sky130_fd_sc_hd__buf_2
X_21596_ _21514_/X _21591_/X _16384_/B _21595_/X VGND VGND VPWR VPWR _21596_/X sky130_fd_sc_hd__o22a_4
X_24384_ _24425_/CLK _24384_/D HRESETn VGND VGND VPWR VPWR _24384_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12109__B _23709_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20547_ _18283_/X _20447_/X _20492_/X _20546_/Y VGND VGND VPWR VPWR _20547_/X sky130_fd_sc_hd__a211o_4
X_23335_ _23079_/CLK _23335_/D VGND VGND VPWR VPWR _23335_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18893__A1 _17181_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14605__A _11976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20478_ _20292_/X _20477_/X _24309_/Q _20305_/X VGND VGND VPWR VPWR _20479_/B sky130_fd_sc_hd__o22a_4
X_23266_ _23522_/CLK _23266_/D VGND VGND VPWR VPWR _15263_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22217_ _22091_/X _22215_/X _16211_/B _22212_/X VGND VGND VPWR VPWR _23383_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23197_ _24059_/CLK _22523_/X VGND VGND VPWR VPWR _12128_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22441__A2 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22148_ _22147_/X _22101_/A _23423_/Q _22071_/X VGND VGND VPWR VPWR _22148_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20342__A _20342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11964__A _11997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15436__A _15436_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14970_ _14970_/A _14909_/B VGND VGND VPWR VPWR _14970_/X sky130_fd_sc_hd__or2_4
X_22079_ _20338_/A VGND VGND VPWR VPWR _22079_/X sky130_fd_sc_hd__buf_2
XFILLER_0_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13921_ _13837_/X _13921_/B VGND VGND VPWR VPWR _13922_/A sky130_fd_sc_hd__or2_4
XFILLER_47_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15155__B _23873_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16640_ _11823_/A VGND VGND VPWR VPWR _16640_/X sky130_fd_sc_hd__buf_2
X_13852_ _13895_/A _23719_/Q VGND VGND VPWR VPWR _13852_/X sky130_fd_sc_hd__or2_4
XANTENNA__22269__A _22269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12803_ _12803_/A _12803_/B VGND VGND VPWR VPWR _12804_/C sky130_fd_sc_hd__or2_4
XFILLER_1_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21173__A _21165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16571_ _16567_/A _16654_/B VGND VGND VPWR VPWR _16573_/B sky130_fd_sc_hd__or2_4
X_13783_ _15398_/A _13783_/B _13782_/X VGND VGND VPWR VPWR _13783_/X sky130_fd_sc_hd__or3_4
XANTENNA__12795__A _12795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18310_ _18171_/X _18293_/X _18202_/X _18309_/X VGND VGND VPWR VPWR _18310_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21704__B2 _21702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15522_ _12233_/X _15522_/B VGND VGND VPWR VPWR _15522_/X sky130_fd_sc_hd__or2_4
X_12734_ _12747_/A VGND VGND VPWR VPWR _12737_/A sky130_fd_sc_hd__buf_2
X_19290_ _24259_/Q _19208_/B _19289_/Y VGND VGND VPWR VPWR _24259_/D sky130_fd_sc_hd__o21a_4
XFILLER_76_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23510__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18241_ _18241_/A _17524_/B VGND VGND VPWR VPWR _18241_/Y sky130_fd_sc_hd__nor2_4
X_15453_ _15453_/A VGND VGND VPWR VPWR _15453_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21901__A _21901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12665_ _12953_/A _24085_/Q VGND VGND VPWR VPWR _12666_/C sky130_fd_sc_hd__or2_4
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _15589_/A _14404_/B _14404_/C VGND VGND VPWR VPWR _14404_/X sky130_fd_sc_hd__or3_4
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21468__B1 _12658_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _11615_/X VGND VGND VPWR VPWR _13595_/A sky130_fd_sc_hd__buf_2
X_18172_ _16945_/Y _16982_/X _18132_/C VGND VGND VPWR VPWR _18172_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ _15384_/A VGND VGND VPWR VPWR _15384_/Y sky130_fd_sc_hd__inv_2
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _12596_/A _12592_/X _12596_/C VGND VGND VPWR VPWR _12596_/X sky130_fd_sc_hd__and3_4
XANTENNA__18333__B1 _18160_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19676__A3 _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17123_ _15120_/Y _17010_/A _17018_/A _17122_/X VGND VGND VPWR VPWR _17160_/A sky130_fd_sc_hd__o22a_4
X_14335_ _11977_/X _14307_/X _14314_/X _14326_/X _14334_/X VGND VGND VPWR VPWR _14335_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11547_ _11544_/X _11547_/B VGND VGND VPWR VPWR _20071_/B sky130_fd_sc_hd__or2_4
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22680__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17054_ _17054_/A _17068_/A _11591_/D _11601_/A VGND VGND VPWR VPWR _17054_/X sky130_fd_sc_hd__or4_4
X_14266_ _14174_/X _14263_/X _14265_/Y VGND VGND VPWR VPWR _14267_/B sky130_fd_sc_hd__a21o_4
XFILLER_13_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16005_ _11851_/X _16004_/X VGND VGND VPWR VPWR _16005_/X sky130_fd_sc_hd__and2_4
X_13217_ _13231_/A _13217_/B _13216_/X VGND VGND VPWR VPWR _13218_/C sky130_fd_sc_hd__and3_4
XFILLER_98_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14197_ _14197_/A VGND VGND VPWR VPWR _14204_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20443__B2 _20374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13148_ _15685_/A _24017_/Q VGND VGND VPWR VPWR _13150_/B sky130_fd_sc_hd__or2_4
XFILLER_97_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11874__A _16147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15346__A _14020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13079_ _13065_/A VGND VGND VPWR VPWR _13080_/A sky130_fd_sc_hd__buf_2
X_17956_ _17090_/X VGND VGND VPWR VPWR _18265_/A sky130_fd_sc_hd__buf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14250__A _13686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22196__B2 _22190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16907_ _16916_/A _16916_/B _16907_/C _16906_/Y VGND VGND VPWR VPWR _16907_/X sky130_fd_sc_hd__or4_4
X_17887_ _11628_/X VGND VGND VPWR VPWR _18129_/A sky130_fd_sc_hd__buf_2
XFILLER_65_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21943__A1 _21823_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20746__A2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18657__A _17090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17561__A _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21943__B2 _21942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19626_ _19625_/Y _19638_/A _19500_/X _19622_/Y VGND VGND VPWR VPWR _19626_/X sky130_fd_sc_hd__o22a_4
XFILLER_96_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16838_ _15915_/X _16835_/X _15920_/Y VGND VGND VPWR VPWR _16838_/X sky130_fd_sc_hd__o21a_4
XFILLER_65_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22179__A _22172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16769_ _16768_/X _16708_/B VGND VGND VPWR VPWR _16769_/X sky130_fd_sc_hd__or2_4
X_19557_ _24151_/Q _19435_/A HRDATA[25] _19431_/X VGND VGND VPWR VPWR _19557_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22499__A2 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18508_ _18224_/A VGND VGND VPWR VPWR _18508_/X sky130_fd_sc_hd__buf_2
XFILLER_34_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19488_ _19499_/A VGND VGND VPWR VPWR _19537_/A sky130_fd_sc_hd__buf_2
XFILLER_62_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22907__A _22899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21171__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14409__B _14330_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18439_ _18438_/X VGND VGND VPWR VPWR _18439_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18392__A _18392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21450_ _21449_/X VGND VGND VPWR VPWR _21455_/A sky130_fd_sc_hd__buf_2
XANTENNA__21459__B1 _23803_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20401_ _20229_/X _20400_/X _20213_/X VGND VGND VPWR VPWR _20401_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_4_10_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21381_ _21265_/X _21376_/X _15577_/B _21380_/X VGND VGND VPWR VPWR _23851_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17678__A2 _17506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14425__A _14425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20332_ _20332_/A _20331_/X VGND VGND VPWR VPWR _20332_/Y sky130_fd_sc_hd__nor2_4
X_23120_ _23473_/CLK _23120_/D VGND VGND VPWR VPWR _13325_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_31_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19935__B _19927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23051_ _23051_/A _16993_/X VGND VGND VPWR VPWR _23053_/B sky130_fd_sc_hd__or2_4
X_20263_ _20251_/X _20262_/X _19235_/Y _20251_/X VGND VGND VPWR VPWR _20263_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17736__A _17736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16640__A _11823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22002_ _22002_/A VGND VGND VPWR VPWR _22002_/X sky130_fd_sc_hd__buf_2
XFILLER_118_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13983__B _23690_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20194_ _20194_/A _11634_/B _16929_/B _20206_/A VGND VGND VPWR VPWR _20195_/D sky130_fd_sc_hd__or4_4
XFILLER_89_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11784__A _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14160__A _15030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22187__B2 _22183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23953_ _24082_/CLK _23953_/D VGND VGND VPWR VPWR _23953_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18567__A _18137_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21934__B2 _21928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22904_ _22899_/X _22902_/X _22904_/C VGND VGND VPWR VPWR _22904_/X sky130_fd_sc_hd__and3_4
XANTENNA__17471__A _12676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23533__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23884_ _23794_/CLK _23884_/D VGND VGND VPWR VPWR _23884_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22089__A _22101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22835_ _17115_/Y _22826_/X _22827_/X VGND VGND VPWR VPWR _22835_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16087__A _13447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13504__A _15892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22766_ _22744_/Y _22765_/B VGND VGND VPWR VPWR _22768_/A sky130_fd_sc_hd__or2_4
XFILLER_0_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17366__A1 _16800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21717_ _21550_/X _21712_/X _23659_/Q _21716_/X VGND VGND VPWR VPWR _23659_/D sky130_fd_sc_hd__o22a_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22697_ _22683_/A VGND VGND VPWR VPWR _22697_/X sky130_fd_sc_hd__buf_2
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _12450_/A VGND VGND VPWR VPWR _12494_/A sky130_fd_sc_hd__buf_2
X_24436_ _23358_/CLK _24436_/D HRESETn VGND VGND VPWR VPWR _24436_/Q sky130_fd_sc_hd__dfrtp_4
X_21648_ _21662_/A VGND VGND VPWR VPWR _21648_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17118__A1 _17115_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17118__B2 _17117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22111__B2 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11959__A _13428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ _12381_/A _12248_/B VGND VGND VPWR VPWR _12382_/C sky130_fd_sc_hd__or2_4
X_24367_ _24334_/CLK _24367_/D HRESETn VGND VGND VPWR VPWR _24367_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22662__A2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21579_ _21578_/X _21532_/A _23743_/Q _21515_/A VGND VGND VPWR VPWR _23743_/D sky130_fd_sc_hd__o22a_4
X_14120_ _15010_/A VGND VGND VPWR VPWR _14121_/A sky130_fd_sc_hd__buf_2
X_23318_ _24082_/CLK _22308_/X VGND VGND VPWR VPWR _12259_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18170__A2_N _18169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24298_ _24299_/CLK _24298_/D HRESETn VGND VGND VPWR VPWR _24298_/Q sky130_fd_sc_hd__dfrtp_4
X_14051_ _14031_/A _13969_/B VGND VGND VPWR VPWR _14053_/B sky130_fd_sc_hd__or2_4
XANTENNA__24374__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23249_ _23217_/CLK _23249_/D VGND VGND VPWR VPWR _13137_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22414__A2 _22404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13002_ _12886_/A _23730_/Q VGND VGND VPWR VPWR _13002_/X sky130_fd_sc_hd__or2_4
XANTENNA__21168__A _21168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20072__A _20071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_30_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_30_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17810_ _17801_/X _17805_/X _17807_/X _17809_/X VGND VGND VPWR VPWR _17810_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_79_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18790_ _13575_/X _18788_/X _24431_/Q _18789_/X VGND VGND VPWR VPWR _24431_/D sky130_fd_sc_hd__o22a_4
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14070__A _14847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12115__B1 _11599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22178__B2 _22176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17741_ _17735_/A _17117_/X _17735_/X _17740_/X VGND VGND VPWR VPWR _17741_/X sky130_fd_sc_hd__o22a_4
X_14953_ _14243_/A _14953_/B _14953_/C VGND VGND VPWR VPWR _14953_/X sky130_fd_sc_hd__and3_4
XANTENNA__20800__A _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21925__B2 _21921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13904_ _13880_/A _13904_/B _13903_/X VGND VGND VPWR VPWR _13904_/X sky130_fd_sc_hd__and3_4
X_17672_ _17672_/A _17497_/X VGND VGND VPWR VPWR _17677_/A sky130_fd_sc_hd__and2_4
X_14884_ _11606_/A _14882_/X _14883_/X VGND VGND VPWR VPWR _14884_/X sky130_fd_sc_hd__and3_4
XFILLER_29_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16623_ _16597_/X _16612_/X _16623_/C VGND VGND VPWR VPWR _16646_/B sky130_fd_sc_hd__and3_4
X_19411_ _19302_/X VGND VGND VPWR VPWR _19411_/X sky130_fd_sc_hd__buf_2
X_13835_ _15450_/A _13834_/X VGND VGND VPWR VPWR _13835_/X sky130_fd_sc_hd__and2_4
XFILLER_63_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16554_ _16689_/A _16554_/B _16553_/X VGND VGND VPWR VPWR _16554_/X sky130_fd_sc_hd__or3_4
X_19342_ _19340_/X _18510_/X _19340_/X _20743_/A VGND VGND VPWR VPWR _24234_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13766_ _12650_/A _13766_/B VGND VGND VPWR VPWR _13766_/X sky130_fd_sc_hd__or2_4
XANTENNA__21153__A2 _21147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15505_ _15512_/A _23852_/Q VGND VGND VPWR VPWR _15506_/C sky130_fd_sc_hd__or2_4
XFILLER_31_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12717_ _12709_/A VGND VGND VPWR VPWR _12720_/A sky130_fd_sc_hd__buf_2
X_19273_ _19217_/B VGND VGND VPWR VPWR _19273_/Y sky130_fd_sc_hd__inv_2
X_16485_ _16471_/X _23610_/Q VGND VGND VPWR VPWR _16487_/B sky130_fd_sc_hd__or2_4
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13697_ _13718_/A VGND VGND VPWR VPWR _13697_/X sky130_fd_sc_hd__buf_2
X_18224_ _18224_/A VGND VGND VPWR VPWR _18224_/X sky130_fd_sc_hd__buf_2
X_15436_ _15436_/A _23468_/Q VGND VGND VPWR VPWR _15438_/B sky130_fd_sc_hd__or2_4
XFILLER_19_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12648_ _12640_/A _12648_/B VGND VGND VPWR VPWR _12648_/X sky130_fd_sc_hd__or2_4
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18306__B1 _18189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22102__A1 _22100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20247__A _20453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22102__B2 _22096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18155_ _18254_/A _18154_/X _17524_/Y VGND VGND VPWR VPWR _18155_/X sky130_fd_sc_hd__o21a_4
X_15367_ _12567_/A _15307_/B VGND VGND VPWR VPWR _15368_/C sky130_fd_sc_hd__or2_4
XANTENNA__18857__A1 _14564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12579_ _12935_/A VGND VGND VPWR VPWR _12980_/A sky130_fd_sc_hd__buf_2
XFILLER_50_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22653__A2 _22650_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18940__A _18940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17106_ _21005_/A _17032_/B _13594_/X _17105_/X VGND VGND VPWR VPWR _17106_/X sky130_fd_sc_hd__o22a_4
XFILLER_7_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20664__A1 _18430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14318_ _14318_/A VGND VGND VPWR VPWR _15574_/A sky130_fd_sc_hd__buf_2
XFILLER_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18086_ _18085_/A _18085_/B _17998_/X VGND VGND VPWR VPWR _18086_/Y sky130_fd_sc_hd__a21oi_4
X_15298_ _12449_/A _15296_/X _15297_/X VGND VGND VPWR VPWR _15298_/X sky130_fd_sc_hd__and3_4
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_112_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR _23539_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23406__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22462__A _21001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17037_ _18864_/C _17032_/X _17105_/B VGND VGND VPWR VPWR _17037_/Y sky130_fd_sc_hd__o21ai_4
X_14249_ _14345_/A _14249_/B _14249_/C VGND VGND VPWR VPWR _14249_/X sky130_fd_sc_hd__and3_4
XANTENNA__17556__A _16077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22405__A2 _22404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14899__B _14899_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15076__A _15114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23556__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18988_ _19002_/A VGND VGND VPWR VPWR _18988_/X sky130_fd_sc_hd__buf_2
XFILLER_86_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15843__A1 _12716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17939_ _17794_/A _17932_/Y _17933_/X _17938_/Y VGND VGND VPWR VPWR _17939_/X sky130_fd_sc_hd__a211o_4
XFILLER_113_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15804__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20950_ _20493_/A _20949_/X _19110_/A _20500_/A VGND VGND VPWR VPWR _20950_/X sky130_fd_sc_hd__o22a_4
XFILLER_96_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21392__A2 _21390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19609_ _19629_/A _19597_/A _19629_/B VGND VGND VPWR VPWR _19609_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15523__B _23499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20881_ _24388_/Q _20405_/A _24420_/Q _20682_/X VGND VGND VPWR VPWR _20881_/X sky130_fd_sc_hd__o22a_4
XFILLER_42_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22620_ _22614_/Y _22619_/X _22388_/X _22619_/X VGND VGND VPWR VPWR _22620_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13324__A _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22341__B2 _22337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13043__B _24082_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22551_ _22439_/X _22550_/X _23177_/Q _22547_/X VGND VGND VPWR VPWR _22551_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16635__A _16622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21502_ _21527_/A VGND VGND VPWR VPWR _21515_/A sky130_fd_sc_hd__buf_2
X_22482_ _22408_/X _22479_/X _12323_/B _22476_/X VGND VGND VPWR VPWR _22482_/X sky130_fd_sc_hd__o22a_4
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24221_ _24187_/CLK _19366_/X HRESETn VGND VGND VPWR VPWR _24221_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11779__A _11821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21433_ _21400_/A VGND VGND VPWR VPWR _21433_/X sky130_fd_sc_hd__buf_2
XANTENNA__22644__A2 _22643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21364_ _21237_/X _21362_/X _16220_/B _21359_/X VGND VGND VPWR VPWR _23863_/D sky130_fd_sc_hd__o22a_4
X_24152_ _24223_/CLK _24152_/D HRESETn VGND VGND VPWR VPWR _24152_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23086__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22372__A _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20315_ _21791_/A VGND VGND VPWR VPWR _20315_/X sky130_fd_sc_hd__buf_2
X_23103_ _23889_/CLK _22663_/X VGND VGND VPWR VPWR _23103_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13994__A _14010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17466__A _12559_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21295_ _23902_/Q VGND VGND VPWR VPWR _21295_/Y sky130_fd_sc_hd__inv_2
X_24083_ _23987_/CLK _20538_/X VGND VGND VPWR VPWR _12909_/B sky130_fd_sc_hd__dfxtp_4
X_20246_ _20525_/A VGND VGND VPWR VPWR _20453_/A sky130_fd_sc_hd__buf_2
X_23034_ _23018_/A _23032_/Y _23033_/X VGND VGND VPWR VPWR _23034_/X sky130_fd_sc_hd__and3_4
XFILLER_46_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21604__B1 _12768_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21080__B2 _21079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_17_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20177_ _20132_/Y _19936_/X _20176_/X VGND VGND VPWR VPWR _20177_/X sky130_fd_sc_hd__o21a_4
XFILLER_44_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21716__A _21702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18297__A _18297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21907__B2 _21905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15714__A _13129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11950_ _11996_/A _21683_/A VGND VGND VPWR VPWR _11965_/B sky130_fd_sc_hd__or2_4
X_23936_ _23104_/CLK _23936_/D VGND VGND VPWR VPWR _14889_/B sky130_fd_sc_hd__dfxtp_4
X_11881_ _14283_/A VGND VGND VPWR VPWR _15706_/A sky130_fd_sc_hd__buf_2
X_23867_ _23867_/CLK _21358_/X VGND VGND VPWR VPWR _23867_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13620_ _13620_/A _13713_/B VGND VGND VPWR VPWR _13621_/C sky130_fd_sc_hd__or2_4
XANTENNA__13234__A _12350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22818_ _22821_/A _14493_/Y VGND VGND VPWR VPWR _22818_/X sky130_fd_sc_hd__or2_4
XFILLER_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23798_ _23473_/CLK _23798_/D VGND VGND VPWR VPWR _12329_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21135__A2 _21133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22547__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13551_ _12980_/A VGND VGND VPWR VPWR _13551_/X sky130_fd_sc_hd__buf_2
X_22749_ SYSTICKCLKDIV[0] _22750_/A _22748_/Y VGND VGND VPWR VPWR _24095_/D sky130_fd_sc_hd__o21a_4
XFILLER_34_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12502_ _12540_/A _12502_/B _12501_/X VGND VGND VPWR VPWR _12502_/X sky130_fd_sc_hd__and3_4
XANTENNA__20894__A1 _20872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16270_ _11980_/X _16269_/X VGND VGND VPWR VPWR _16270_/X sky130_fd_sc_hd__and2_4
XFILLER_51_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13482_ _13442_/X _13480_/X _13482_/C VGND VGND VPWR VPWR _13483_/C sky130_fd_sc_hd__and3_4
XFILLER_16_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20894__B2 _20839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16264__B _23577_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15221_ _14186_/A _23585_/Q VGND VGND VPWR VPWR _15221_/X sky130_fd_sc_hd__or2_4
XFILLER_90_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12433_ _12432_/X VGND VGND VPWR VPWR _12433_/Y sky130_fd_sc_hd__inv_2
X_24419_ _24320_/CLK _24419_/D HRESETn VGND VGND VPWR VPWR _20901_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18839__A1 _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11689__A _12837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22635__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17079__C _18728_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18760__A _17040_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15152_ _14119_/X _15148_/X _15151_/X VGND VGND VPWR VPWR _15153_/B sky130_fd_sc_hd__or3_4
X_12364_ _13133_/A _12354_/X _12364_/C VGND VGND VPWR VPWR _12364_/X sky130_fd_sc_hd__and3_4
XANTENNA__24213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14103_ _14992_/A VGND VGND VPWR VPWR _14315_/A sky130_fd_sc_hd__buf_2
X_15083_ _15107_/A _15083_/B _15083_/C VGND VGND VPWR VPWR _15084_/C sky130_fd_sc_hd__and3_4
X_19960_ _19960_/A VGND VGND VPWR VPWR _19960_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12295_ _12695_/A _12293_/X _12294_/X VGND VGND VPWR VPWR _12295_/X sky130_fd_sc_hd__and3_4
X_14034_ _11647_/A _22320_/A VGND VGND VPWR VPWR _14036_/B sky130_fd_sc_hd__or2_4
X_18911_ _14425_/A _18905_/X _19072_/A _18906_/X VGND VGND VPWR VPWR _24358_/D sky130_fd_sc_hd__o22a_4
XFILLER_113_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17095__B _18421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19891_ _20218_/A VGND VGND VPWR VPWR _20849_/B sky130_fd_sc_hd__buf_2
XFILLER_79_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18842_ _18842_/A VGND VGND VPWR VPWR _18842_/X sky130_fd_sc_hd__buf_2
XFILLER_84_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21071__B2 _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21626__A _21590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15985_ _15957_/A _23416_/Q VGND VGND VPWR VPWR _15986_/C sky130_fd_sc_hd__or2_4
X_18773_ _16514_/X _18765_/X _24442_/Q _18768_/X VGND VGND VPWR VPWR _18773_/X sky130_fd_sc_hd__o22a_4
XFILLER_114_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14936_ _12340_/A _14879_/B VGND VGND VPWR VPWR _14938_/B sky130_fd_sc_hd__or2_4
X_17724_ _17720_/A VGND VGND VPWR VPWR _17724_/X sky130_fd_sc_hd__buf_2
XFILLER_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17578__A1 _16814_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17578__B2 _17577_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21374__A2 _21369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14867_ _14880_/A VGND VGND VPWR VPWR _14867_/X sky130_fd_sc_hd__buf_2
X_17655_ _17652_/A _17652_/B VGND VGND VPWR VPWR _17658_/A sky130_fd_sc_hd__or2_4
XANTENNA__13144__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_37_0_HCLK clkbuf_6_18_0_HCLK/X VGND VGND VPWR VPWR _23557_/CLK sky130_fd_sc_hd__clkbuf_1
X_13818_ _13630_/A _23399_/Q VGND VGND VPWR VPWR _13819_/C sky130_fd_sc_hd__or2_4
X_16606_ _11748_/X VGND VGND VPWR VPWR _16616_/A sky130_fd_sc_hd__buf_2
XFILLER_56_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17586_ _17447_/X _17455_/X _17586_/C _18152_/A VGND VGND VPWR VPWR _17590_/A sky130_fd_sc_hd__or4_4
XANTENNA__11590__C _17040_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14798_ _13862_/A _14798_/B VGND VGND VPWR VPWR _14798_/X sky130_fd_sc_hd__or2_4
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16537_ _12011_/A _16537_/B _16537_/C VGND VGND VPWR VPWR _16542_/B sky130_fd_sc_hd__and3_4
X_19325_ _19328_/A VGND VGND VPWR VPWR _19325_/X sky130_fd_sc_hd__buf_2
X_13749_ _13697_/X _13662_/B VGND VGND VPWR VPWR _13749_/X sky130_fd_sc_hd__or2_4
XFILLER_71_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16455__A _11702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16468_ _16159_/X _16408_/B VGND VGND VPWR VPWR _16468_/X sky130_fd_sc_hd__or2_4
X_19256_ _19225_/A _19257_/A _19255_/Y VGND VGND VPWR VPWR _24276_/D sky130_fd_sc_hd__o21a_4
X_15419_ _13647_/A _15419_/B _15419_/C VGND VGND VPWR VPWR _15419_/X sky130_fd_sc_hd__or3_4
X_18207_ _18266_/A _17452_/X VGND VGND VPWR VPWR _18207_/X sky130_fd_sc_hd__and2_4
XANTENNA__11599__A _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22087__B1 _16267_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19187_ _19116_/B VGND VGND VPWR VPWR _19187_/Y sky130_fd_sc_hd__inv_2
X_16399_ _16083_/A _16396_/X _16398_/X VGND VGND VPWR VPWR _16399_/X sky130_fd_sc_hd__and3_4
Xclkbuf_3_6_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18138_ _18266_/A _18138_/B VGND VGND VPWR VPWR _18139_/D sky130_fd_sc_hd__and2_4
XFILLER_105_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18069_ _17824_/X _17820_/Y _17812_/A _17829_/Y VGND VGND VPWR VPWR _18069_/X sky130_fd_sc_hd__o22a_4
X_20100_ _20099_/Y _11538_/X _11553_/X VGND VGND VPWR VPWR _20100_/Y sky130_fd_sc_hd__a21oi_4
X_21080_ _20487_/X _21075_/X _24021_/Q _21079_/X VGND VGND VPWR VPWR _21080_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15518__B _15517_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22920__A _22899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20031_ _20018_/X _17893_/X _20024_/X _20030_/X VGND VGND VPWR VPWR _20031_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12223__A _12211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21536__A _20574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21982_ _21804_/X _21981_/X _23512_/Q _21978_/X VGND VGND VPWR VPWR _23512_/D sky130_fd_sc_hd__o22a_4
XFILLER_96_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21365__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22562__B2 _22518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23721_ _23978_/CLK _23721_/D VGND VGND VPWR VPWR _23721_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20933_ _20283_/X _20924_/Y _20931_/X _20932_/Y _20459_/A VGND VGND VPWR VPWR _20933_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_76_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15253__B _15253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13054__A _13054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ _23363_/CLK _21727_/X VGND VGND VPWR VPWR _14679_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ _20864_/A VGND VGND VPWR VPWR _20864_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22603_ _22444_/X _22600_/X _13873_/B _22597_/X VGND VGND VPWR VPWR _22603_/X sky130_fd_sc_hd__o22a_4
XFILLER_74_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23583_ _23487_/CLK _23583_/D VGND VGND VPWR VPWR _23583_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20795_ _24200_/Q _20751_/X _20794_/Y VGND VGND VPWR VPWR _22127_/A sky130_fd_sc_hd__o21a_4
XANTENNA__16365__A _16365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22534_ _22410_/X _22529_/X _12462_/B _22533_/X VGND VGND VPWR VPWR _22534_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16084__B _16158_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22078__B1 _12140_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22465_ _20199_/A _21784_/D VGND VGND VPWR VPWR _22465_/X sky130_fd_sc_hd__or2_4
XFILLER_6_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24204_ _24208_/CLK _19395_/X HRESETn VGND VGND VPWR VPWR _24204_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20628__A1 _20494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21416_ _21416_/A VGND VGND VPWR VPWR _21416_/X sky130_fd_sc_hd__buf_2
XFILLER_33_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22396_ _20355_/A VGND VGND VPWR VPWR _22396_/X sky130_fd_sc_hd__buf_2
XFILLER_68_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24135_ _24241_/CLK _24135_/D HRESETn VGND VGND VPWR VPWR _24135_/Q sky130_fd_sc_hd__dfrtp_4
X_21347_ _23870_/Q VGND VGND VPWR VPWR _21347_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15709__A _13004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14613__A _14146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12080_ _11999_/A _12080_/B _12080_/C VGND VGND VPWR VPWR _12081_/B sky130_fd_sc_hd__or3_4
X_24066_ _24066_/CLK _24066_/D VGND VGND VPWR VPWR _15297_/B sky130_fd_sc_hd__dfxtp_4
X_21278_ _21242_/A VGND VGND VPWR VPWR _21278_/X sky130_fd_sc_hd__buf_2
X_23017_ _18162_/X _23017_/B VGND VGND VPWR VPWR _23018_/C sky130_fd_sc_hd__or2_4
XFILLER_1_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21053__B2 _21048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20229_ _20229_/A VGND VGND VPWR VPWR _20229_/X sky130_fd_sc_hd__buf_2
XANTENNA__12133__A _12169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17643__B _17274_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23101__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11972__A _11966_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15770_ _15751_/A _15697_/B VGND VGND VPWR VPWR _15770_/X sky130_fd_sc_hd__or2_4
X_12982_ _12982_/A _12982_/B _12981_/X VGND VGND VPWR VPWR _12982_/X sky130_fd_sc_hd__and3_4
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24179__D _19717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14721_ _14640_/X _14723_/B VGND VGND VPWR VPWR _15387_/A sky130_fd_sc_hd__or2_4
XANTENNA__22553__B2 _22547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11933_ _12914_/A VGND VGND VPWR VPWR _11933_/X sky130_fd_sc_hd__buf_2
X_23919_ _23859_/CLK _23919_/D VGND VGND VPWR VPWR _13453_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15163__B _23809_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17440_ _12101_/X _17467_/B VGND VGND VPWR VPWR _17440_/X sky130_fd_sc_hd__and2_4
X_14652_ _14679_/A _14652_/B VGND VGND VPWR VPWR _14652_/X sky130_fd_sc_hd__or2_4
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11864_ _16113_/A VGND VGND VPWR VPWR _11924_/A sky130_fd_sc_hd__buf_2
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21108__A2 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13603_ _13603_/A VGND VGND VPWR VPWR _15404_/A sky130_fd_sc_hd__buf_2
X_17371_ _15782_/B _17371_/B VGND VGND VPWR VPWR _17371_/X sky130_fd_sc_hd__and2_4
XANTENNA__13899__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14583_ _15028_/A VGND VGND VPWR VPWR _14727_/A sky130_fd_sc_hd__buf_2
XANTENNA__24465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11795_ _16045_/A _11763_/X _11794_/X VGND VGND VPWR VPWR _11837_/B sky130_fd_sc_hd__or3_4
X_16322_ _16322_/A _16263_/B VGND VGND VPWR VPWR _16322_/X sky130_fd_sc_hd__or2_4
X_19110_ _19110_/A _19110_/B VGND VGND VPWR VPWR _19197_/A sky130_fd_sc_hd__and2_4
XFILLER_41_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13534_ _13562_/A _23535_/Q VGND VGND VPWR VPWR _13534_/X sky130_fd_sc_hd__or2_4
X_19041_ _24331_/Q VGND VGND VPWR VPWR _19041_/Y sky130_fd_sc_hd__inv_2
X_16253_ _16252_/X _16253_/B VGND VGND VPWR VPWR _16253_/X sky130_fd_sc_hd__or2_4
XFILLER_51_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13349__A2 _11618_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13465_ _13437_/X _23599_/Q VGND VGND VPWR VPWR _13467_/B sky130_fd_sc_hd__or2_4
XANTENNA__22608__A2 _22607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12308__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15204_ _14251_/A _15149_/B VGND VGND VPWR VPWR _15204_/X sky130_fd_sc_hd__or2_4
X_12416_ _12413_/X _12414_/X _12416_/C VGND VGND VPWR VPWR _12416_/X sky130_fd_sc_hd__and3_4
XFILLER_51_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16184_ _11700_/X VGND VGND VPWR VPWR _16185_/A sky130_fd_sc_hd__buf_2
X_13396_ _13395_/X _23600_/Q VGND VGND VPWR VPWR _13399_/B sky130_fd_sc_hd__or2_4
X_15135_ _11879_/A _15196_/B VGND VGND VPWR VPWR _15135_/X sky130_fd_sc_hd__or2_4
X_12347_ _12828_/A _12213_/B VGND VGND VPWR VPWR _12348_/C sky130_fd_sc_hd__or2_4
XANTENNA__21292__B2 _21230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15066_ _15104_/A _15064_/X _15065_/X VGND VGND VPWR VPWR _15066_/X sky130_fd_sc_hd__and3_4
X_19943_ _18066_/A _19943_/B VGND VGND VPWR VPWR _19944_/D sky130_fd_sc_hd__and2_4
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12278_ _13025_/A _12278_/B _12277_/X VGND VGND VPWR VPWR _12278_/X sky130_fd_sc_hd__or3_4
XANTENNA__22740__A SYSTICKCLKDIV[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19360__A2_N _18754_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14017_ _12599_/A _14017_/B _14016_/X VGND VGND VPWR VPWR _14018_/C sky130_fd_sc_hd__and3_4
XFILLER_96_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13139__A _15654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19874_ _19494_/X _19706_/A _19873_/X VGND VGND VPWR VPWR _19874_/X sky130_fd_sc_hd__o21a_4
XFILLER_64_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18825_ _17277_/X _18818_/X _24411_/Q _18821_/X VGND VGND VPWR VPWR _18825_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20260__A _20449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12978__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11882__A _15706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18756_ _18650_/X _18755_/X _24447_/Q _18650_/X VGND VGND VPWR VPWR _24447_/D sky130_fd_sc_hd__a2bb2o_4
X_15968_ _13477_/X VGND VGND VPWR VPWR _15997_/A sky130_fd_sc_hd__buf_2
XANTENNA__18748__B1 _17057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22544__B2 _22540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17707_ _17708_/A VGND VGND VPWR VPWR _18348_/A sky130_fd_sc_hd__buf_2
XFILLER_64_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14919_ _14177_/A VGND VGND VPWR VPWR _15063_/A sky130_fd_sc_hd__buf_2
X_15899_ _15892_/A _15829_/B VGND VGND VPWR VPWR _15900_/C sky130_fd_sc_hd__or2_4
X_18687_ _18684_/Y _18686_/X _18684_/Y _18686_/X VGND VGND VPWR VPWR _18687_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17638_ _16924_/X VGND VGND VPWR VPWR _17639_/A sky130_fd_sc_hd__buf_2
XFILLER_97_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14785__A1 _11841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17569_ _17569_/A _18047_/A _18085_/A _17568_/Y VGND VGND VPWR VPWR _17569_/X sky130_fd_sc_hd__or4_4
XFILLER_17_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16185__A _16185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19308_ _19308_/A VGND VGND VPWR VPWR _19308_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13602__A _14778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20580_ _20448_/X _20579_/X _24368_/Q _20407_/X VGND VGND VPWR VPWR _20580_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24135__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22915__A _23038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19239_ _19234_/B VGND VGND VPWR VPWR _19239_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19496__A _19545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12218__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19927__C _18812_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22250_ _11732_/B VGND VGND VPWR VPWR _22250_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17728__B _17300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21201_ _21180_/A VGND VGND VPWR VPWR _21201_/X sky130_fd_sc_hd__buf_2
X_22181_ _22115_/X _22179_/X _15825_/B _22176_/X VGND VGND VPWR VPWR _22181_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15529__A _12257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22480__B1 _15992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14433__A _15571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21132_ _20509_/X _21126_/X _23988_/Q _21130_/X VGND VGND VPWR VPWR _21132_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23024__A2 _16985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22650__A _22621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21063_ _21067_/A VGND VGND VPWR VPWR _21079_/A sky130_fd_sc_hd__inv_2
XFILLER_87_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23124__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13049__A _13022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21035__B2 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20014_ _24466_/Q VGND VGND VPWR VPWR _20014_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21266__A _21242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20170__A _18940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12888__A _12518_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11792__A _11823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15264__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22535__A1 _22413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21338__A2 _21333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16079__B _16077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22535__B2 _22533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21965_ _21863_/X _21938_/A _23519_/Q _21920_/X VGND VGND VPWR VPWR _23519_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19400__B2 _24201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12400__B _12293_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23704_ _23316_/CLK _23704_/D VGND VGND VPWR VPWR _23704_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_76_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _21855_/A VGND VGND VPWR VPWR _20916_/X sky130_fd_sc_hd__buf_2
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21896_ _21831_/X _21894_/X _15861_/B _21891_/X VGND VGND VPWR VPWR _21896_/X sky130_fd_sc_hd__o22a_4
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_20_0_HCLK clkbuf_6_10_0_HCLK/X VGND VGND VPWR VPWR _24223_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23635_/CLK _21756_/X VGND VGND VPWR VPWR _12912_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_74_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22299__B1 _15056_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _20846_/X VGND VGND VPWR VPWR _20847_/X sky130_fd_sc_hd__buf_2
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16095__A _16095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14608__A _14143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_83_0_HCLK clkbuf_7_82_0_HCLK/A VGND VGND VPWR VPWR _24334_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13512__A _12591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ _17024_/A VGND VGND VPWR VPWR _11580_/Y sky130_fd_sc_hd__inv_2
X_23566_ _23564_/CLK _21895_/X VGND VGND VPWR VPWR _15674_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_22_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20778_ _20778_/A VGND VGND VPWR VPWR _21555_/A sky130_fd_sc_hd__buf_2
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22517_ _22521_/A VGND VGND VPWR VPWR _22533_/A sky130_fd_sc_hd__inv_2
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23497_ _23561_/CLK _22003_/X VGND VGND VPWR VPWR _23497_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13250_ _12350_/A _13248_/X _13250_/C VGND VGND VPWR VPWR _13251_/C sky130_fd_sc_hd__and3_4
XFILLER_52_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22448_ _22446_/X _22440_/X _14268_/B _22447_/X VGND VGND VPWR VPWR _23238_/D sky130_fd_sc_hd__o22a_4
XFILLER_100_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12201_ _13983_/A VGND VGND VPWR VPWR _12202_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15439__A _15436_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11967__A _11886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21274__A1 _21273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13181_ _15696_/A _13181_/B VGND VGND VPWR VPWR _13181_/X sky130_fd_sc_hd__or2_4
XANTENNA__21274__B2 _21266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22379_ _22143_/X _22375_/X _15197_/B _22344_/A VGND VGND VPWR VPWR _22379_/X sky130_fd_sc_hd__o22a_4
X_12132_ _12168_/A _12132_/B VGND VGND VPWR VPWR _12133_/C sky130_fd_sc_hd__or2_4
X_24118_ _24203_/CLK _24118_/D HRESETn VGND VGND VPWR VPWR _24118_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15158__B _23585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21026__B2 _21020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12063_ _11943_/A VGND VGND VPWR VPWR _12093_/A sky130_fd_sc_hd__buf_2
X_16940_ _17644_/A VGND VGND VPWR VPWR _17645_/A sky130_fd_sc_hd__inv_2
X_24049_ _23155_/CLK _24049_/D VGND VGND VPWR VPWR _24049_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21577__A2 _21568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14997__B _23743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21176__A _21183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16871_ _16824_/D _13593_/B _16824_/D _13593_/B VGND VGND VPWR VPWR _16872_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23617__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18610_ _18610_/A _17735_/A _18609_/Y VGND VGND VPWR VPWR _18610_/X sky130_fd_sc_hd__or3_4
XANTENNA__15174__A _14737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15822_ _12895_/A _23821_/Q VGND VGND VPWR VPWR _15823_/C sky130_fd_sc_hd__or2_4
X_19590_ _19839_/A VGND VGND VPWR VPWR _19612_/A sky130_fd_sc_hd__buf_2
XANTENNA__21329__A2 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15753_ _11741_/X _15753_/B _15752_/X VGND VGND VPWR VPWR _15753_/X sky130_fd_sc_hd__or3_4
X_18541_ _17422_/B _18539_/X VGND VGND VPWR VPWR _18541_/X sky130_fd_sc_hd__or2_4
X_12965_ _12965_/A _12965_/B VGND VGND VPWR VPWR _12965_/X sky130_fd_sc_hd__or2_4
XFILLER_98_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18485__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17402__B1 _11886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11916_ _15986_/A VGND VGND VPWR VPWR _11916_/X sky130_fd_sc_hd__buf_2
X_14704_ _14666_/X _14632_/B VGND VGND VPWR VPWR _14704_/X sky130_fd_sc_hd__or2_4
XFILLER_59_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15684_ _12720_/A _15684_/B _15684_/C VGND VGND VPWR VPWR _15688_/B sky130_fd_sc_hd__and3_4
X_18472_ _17261_/X _18400_/X _17261_/X _18395_/C VGND VGND VPWR VPWR _18473_/B sky130_fd_sc_hd__a2bb2o_4
X_12896_ _12464_/A _12894_/X _12895_/X VGND VGND VPWR VPWR _12896_/X sky130_fd_sc_hd__and3_4
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14635_ _15037_/A _14635_/B VGND VGND VPWR VPWR _14636_/C sky130_fd_sc_hd__or2_4
X_17423_ _17382_/X _17423_/B VGND VGND VPWR VPWR _17423_/Y sky130_fd_sc_hd__nor2_4
X_11847_ _11847_/A VGND VGND VPWR VPWR _13682_/A sky130_fd_sc_hd__buf_2
XANTENNA__15621__B _23115_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14518__A _13695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13422__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14566_ _14492_/X _14565_/Y VGND VGND VPWR VPWR _14566_/X sky130_fd_sc_hd__or2_4
X_17354_ _17363_/A _17354_/B VGND VGND VPWR VPWR _17354_/X sky130_fd_sc_hd__or2_4
XFILLER_57_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11778_ _11754_/X VGND VGND VPWR VPWR _11821_/A sky130_fd_sc_hd__buf_2
XFILLER_105_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13517_ _13507_/X _13510_/X _13517_/C VGND VGND VPWR VPWR _13518_/C sky130_fd_sc_hd__or3_4
X_16305_ _16188_/A _23513_/Q VGND VGND VPWR VPWR _16306_/C sky130_fd_sc_hd__or2_4
X_17285_ _17285_/A _17342_/A VGND VGND VPWR VPWR _17286_/A sky130_fd_sc_hd__and2_4
X_14497_ _14533_/A _14497_/B VGND VGND VPWR VPWR _14497_/X sky130_fd_sc_hd__or2_4
XANTENNA__12038__A _11875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16236_ _16155_/X _16234_/Y VGND VGND VPWR VPWR _16236_/X sky130_fd_sc_hd__or2_4
X_19024_ _18994_/A VGND VGND VPWR VPWR _19024_/X sky130_fd_sc_hd__buf_2
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13448_ _12872_/A VGND VGND VPWR VPWR _13448_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20255__A _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16167_ _16162_/X _16164_/X _16167_/C VGND VGND VPWR VPWR _16168_/C sky130_fd_sc_hd__and3_4
XFILLER_115_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13379_ _13378_/X _13312_/B VGND VGND VPWR VPWR _13380_/C sky130_fd_sc_hd__or2_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15118_ _14073_/A _15086_/X _15118_/C VGND VGND VPWR VPWR _15118_/X sky130_fd_sc_hd__and3_4
X_16098_ _15986_/A _16098_/B _16098_/C VGND VGND VPWR VPWR _16098_/X sky130_fd_sc_hd__and3_4
X_15049_ _11839_/X _11615_/X _15018_/X _11592_/X _15048_/X VGND VGND VPWR VPWR _15050_/A
+ sky130_fd_sc_hd__a32o_4
X_19926_ _12101_/X _19926_/B VGND VGND VPWR VPWR _19926_/X sky130_fd_sc_hd__or2_4
XANTENNA__17564__A _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21017__B2 _21013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22214__B1 _16282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21086__A _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19857_ _19670_/X _19442_/B _19857_/C _19672_/C VGND VGND VPWR VPWR _19857_/X sky130_fd_sc_hd__and4_4
XFILLER_96_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15084__A _15108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18808_ _15249_/X _18802_/X _11541_/A _18803_/X VGND VGND VPWR VPWR _24417_/D sky130_fd_sc_hd__o22a_4
XFILLER_95_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19788_ _19866_/B _19786_/Y _19787_/Y VGND VGND VPWR VPWR _19788_/X sky130_fd_sc_hd__a21o_4
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18739_ _18203_/A _18160_/A _17613_/Y _18736_/X VGND VGND VPWR VPWR _18751_/B sky130_fd_sc_hd__a211o_4
XFILLER_37_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24387__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15812__A _15812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21750_ _21522_/X _21748_/X _23639_/Q _21745_/X VGND VGND VPWR VPWR _23639_/D sky130_fd_sc_hd__o22a_4
XFILLER_110_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20701_ _20641_/X _20699_/X _20701_/C VGND VGND VPWR VPWR _20701_/X sky130_fd_sc_hd__and3_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21681_ _21576_/X _21676_/X _14912_/B _21637_/X VGND VGND VPWR VPWR _23680_/D sky130_fd_sc_hd__o22a_4
XFILLER_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23420_ _23100_/CLK _23420_/D VGND VGND VPWR VPWR _16658_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20632_ _24238_/Q VGND VGND VPWR VPWR _20632_/Y sky130_fd_sc_hd__inv_2
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23351_ _23473_/CLK _22267_/X VGND VGND VPWR VPWR _16092_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20563_ _20468_/X _20561_/Y _24273_/Q _20562_/X VGND VGND VPWR VPWR _20563_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16643__A _16640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22302_ _16550_/B VGND VGND VPWR VPWR _22302_/X sky130_fd_sc_hd__buf_2
X_23282_ _23314_/CLK _22356_/X VGND VGND VPWR VPWR _23282_/Q sky130_fd_sc_hd__dfxtp_4
X_20494_ _20494_/A VGND VGND VPWR VPWR _20494_/X sky130_fd_sc_hd__buf_2
XFILLER_30_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17886__A1_N _11629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22233_ _22219_/A VGND VGND VPWR VPWR _22233_/X sky130_fd_sc_hd__buf_2
XANTENNA__15259__A _14315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18121__A1 _18107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14163__A _14146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18121__B2 _17531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22164_ _22086_/X _22158_/X _16283_/B _22162_/X VGND VGND VPWR VPWR _23417_/D sky130_fd_sc_hd__o22a_4
XFILLER_65_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21115_ _21130_/A VGND VGND VPWR VPWR _21115_/X sky130_fd_sc_hd__buf_2
X_22095_ _20486_/A VGND VGND VPWR VPWR _22095_/X sky130_fd_sc_hd__buf_2
XANTENNA__21559__A2 _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21046_ _20797_/X _21044_/X _13745_/B _21041_/X VGND VGND VPWR VPWR _24040_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17632__B1 _18107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13507__A _12964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22508__B2 _22504_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22997_ _22967_/A VGND VGND VPWR VPWR _22997_/X sky130_fd_sc_hd__buf_2
X_12750_ _12716_/X _12724_/X _12732_/X _12741_/X _12749_/X VGND VGND VPWR VPWR _12750_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15722__A _13130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21948_ _21833_/X _21945_/X _15410_/B _21942_/X VGND VGND VPWR VPWR _21948_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21192__B1 _15815_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21731__A2 _21726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11700_/X VGND VGND VPWR VPWR _11702_/A sky130_fd_sc_hd__buf_2
XFILLER_42_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _11618_/A VGND VGND VPWR VPWR _12681_/X sky130_fd_sc_hd__buf_2
XANTENNA__21162__C _21162_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21879_ _21802_/X _21873_/X _23577_/Q _21877_/X VGND VGND VPWR VPWR _23577_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14338__A _13686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _15604_/A _14416_/X _14420_/C VGND VGND VPWR VPWR _14421_/C sky130_fd_sc_hd__or3_4
XANTENNA__13242__A _13242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _17054_/A _17052_/A VGND VGND VPWR VPWR _11632_/X sky130_fd_sc_hd__and2_4
X_23618_ _23363_/CLK _23618_/D VGND VGND VPWR VPWR _15300_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_93_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _15589_/A _14344_/X _14351_/C VGND VGND VPWR VPWR _14351_/X sky130_fd_sc_hd__or3_4
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ _24434_/Q IRQ[19] _20156_/A VGND VGND VPWR VPWR _20098_/B sky130_fd_sc_hd__a21o_4
X_23549_ _23485_/CLK _21925_/X VGND VGND VPWR VPWR _23549_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21495__B2 _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13281_/X _13300_/X _13302_/C VGND VGND VPWR VPWR _13302_/X sky130_fd_sc_hd__and3_4
XFILLER_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17070_ _17069_/X VGND VGND VPWR VPWR _17070_/Y sky130_fd_sc_hd__inv_2
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _14322_/A VGND VGND VPWR VPWR _15534_/A sky130_fd_sc_hd__buf_2
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20075__A NMI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16272__B _16272_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16021_ _16048_/A _16021_/B _16020_/X VGND VGND VPWR VPWR _16028_/B sky130_fd_sc_hd__and3_4
XFILLER_100_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13233_ _13257_/A _23537_/Q VGND VGND VPWR VPWR _13233_/X sky130_fd_sc_hd__or2_4
XANTENNA__15169__A _14113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14073__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21798__A2 _21793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13164_ _12709_/A _13162_/X _13164_/C VGND VGND VPWR VPWR _13164_/X sky130_fd_sc_hd__and3_4
XANTENNA__22290__A _22269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12115_ _11844_/X _11620_/X _12082_/X _11599_/X _12114_/X VGND VGND VPWR VPWR _12115_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_65_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13095_ _13080_/A _23986_/Q VGND VGND VPWR VPWR _13095_/X sky130_fd_sc_hd__or2_4
X_17972_ _17818_/X _17819_/X _17813_/X _17805_/X VGND VGND VPWR VPWR _17973_/A sky130_fd_sc_hd__o22a_4
XFILLER_65_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14801__A _11669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19711_ HRDATA[21] VGND VGND VPWR VPWR _20490_/B sky130_fd_sc_hd__buf_2
X_12046_ _12083_/A _12123_/B VGND VGND VPWR VPWR _12049_/B sky130_fd_sc_hd__or2_4
X_16923_ _16923_/A _17105_/A VGND VGND VPWR VPWR _16923_/X sky130_fd_sc_hd__and2_4
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19642_ _19744_/B VGND VGND VPWR VPWR _19643_/A sky130_fd_sc_hd__buf_2
X_16854_ _16840_/C _16840_/B _13922_/A VGND VGND VPWR VPWR _16854_/X sky130_fd_sc_hd__o21a_4
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12321__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15805_ _12850_/A _15805_/B VGND VGND VPWR VPWR _15807_/B sky130_fd_sc_hd__or2_4
X_19573_ _19573_/A VGND VGND VPWR VPWR _19573_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13136__B _13135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13997_ _14050_/A _13995_/X _13997_/C VGND VGND VPWR VPWR _13997_/X sky130_fd_sc_hd__and3_4
X_16785_ _16768_/X _24059_/Q VGND VGND VPWR VPWR _16786_/C sky130_fd_sc_hd__or2_4
XFILLER_81_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19376__B1 _19374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18524_ _18714_/A _17416_/A _18442_/A VGND VGND VPWR VPWR _18524_/X sky130_fd_sc_hd__a21o_4
X_12948_ _12948_/A _12948_/B _12948_/C VGND VGND VPWR VPWR _12948_/X sky130_fd_sc_hd__or3_4
X_15736_ _13088_/A VGND VGND VPWR VPWR _15750_/A sky130_fd_sc_hd__buf_2
XFILLER_34_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21722__A2 _21719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18455_ _17701_/X _17751_/X _17701_/X _17751_/X VGND VGND VPWR VPWR _18455_/X sky130_fd_sc_hd__a2bb2o_4
X_12879_ _12879_/A _23923_/Q VGND VGND VPWR VPWR _12879_/X sky130_fd_sc_hd__or2_4
X_15667_ _15667_/A _15667_/B VGND VGND VPWR VPWR _15667_/X sky130_fd_sc_hd__or2_4
XFILLER_60_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13152__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17406_ _17171_/X _17407_/B VGND VGND VPWR VPWR _17409_/A sky130_fd_sc_hd__and2_4
X_14618_ _12439_/A _14698_/B VGND VGND VPWR VPWR _14618_/X sky130_fd_sc_hd__or2_4
X_15598_ _15598_/A _23915_/Q VGND VGND VPWR VPWR _15600_/B sky130_fd_sc_hd__or2_4
X_18386_ _18204_/A _17372_/X VGND VGND VPWR VPWR _18386_/X sky130_fd_sc_hd__or2_4
XANTENNA__21486__A1 _21273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14549_ _14494_/X _14547_/X _14549_/C VGND VGND VPWR VPWR _14549_/X sky130_fd_sc_hd__and3_4
X_17337_ _17337_/A VGND VGND VPWR VPWR _17337_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21486__B2 _21481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12991__A _12990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17268_ _17266_/X _17781_/B VGND VGND VPWR VPWR _17785_/B sky130_fd_sc_hd__or2_4
XANTENNA__16901__A2 _16900_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19007_ _24337_/Q VGND VGND VPWR VPWR _19007_/Y sky130_fd_sc_hd__inv_2
X_16219_ _16219_/A _16219_/B VGND VGND VPWR VPWR _16221_/B sky130_fd_sc_hd__or2_4
XFILLER_31_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21238__B2 _21230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17199_ _17227_/A _17185_/Y _17251_/A _17198_/Y VGND VGND VPWR VPWR _17199_/X sky130_fd_sc_hd__o22a_4
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21809__A _20464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17294__A _14565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15807__A _11912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19909_ _19909_/A VGND VGND VPWR VPWR _19909_/X sky130_fd_sc_hd__buf_2
XFILLER_29_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15526__B _23723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22920_ _22899_/X _16960_/A VGND VGND VPWR VPWR _22920_/X sky130_fd_sc_hd__or2_4
XFILLER_99_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21410__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12231__A _12198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21961__A2 _21959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21544__A _21532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22851_ _12338_/Y _22824_/X _22777_/X _22850_/X VGND VGND VPWR VPWR _22852_/A sky130_fd_sc_hd__a211o_4
XFILLER_72_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21802_ _21802_/A VGND VGND VPWR VPWR _21802_/X sky130_fd_sc_hd__buf_2
XFILLER_37_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15542__A _12533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22782_ _22781_/X VGND VGND VPWR VPWR _22782_/X sky130_fd_sc_hd__buf_2
XFILLER_52_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21713__A2 _21712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22910__A1 _18640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21733_ _23646_/Q VGND VGND VPWR VPWR _21733_/Y sky130_fd_sc_hd__inv_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14158__A _14158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23312__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13062__A _13726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24452_ _24203_/CLK _24452_/D HRESETn VGND VGND VPWR VPWR _20093_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21664_ _21546_/X _21662_/X _15838_/B _21659_/X VGND VGND VPWR VPWR _21664_/X sky130_fd_sc_hd__o22a_4
XFILLER_75_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22375__A _22368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23403_ _23688_/CLK _23403_/D VGND VGND VPWR VPWR _23403_/Q sky130_fd_sc_hd__dfxtp_4
X_20615_ _20399_/A VGND VGND VPWR VPWR _20634_/A sky130_fd_sc_hd__buf_2
XANTENNA__17469__A _17662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13997__A _14050_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24383_ _24425_/CLK _24383_/D HRESETn VGND VGND VPWR VPWR _24383_/Q sky130_fd_sc_hd__dfrtp_4
X_21595_ _21595_/A VGND VGND VPWR VPWR _21595_/X sky130_fd_sc_hd__buf_2
XANTENNA__16373__A _11658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23334_ _23270_/CLK _22291_/X VGND VGND VPWR VPWR _14271_/B sky130_fd_sc_hd__dfxtp_4
X_20546_ _20502_/A _20546_/B VGND VGND VPWR VPWR _20546_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16092__B _16092_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23265_ _24032_/CLK _22379_/X VGND VGND VPWR VPWR _15197_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20477_ _20293_/X _20476_/X _18982_/A _20303_/X VGND VGND VPWR VPWR _20477_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12406__A _15889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22216_ _22088_/X _22215_/X _15984_/B _22212_/X VGND VGND VPWR VPWR _23384_/D sky130_fd_sc_hd__o22a_4
XFILLER_69_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21719__A _21690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23196_ _23324_/CLK _22524_/X VGND VGND VPWR VPWR _16614_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20988__B1 _19770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12125__B _23741_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22147_ _21001_/A VGND VGND VPWR VPWR _22147_/X sky130_fd_sc_hd__buf_2
XANTENNA__15717__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20342__B _20342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22078_ _22075_/X _22077_/X _12140_/B _22072_/X VGND VGND VPWR VPWR _23453_/D sky130_fd_sc_hd__o22a_4
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13237__A _11664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13920_ _13921_/B VGND VGND VPWR VPWR _13920_/X sky130_fd_sc_hd__buf_2
X_21029_ _20509_/X _21023_/X _24052_/Q _21027_/X VGND VGND VPWR VPWR _24052_/D sky130_fd_sc_hd__o22a_4
XFILLER_101_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_12_0_HCLK_A clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13851_ _13851_/A VGND VGND VPWR VPWR _13895_/A sky130_fd_sc_hd__buf_2
XFILLER_25_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16548__A _16569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12802_ _12802_/A _23316_/Q VGND VGND VPWR VPWR _12804_/B sky130_fd_sc_hd__or2_4
XANTENNA__11980__A _11980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13782_ _12450_/A _13782_/B _13781_/X VGND VGND VPWR VPWR _13782_/X sky130_fd_sc_hd__and3_4
X_16570_ _16542_/A _16570_/B _16570_/C VGND VGND VPWR VPWR _16570_/X sky130_fd_sc_hd__or3_4
XANTENNA__21704__A2 _21698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24334__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16267__B _16267_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12733_ _12713_/A VGND VGND VPWR VPWR _15820_/A sky130_fd_sc_hd__buf_2
X_15521_ _15518_/X _15520_/Y VGND VGND VPWR VPWR _15914_/A sky130_fd_sc_hd__or2_4
XANTENNA__20912__B1 _20911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15452_ _13594_/X _13595_/X _15421_/X _11595_/A _15451_/X VGND VGND VPWR VPWR _15453_/A
+ sky130_fd_sc_hd__a32o_4
X_18240_ _18240_/A VGND VGND VPWR VPWR _18244_/A sky130_fd_sc_hd__buf_2
XFILLER_71_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12664_ _12976_/A _12542_/B VGND VGND VPWR VPWR _12664_/X sky130_fd_sc_hd__or2_4
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _15626_/A _14401_/X _14402_/X VGND VGND VPWR VPWR _14404_/C sky130_fd_sc_hd__and3_4
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11614_/X VGND VGND VPWR VPWR _11615_/X sky130_fd_sc_hd__buf_2
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_53_0_HCLK clkbuf_6_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15383_ _15312_/X _15380_/Y _15185_/X _15251_/A VGND VGND VPWR VPWR _15384_/A sky130_fd_sc_hd__o22a_4
X_18171_ _18171_/A VGND VGND VPWR VPWR _18171_/X sky130_fd_sc_hd__buf_2
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17379__A _15909_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21468__B2 _21467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12595_ _12640_/A _12463_/B VGND VGND VPWR VPWR _12596_/C sky130_fd_sc_hd__or2_4
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ _13682_/A _14333_/X VGND VGND VPWR VPWR _14334_/X sky130_fd_sc_hd__and2_4
X_17122_ _11912_/A _17105_/X _21007_/A _17033_/A VGND VGND VPWR VPWR _17122_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13700__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _24436_/Q IRQ[21] _20158_/A VGND VGND VPWR VPWR _11547_/B sky130_fd_sc_hd__a21o_4
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17053_ _17052_/X VGND VGND VPWR VPWR _17068_/A sky130_fd_sc_hd__buf_2
X_14265_ _14265_/A VGND VGND VPWR VPWR _14265_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12316__A _15693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16004_ _15929_/X _16004_/B _16003_/X VGND VGND VPWR VPWR _16004_/X sky130_fd_sc_hd__or3_4
XFILLER_13_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13216_ _13239_/A _13149_/B VGND VGND VPWR VPWR _13216_/X sky130_fd_sc_hd__or2_4
X_14196_ _14207_/A VGND VGND VPWR VPWR _14215_/A sky130_fd_sc_hd__buf_2
XFILLER_97_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13147_ _12744_/A VGND VGND VPWR VPWR _15687_/A sky130_fd_sc_hd__buf_2
XANTENNA__15627__A _15611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21348__B _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14531__A _11664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13078_ _13119_/A _24018_/Q VGND VGND VPWR VPWR _13078_/X sky130_fd_sc_hd__or2_4
X_17955_ _18205_/A _17570_/Y VGND VGND VPWR VPWR _17959_/B sky130_fd_sc_hd__and2_4
XANTENNA__22196__A2 _22193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12029_ _11844_/X _11619_/X _11991_/X _11598_/X _12028_/X VGND VGND VPWR VPWR _12029_/X
+ sky130_fd_sc_hd__a32o_4
X_16906_ _16905_/X VGND VGND VPWR VPWR _16906_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13147__A _12744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17886_ _11629_/X _17885_/X _24476_/Q _11629_/X VGND VGND VPWR VPWR _24476_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21943__A2 _21938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19625_ _19866_/B VGND VGND VPWR VPWR _19625_/Y sky130_fd_sc_hd__inv_2
X_16837_ _15914_/A _16836_/X _15914_/A _16836_/X VGND VGND VPWR VPWR _16837_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12986__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16458__A _12837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23335__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15362__A _14020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19556_ _19877_/B VGND VGND VPWR VPWR _19556_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16768_ _12153_/A VGND VGND VPWR VPWR _16768_/X sky130_fd_sc_hd__buf_2
XFILLER_34_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16177__B _16103_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18507_ _18458_/X _18484_/Y _18485_/X _18506_/X VGND VGND VPWR VPWR _18507_/X sky130_fd_sc_hd__o22a_4
XFILLER_62_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15719_ _12765_/X _15719_/B _15719_/C VGND VGND VPWR VPWR _15719_/X sky130_fd_sc_hd__and3_4
XANTENNA__19769__A HRDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19487_ _19483_/X _19481_/A _19486_/Y VGND VGND VPWR VPWR _19499_/A sky130_fd_sc_hd__o21a_4
X_16699_ _12088_/A _16697_/X _16699_/C VGND VGND VPWR VPWR _16703_/B sky130_fd_sc_hd__and3_4
XANTENNA__18673__A _18392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18438_ _18011_/X _18352_/B _18436_/Y _18016_/X _18437_/Y VGND VGND VPWR VPWR _18438_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_72_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23485__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21459__A1 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21459__B2 _21453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18369_ _17796_/X _18368_/X _17868_/X VGND VGND VPWR VPWR _18392_/B sky130_fd_sc_hd__o21a_4
XANTENNA__19521__B1 HRDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20400_ _20342_/A _20400_/B VGND VGND VPWR VPWR _20400_/X sky130_fd_sc_hd__and2_4
X_21380_ _21373_/A VGND VGND VPWR VPWR _21380_/X sky130_fd_sc_hd__buf_2
XFILLER_30_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20131__A1 _19884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22923__A _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20331_ _20321_/X _20329_/X _19137_/A _20330_/X VGND VGND VPWR VPWR _20331_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16921__A _16919_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12226__A _12556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23050_ _23050_/A VGND VGND VPWR VPWR HADDR[29] sky130_fd_sc_hd__inv_2
XANTENNA__19852__A1_N _19730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20262_ _20255_/X _20261_/X _24382_/Q _18872_/B VGND VGND VPWR VPWR _20262_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21539__A _21527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22001_ _21838_/X _21995_/X _23498_/Q _21999_/X VGND VGND VPWR VPWR _23498_/D sky130_fd_sc_hd__o22a_4
XFILLER_116_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15537__A _15556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20193_ _20193_/A VGND VGND VPWR VPWR _20196_/B sky130_fd_sc_hd__inv_2
XFILLER_118_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21631__B2 _21595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15256__B _15256_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24110__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22187__A2 _22186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23952_ _23983_/CLK _21188_/X VGND VGND VPWR VPWR _23952_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21395__B1 _23840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22903_ _18664_/X _22889_/X VGND VGND VPWR VPWR _22904_/C sky130_fd_sc_hd__or2_4
X_23883_ _23915_/CLK _21331_/X VGND VGND VPWR VPWR _23883_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12896__A _12464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16368__A _11715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15272__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22834_ _22834_/A VGND VGND VPWR VPWR HWDATA[17] sky130_fd_sc_hd__inv_2
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22765_ _22763_/Y _22765_/B _22754_/X VGND VGND VPWR VPWR _24100_/D sky130_fd_sc_hd__and3_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18583__A _17792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19760__B1 _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21716_ _21702_/A VGND VGND VPWR VPWR _21716_/X sky130_fd_sc_hd__buf_2
XFILLER_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22696_ _21263_/A _22693_/X _23084_/Q _22690_/X VGND VGND VPWR VPWR _22696_/X sky130_fd_sc_hd__o22a_4
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24435_ _24435_/CLK _18784_/X HRESETn VGND VGND VPWR VPWR _20520_/A sky130_fd_sc_hd__dfrtp_4
X_21647_ _21517_/X _21641_/X _16296_/B _21645_/X VGND VGND VPWR VPWR _21647_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22111__A2 _22101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12380_ _12360_/A _12246_/B VGND VGND VPWR VPWR _12382_/B sky130_fd_sc_hd__or2_4
X_24366_ _24334_/CLK _24366_/D HRESETn VGND VGND VPWR VPWR _24366_/Q sky130_fd_sc_hd__dfstp_4
X_21578_ _21293_/A VGND VGND VPWR VPWR _21578_/X sky130_fd_sc_hd__buf_2
X_23317_ _24021_/CLK _23317_/D VGND VGND VPWR VPWR _23317_/Q sky130_fd_sc_hd__dfxtp_4
X_20529_ _20603_/A _20529_/B VGND VGND VPWR VPWR _20529_/Y sky130_fd_sc_hd__nor2_4
XFILLER_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24297_ _24299_/CLK _19182_/X HRESETn VGND VGND VPWR VPWR _24297_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14050_ _14050_/A _14048_/X _14050_/C VGND VGND VPWR VPWR _14050_/X sky130_fd_sc_hd__and3_4
X_23248_ _23920_/CLK _22424_/X VGND VGND VPWR VPWR _13282_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23208__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17646__B _17646_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19815__B2 _19730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13001_ _12879_/A _13069_/B VGND VGND VPWR VPWR _13003_/B sky130_fd_sc_hd__or2_4
X_23179_ _23336_/CLK _23179_/D VGND VGND VPWR VPWR _23179_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21622__B2 _21616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12115__A1 _11844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22178__A2 _22172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17740_ _16997_/A _17122_/X _17738_/X _17739_/X VGND VGND VPWR VPWR _17740_/X sky130_fd_sc_hd__o22a_4
X_14952_ _14642_/A _14952_/B _14952_/C VGND VGND VPWR VPWR _14953_/C sky130_fd_sc_hd__or3_4
XFILLER_62_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21925__A2 _21924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13903_ _13879_/A _13829_/B VGND VGND VPWR VPWR _13903_/X sky130_fd_sc_hd__or2_4
X_17671_ _16948_/Y VGND VGND VPWR VPWR _17672_/A sky130_fd_sc_hd__buf_2
X_14883_ _14880_/A _14883_/B VGND VGND VPWR VPWR _14883_/X sky130_fd_sc_hd__or2_4
XANTENNA__16278__A _15980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19410_ _19406_/X _18702_/X _19406_/X _24193_/Q VGND VGND VPWR VPWR _24193_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15182__A _15032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16622_ _16622_/A _16616_/X _16622_/C VGND VGND VPWR VPWR _16623_/C sky130_fd_sc_hd__or3_4
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13834_ _15449_/A _13830_/X _13833_/X VGND VGND VPWR VPWR _13834_/X sky130_fd_sc_hd__or3_4
XFILLER_75_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19341_ _19340_/X _18477_/X _19340_/X _24235_/Q VGND VGND VPWR VPWR _24235_/D sky130_fd_sc_hd__a2bb2o_4
X_13765_ _13765_/A _13765_/B _13765_/C VGND VGND VPWR VPWR _13769_/B sky130_fd_sc_hd__and3_4
X_16553_ _16715_/A _16550_/X _16553_/C VGND VGND VPWR VPWR _16553_/X sky130_fd_sc_hd__and3_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21689__B2 _21688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22350__A2 _22347_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15504_ _15480_/A _15504_/B VGND VGND VPWR VPWR _15504_/X sky130_fd_sc_hd__or2_4
XANTENNA__15910__A _15844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12716_ _13026_/A VGND VGND VPWR VPWR _12716_/X sky130_fd_sc_hd__buf_2
X_19272_ _19217_/A _19217_/B _19271_/Y VGND VGND VPWR VPWR _24268_/D sky130_fd_sc_hd__o21a_4
X_13696_ _13695_/X _13696_/B VGND VGND VPWR VPWR _13696_/X sky130_fd_sc_hd__or2_4
X_16484_ _16506_/A _16482_/X _16484_/C VGND VGND VPWR VPWR _16484_/X sky130_fd_sc_hd__and3_4
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18223_ _18171_/X _19382_/A _18202_/X _18222_/X VGND VGND VPWR VPWR _18223_/X sky130_fd_sc_hd__o22a_4
XFILLER_62_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12647_ _12591_/X _12647_/B VGND VGND VPWR VPWR _12647_/X sky130_fd_sc_hd__or2_4
X_15435_ _15435_/A _15435_/B _15435_/C VGND VGND VPWR VPWR _15435_/X sky130_fd_sc_hd__or3_4
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14526__A _13695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22102__A2 _22101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15366_ _14000_/A _15306_/B VGND VGND VPWR VPWR _15368_/B sky130_fd_sc_hd__or2_4
X_18154_ _18153_/Y _17514_/B _17521_/X VGND VGND VPWR VPWR _18154_/X sky130_fd_sc_hd__o21a_4
X_12578_ _12578_/A VGND VGND VPWR VPWR _12935_/A sky130_fd_sc_hd__buf_2
XFILLER_89_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22743__A SYSTICKCLKDIV[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17105_ _17105_/A _17105_/B VGND VGND VPWR VPWR _17105_/X sky130_fd_sc_hd__and2_4
X_11529_ _24344_/Q _11528_/X VGND VGND VPWR VPWR _18959_/A sky130_fd_sc_hd__or2_4
X_14317_ _14431_/A _14317_/B VGND VGND VPWR VPWR _14317_/X sky130_fd_sc_hd__or2_4
X_15297_ _14756_/A _15297_/B VGND VGND VPWR VPWR _15297_/X sky130_fd_sc_hd__or2_4
X_18085_ _18085_/A _18085_/B VGND VGND VPWR VPWR _18085_/X sky130_fd_sc_hd__or2_4
XANTENNA__16741__A _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14248_ _14218_/X _23849_/Q VGND VGND VPWR VPWR _14249_/C sky130_fd_sc_hd__or2_4
X_17036_ _17036_/A _17342_/A VGND VGND VPWR VPWR _17105_/B sky130_fd_sc_hd__or2_4
XANTENNA__21359__A _21359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16460__B _16391_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11885__A _11884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14179_ _14197_/A VGND VGND VPWR VPWR _14225_/A sky130_fd_sc_hd__buf_2
XANTENNA__21613__B2 _21609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14261__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18987_ _18987_/A VGND VGND VPWR VPWR _19002_/A sky130_fd_sc_hd__buf_2
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17572__A _17165_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17938_ _17794_/A _17937_/X VGND VGND VPWR VPWR _17938_/Y sky130_fd_sc_hd__nor2_4
XFILLER_97_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17045__A1 _12116_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17045__B2 _17044_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17869_ _17868_/X VGND VGND VPWR VPWR _17869_/X sky130_fd_sc_hd__buf_2
XFILLER_38_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16188__A _16188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18793__A1 _17191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19608_ _19481_/B _19600_/B VGND VGND VPWR VPWR _19862_/A sky130_fd_sc_hd__and2_4
XANTENNA__13605__A _13959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20880_ _20877_/X _20879_/X _20240_/X VGND VGND VPWR VPWR _20880_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21129__B1 _12248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19539_ _19428_/A _19872_/B VGND VGND VPWR VPWR _19637_/A sky130_fd_sc_hd__or2_4
XFILLER_39_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15820__A _15820_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22550_ _22521_/A VGND VGND VPWR VPWR _22550_/X sky130_fd_sc_hd__buf_2
XANTENNA__24380__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21501_ _21556_/A VGND VGND VPWR VPWR _21527_/A sky130_fd_sc_hd__inv_2
X_22481_ _22406_/X _22479_/X _16226_/B _22476_/X VGND VGND VPWR VPWR _22481_/X sky130_fd_sc_hd__o22a_4
XFILLER_72_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14436__A _14463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24220_ _24187_/CLK _19368_/X HRESETn VGND VGND VPWR VPWR _24220_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13340__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21432_ _21268_/X _21426_/X _23818_/Q _21430_/X VGND VGND VPWR VPWR _21432_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16859__A1 _15051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24151_ _24223_/CLK _19912_/X HRESETn VGND VGND VPWR VPWR _24151_/Q sky130_fd_sc_hd__dfrtp_4
X_21363_ _21234_/X _21362_/X _23864_/Q _21359_/X VGND VGND VPWR VPWR _23864_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19665__C _19672_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23102_ _23774_/CLK _22670_/X VGND VGND VPWR VPWR _23102_/Q sky130_fd_sc_hd__dfxtp_4
X_20314_ _20314_/A VGND VGND VPWR VPWR _21791_/A sky130_fd_sc_hd__buf_2
X_24082_ _24082_/CLK _20554_/X VGND VGND VPWR VPWR _24082_/Q sky130_fd_sc_hd__dfxtp_4
X_21294_ _21293_/X _21247_/A _23903_/Q _21230_/A VGND VGND VPWR VPWR _21294_/X sky130_fd_sc_hd__o22a_4
XFILLER_11_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23033_ _18050_/X _23017_/B VGND VGND VPWR VPWR _23033_/X sky130_fd_sc_hd__or2_4
XANTENNA__15267__A _11894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11795__A _16045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20245_ _20248_/A _20073_/X VGND VGND VPWR VPWR _20525_/A sky130_fd_sc_hd__or2_4
XANTENNA__21604__B2 _21602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14171__A _15032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20176_ _20176_/A _20175_/X VGND VGND VPWR VPWR _20176_/X sky130_fd_sc_hd__or2_4
XANTENNA__19681__B HRDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21368__B1 _23860_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21907__A2 _21901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23935_ _23130_/CLK _23935_/D VGND VGND VPWR VPWR _15088_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15714__B _15652_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18784__A1 _12990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22580__A2 _22579_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11880_ _15543_/A VGND VGND VPWR VPWR _14283_/A sky130_fd_sc_hd__buf_2
X_23866_ _23706_/CLK _21360_/X VGND VGND VPWR VPWR _16438_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22817_ _22813_/X _22817_/B VGND VGND VPWR VPWR HWDATA[13] sky130_fd_sc_hd__nor2_4
XFILLER_60_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23797_ _23315_/CLK _21468_/X VGND VGND VPWR VPWR _12658_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13550_ _13550_/A _13547_/X _13549_/X VGND VGND VPWR VPWR _13550_/X sky130_fd_sc_hd__and3_4
XFILLER_41_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15730__A _15725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22748_ _22747_/X VGND VGND VPWR VPWR _22748_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18000__A3 _17987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12501_ _12500_/X _12633_/B VGND VGND VPWR VPWR _12501_/X sky130_fd_sc_hd__or2_4
XFILLER_40_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13481_ _13477_/X _13569_/B VGND VGND VPWR VPWR _13482_/C sky130_fd_sc_hd__or2_4
X_22679_ _22686_/A VGND VGND VPWR VPWR _22679_/X sky130_fd_sc_hd__buf_2
XFILLER_9_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15220_ _14195_/A _15220_/B _15219_/X VGND VGND VPWR VPWR _15220_/X sky130_fd_sc_hd__and3_4
XFILLER_16_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13250__A _12350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12432_ _12338_/Y _12429_/X VGND VGND VPWR VPWR _12432_/X sky130_fd_sc_hd__or2_4
X_24418_ _24425_/CLK _24418_/D HRESETn VGND VGND VPWR VPWR _24418_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24156__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15151_ _11608_/A _15149_/X _15151_/C VGND VGND VPWR VPWR _15151_/X sky130_fd_sc_hd__and3_4
X_12363_ _11741_/X _12363_/B _12362_/X VGND VGND VPWR VPWR _12364_/C sky130_fd_sc_hd__or3_4
X_24349_ _24344_/CLK _24349_/D HRESETn VGND VGND VPWR VPWR _11533_/D sky130_fd_sc_hd__dfstp_4
XFILLER_103_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16561__A _11936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14102_ _15010_/A VGND VGND VPWR VPWR _14992_/A sky130_fd_sc_hd__buf_2
X_15082_ _11710_/A _23519_/Q VGND VGND VPWR VPWR _15083_/C sky130_fd_sc_hd__or2_4
X_12294_ _12726_/A _12294_/B VGND VGND VPWR VPWR _12294_/X sky130_fd_sc_hd__or2_4
XFILLER_10_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12336__A1 _12892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16280__B _16280_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14033_ _12599_/A _14033_/B _14033_/C VGND VGND VPWR VPWR _14033_/X sky130_fd_sc_hd__and3_4
X_18910_ _13918_/X _18905_/X _19068_/A _18906_/X VGND VGND VPWR VPWR _24359_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15177__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19890_ _24158_/Q VGND VGND VPWR VPWR _20218_/A sky130_fd_sc_hd__inv_2
XANTENNA__14081__A _12196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17275__A1 _17272_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18841_ _18841_/A VGND VGND VPWR VPWR _18841_/X sky130_fd_sc_hd__buf_2
XANTENNA__17275__B2 _17274_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18472__B1 _17261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15905__A _13572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18772_ _17277_/X _18765_/X _24443_/Q _18768_/X VGND VGND VPWR VPWR _18772_/X sky130_fd_sc_hd__o22a_4
XFILLER_114_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15984_ _15984_/A _15984_/B VGND VGND VPWR VPWR _15986_/B sky130_fd_sc_hd__or2_4
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13836__A1 _12269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17723_ _17723_/A _17723_/B VGND VGND VPWR VPWR _17745_/A sky130_fd_sc_hd__or2_4
X_14935_ _14202_/A _14935_/B _14934_/X VGND VGND VPWR VPWR _14954_/B sky130_fd_sc_hd__and3_4
XANTENNA__15624__B _23371_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13425__A _11658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17654_ _17653_/X VGND VGND VPWR VPWR _17654_/Y sky130_fd_sc_hd__inv_2
X_14866_ _13983_/A _14866_/B VGND VGND VPWR VPWR _14869_/B sky130_fd_sc_hd__or2_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20582__A1 _20494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22738__A SYSTICKCLKDIV[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16605_ _16621_/A _16602_/X _16605_/C VGND VGND VPWR VPWR _16612_/B sky130_fd_sc_hd__and3_4
XFILLER_51_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13817_ _13794_/A _23367_/Q VGND VGND VPWR VPWR _13819_/B sky130_fd_sc_hd__or2_4
XANTENNA__22859__B1 _13685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17585_ _17471_/X _17584_/Y _17464_/B _17473_/X VGND VGND VPWR VPWR _17626_/B sky130_fd_sc_hd__a211o_4
XFILLER_17_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14797_ _13694_/A _14797_/B VGND VGND VPWR VPWR _14799_/B sky130_fd_sc_hd__or2_4
XFILLER_1_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16736__A _11875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19324_ _19321_/X _18168_/X _19321_/X _24246_/Q VGND VGND VPWR VPWR _19324_/X sky130_fd_sc_hd__a2bb2o_4
X_16536_ _16536_/A _23772_/Q VGND VGND VPWR VPWR _16537_/C sky130_fd_sc_hd__or2_4
X_13748_ _11648_/X _13660_/B VGND VGND VPWR VPWR _13750_/B sky130_fd_sc_hd__or2_4
XFILLER_56_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12983__B _12983_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16455__B _16387_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19255_ _19225_/X VGND VGND VPWR VPWR _19255_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16467_ _16158_/A _16407_/B VGND VGND VPWR VPWR _16467_/X sky130_fd_sc_hd__or2_4
X_13679_ _15447_/A _13760_/B VGND VGND VPWR VPWR _13680_/C sky130_fd_sc_hd__or2_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18206_ _18206_/A _17454_/A VGND VGND VPWR VPWR _18208_/C sky130_fd_sc_hd__and2_4
XANTENNA__13160__A _12737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15418_ _13654_/A _15418_/B _15418_/C VGND VGND VPWR VPWR _15419_/C sky130_fd_sc_hd__and3_4
X_19186_ _24295_/Q _19116_/B _19185_/Y VGND VGND VPWR VPWR _24295_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_5_23_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_23_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16398_ _16397_/X _16398_/B VGND VGND VPWR VPWR _16398_/X sky130_fd_sc_hd__or2_4
X_18137_ _18137_/A VGND VGND VPWR VPWR _18266_/A sky130_fd_sc_hd__buf_2
X_15349_ _15314_/A _15283_/B VGND VGND VPWR VPWR _15350_/C sky130_fd_sc_hd__or2_4
XFILLER_69_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21834__B2 _21824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20705__B _20595_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21089__A _21075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18068_ _18068_/A VGND VGND VPWR VPWR _18068_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17019_ _17018_/X VGND VGND VPWR VPWR _17020_/A sky130_fd_sc_hd__buf_2
XANTENNA__12504__A _12518_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20030_ _18379_/X _20009_/X _20029_/Y _20020_/X VGND VGND VPWR VPWR _20030_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21817__A _21817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18398__A _18713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11550__A2 IRQ[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15815__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22011__B2 _22006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21981_ _21988_/A VGND VGND VPWR VPWR _21981_/X sky130_fd_sc_hd__buf_2
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23720_ _23304_/CLK _21621_/X VGND VGND VPWR VPWR _13703_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13335__A _12849_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22562__A2 _22557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20932_ _20932_/A VGND VGND VPWR VPWR _20932_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23651_ _23270_/CLK _21728_/X VGND VGND VPWR VPWR _14739_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ _18624_/X _20653_/X _20758_/X _20862_/Y VGND VGND VPWR VPWR _20864_/A sky130_fd_sc_hd__a211o_4
XFILLER_74_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16646__A _16045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22602_ _22442_/X _22600_/X _13727_/B _22597_/X VGND VGND VPWR VPWR _23144_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15550__A _12269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23582_ _23320_/CLK _21871_/X VGND VGND VPWR VPWR _23582_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20794_ _20634_/A _20793_/X VGND VGND VPWR VPWR _20794_/Y sky130_fd_sc_hd__nand2_4
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22533_ _22533_/A VGND VGND VPWR VPWR _22533_/X sky130_fd_sc_hd__buf_2
XFILLER_10_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19957__A _19929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17741__A2 _17117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22464_ _12014_/B VGND VGND VPWR VPWR _22464_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22078__B2 _22072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24203_ _24203_/CLK _24203_/D HRESETn VGND VGND VPWR VPWR _24203_/Q sky130_fd_sc_hd__dfrtp_4
X_21415_ _21239_/X _21412_/X _12294_/B _21409_/X VGND VGND VPWR VPWR _21415_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21825__A1 _21823_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17477__A _13493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21825__B2 _21824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22395_ _22394_/X _22392_/X _16602_/B _22387_/X VGND VGND VPWR VPWR _22395_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16381__A _15997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24134_ _24239_/CLK _19989_/Y HRESETn VGND VGND VPWR VPWR _17652_/A sky130_fd_sc_hd__dfrtp_4
X_21346_ _21293_/X _21319_/A _23871_/Q _21301_/X VGND VGND VPWR VPWR _21346_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24065_ _24065_/CLK _20959_/X VGND VGND VPWR VPWR _15241_/B sky130_fd_sc_hd__dfxtp_4
X_21277_ _20838_/A VGND VGND VPWR VPWR _21277_/X sky130_fd_sc_hd__buf_2
X_23016_ _23003_/A _23016_/B VGND VGND VPWR VPWR _23018_/B sky130_fd_sc_hd__nand2_4
XFILLER_81_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20228_ _20286_/A VGND VGND VPWR VPWR _20229_/A sky130_fd_sc_hd__buf_2
XFILLER_85_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21053__A2 _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_43_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR _23368_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_77_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15725__A _15725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20159_ _24436_/Q IRQ[21] _20158_/X VGND VGND VPWR VPWR _20159_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_77_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12981_ _12981_/A _12909_/B VGND VGND VPWR VPWR _12981_/X sky130_fd_sc_hd__or2_4
XANTENNA__15444__B _23788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14491__A1 _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22553__A2 _22550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14720_ _14719_/X VGND VGND VPWR VPWR _14723_/B sky130_fd_sc_hd__inv_2
XFILLER_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11932_ _13048_/A VGND VGND VPWR VPWR _12914_/A sky130_fd_sc_hd__buf_2
X_23918_ _23922_/CLK _23918_/D VGND VGND VPWR VPWR _15729_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20564__A1 _20518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20564__B2 _20525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11863_ _16152_/A VGND VGND VPWR VPWR _16113_/A sky130_fd_sc_hd__buf_2
X_14651_ _15201_/A VGND VGND VPWR VPWR _14679_/A sky130_fd_sc_hd__buf_2
X_23849_ _23847_/CLK _23849_/D VGND VGND VPWR VPWR _23849_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16556__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13602_ _14778_/A VGND VGND VPWR VPWR _13603_/A sky130_fd_sc_hd__buf_2
XFILLER_57_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15460__A _12638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17370_ _15780_/B _18387_/B VGND VGND VPWR VPWR _17370_/X sky130_fd_sc_hd__and2_4
X_11794_ _11772_/X _11783_/X _11793_/X VGND VGND VPWR VPWR _11794_/X sky130_fd_sc_hd__and3_4
X_14582_ _15015_/A VGND VGND VPWR VPWR _15028_/A sky130_fd_sc_hd__buf_2
XFILLER_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16321_ _11673_/X _16313_/X _16320_/X VGND VGND VPWR VPWR _16321_/X sky130_fd_sc_hd__and3_4
X_13533_ _13561_/A _23311_/Q VGND VGND VPWR VPWR _13535_/B sky130_fd_sc_hd__or2_4
XANTENNA__17193__B1 _13278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19040_ _19030_/X _19039_/X _19030_/X _24332_/Q VGND VGND VPWR VPWR _24332_/D sky130_fd_sc_hd__a2bb2o_4
X_13464_ _11913_/X _13462_/X _13464_/C VGND VGND VPWR VPWR _13464_/X sky130_fd_sc_hd__and3_4
X_16252_ _11959_/X VGND VGND VPWR VPWR _16252_/X sky130_fd_sc_hd__buf_2
XANTENNA__22293__A _22286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12415_ _12386_/X _12332_/B VGND VGND VPWR VPWR _12416_/C sky130_fd_sc_hd__or2_4
X_15203_ _15203_/A _15201_/X _15203_/C VGND VGND VPWR VPWR _15207_/B sky130_fd_sc_hd__and3_4
XANTENNA__17387__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13395_ _12827_/A VGND VGND VPWR VPWR _13395_/X sky130_fd_sc_hd__buf_2
X_16183_ _16203_/A _16183_/B _16183_/C VGND VGND VPWR VPWR _16183_/X sky130_fd_sc_hd__and3_4
XANTENNA__24434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14804__A _12575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17496__A1 _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12346_ _12794_/A VGND VGND VPWR VPWR _12828_/A sky130_fd_sc_hd__buf_2
X_15134_ _12252_/A _15132_/X _15134_/C VGND VGND VPWR VPWR _15134_/X sky130_fd_sc_hd__and3_4
XANTENNA__21292__A2 _21283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15065_ _12583_/A _23263_/Q VGND VGND VPWR VPWR _15065_/X sky130_fd_sc_hd__or2_4
X_19942_ _18265_/A _18743_/X VGND VGND VPWR VPWR _19944_/C sky130_fd_sc_hd__nor2_4
X_12277_ _12198_/X _12274_/X _12276_/X VGND VGND VPWR VPWR _12277_/X sky130_fd_sc_hd__and3_4
XANTENNA__12324__A _12739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14016_ _14045_/A _13939_/B VGND VGND VPWR VPWR _14016_/X sky130_fd_sc_hd__or2_4
XANTENNA__21637__A _21659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19873_ _19580_/X _19873_/B _19839_/B _19872_/X VGND VGND VPWR VPWR _19873_/X sky130_fd_sc_hd__or4_4
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22241__B2 _22240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18824_ _17266_/X _18818_/X _24412_/Q _18821_/X VGND VGND VPWR VPWR _24412_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18011__A _18174_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18755_ _16927_/A _18753_/X _17639_/A _18754_/Y VGND VGND VPWR VPWR _18755_/X sky130_fd_sc_hd__o22a_4
XFILLER_83_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_0_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15967_ _15959_/A _15967_/B VGND VGND VPWR VPWR _15970_/B sky130_fd_sc_hd__or2_4
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22544__A2 _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18946__A _18999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17706_ _17704_/X _17705_/Y VGND VGND VPWR VPWR _17706_/X sky130_fd_sc_hd__or2_4
XANTENNA__13155__A _12740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14918_ _11838_/Y _11614_/X _14887_/X _11592_/X _14917_/X VGND VGND VPWR VPWR _14918_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_3_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18686_ _18610_/A _17111_/X _18685_/Y VGND VGND VPWR VPWR _18686_/X sky130_fd_sc_hd__o21a_4
XFILLER_75_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15898_ _15879_/A _15828_/B VGND VGND VPWR VPWR _15900_/B sky130_fd_sc_hd__or2_4
XANTENNA__22468__A _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23076__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17637_ _16935_/X _17004_/X _17006_/X _17636_/X VGND VGND VPWR VPWR _17637_/X sky130_fd_sc_hd__o22a_4
X_14849_ _14040_/X _14833_/X _14848_/X VGND VGND VPWR VPWR _14850_/C sky130_fd_sc_hd__or3_4
XFILLER_90_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15370__A _14010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17568_ _17567_/X VGND VGND VPWR VPWR _17568_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14785__A2 _13595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19307_ _18864_/C _24140_/Q _17040_/A _19306_/Y VGND VGND VPWR VPWR _19308_/A sky130_fd_sc_hd__o22a_4
X_16519_ _16519_/A _16518_/X VGND VGND VPWR VPWR _16520_/B sky130_fd_sc_hd__or2_4
XFILLER_17_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17499_ _17175_/Y _17498_/X VGND VGND VPWR VPWR _17499_/X sky130_fd_sc_hd__or2_4
XFILLER_20_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18920__A1 _15119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18920__B2 _18892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19238_ _24285_/Q _19234_/B _19236_/Y VGND VGND VPWR VPWR _24285_/D sky130_fd_sc_hd__o21a_4
XFILLER_118_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19927__D _19926_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17297__A _14719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19169_ _19169_/A VGND VGND VPWR VPWR _19169_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21200_ _20819_/X _21197_/X _23943_/Q _21194_/X VGND VGND VPWR VPWR _21200_/X sky130_fd_sc_hd__o22a_4
X_22180_ _22112_/X _22179_/X _15758_/B _22176_/X VGND VGND VPWR VPWR _22180_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21131_ _20487_/X _21126_/X _12628_/B _21130_/X VGND VGND VPWR VPWR _21131_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20491__B1 _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12234__A _12233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22232__A1 _22117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21035__A2 _21030_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21062_ _21061_/X VGND VGND VPWR VPWR _21067_/A sky130_fd_sc_hd__buf_2
XFILLER_8_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22232__B2 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20013_ _20013_/A VGND VGND VPWR VPWR _20013_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20170__B _20169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12888__B _12945_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18739__A1 _18203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22535__A2 _22529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21964_ _21861_/X _21959_/X _23520_/Q _21920_/X VGND VGND VPWR VPWR _23520_/D sky130_fd_sc_hd__o22a_4
XFILLER_66_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20915_ _20915_/A VGND VGND VPWR VPWR _21855_/A sky130_fd_sc_hd__buf_2
X_23703_ _23316_/CLK _23703_/D VGND VGND VPWR VPWR _16219_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_82_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21895_ _21828_/X _21894_/X _15674_/B _21891_/X VGND VGND VPWR VPWR _21895_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23569__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15280__A _11976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23634_ _23155_/CLK _23634_/D VGND VGND VPWR VPWR _13046_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _20644_/A _20846_/B VGND VGND VPWR VPWR _20846_/X sky130_fd_sc_hd__and2_4
XANTENNA__22299__B2 _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15973__A1 _11852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14608__B _14689_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23565_ _23826_/CLK _21896_/X VGND VGND VPWR VPWR _15861_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19687__A _19873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20777_ _24201_/Q _20751_/X _20776_/X VGND VGND VPWR VPWR _20778_/A sky130_fd_sc_hd__o21a_4
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18911__A1 _14425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22516_ _22516_/A VGND VGND VPWR VPWR _22521_/A sky130_fd_sc_hd__buf_2
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23496_ _23079_/CLK _22004_/X VGND VGND VPWR VPWR _13698_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23002__A _23001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22447_ _22423_/A VGND VGND VPWR VPWR _22447_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12200_ _11610_/A VGND VGND VPWR VPWR _13983_/A sky130_fd_sc_hd__buf_2
XANTENNA__17478__A1 _16640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13180_ _15687_/A _13178_/X _13179_/X VGND VGND VPWR VPWR _13180_/X sky130_fd_sc_hd__and3_4
XANTENNA__18675__B1 _18206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21274__A2 _21271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22378_ _22141_/X _22375_/X _15263_/B _22372_/X VGND VGND VPWR VPWR _23266_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14343__B _14269_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12131_ _12167_/A _24029_/Q VGND VGND VPWR VPWR _12131_/X sky130_fd_sc_hd__or2_4
X_24117_ _24202_/CLK _20069_/Y HRESETn VGND VGND VPWR VPWR _24117_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20482__B1 _20288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21329_ _21263_/X _21326_/X _23884_/Q _21323_/X VGND VGND VPWR VPWR _23884_/D sky130_fd_sc_hd__o22a_4
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12062_ _11924_/A VGND VGND VPWR VPWR _12096_/A sky130_fd_sc_hd__buf_2
X_24048_ _23983_/CLK _24048_/D VGND VGND VPWR VPWR _24048_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18427__B1 _17261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22223__A1 _22100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22223__B2 _22219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15455__A _15487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16870_ _16870_/A _16870_/B _16868_/X _16870_/D VGND VGND VPWR VPWR _16870_/X sky130_fd_sc_hd__and4_4
XFILLER_46_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22338__A2_N _22337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15821_ _12851_/A _15821_/B VGND VGND VPWR VPWR _15821_/X sky130_fd_sc_hd__or2_4
XFILLER_93_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18540_ _17422_/B _18539_/X VGND VGND VPWR VPWR _18540_/Y sky130_fd_sc_hd__nand2_4
XFILLER_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15752_ _12777_/X _15752_/B _15751_/X VGND VGND VPWR VPWR _15752_/X sky130_fd_sc_hd__and3_4
X_12964_ _12964_/A _12964_/B _12963_/X VGND VGND VPWR VPWR _12972_/B sky130_fd_sc_hd__or3_4
X_14703_ _11697_/A _14703_/B VGND VGND VPWR VPWR _14703_/X sky130_fd_sc_hd__or2_4
XFILLER_61_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11915_ _11915_/A VGND VGND VPWR VPWR _15986_/A sky130_fd_sc_hd__buf_2
X_18471_ _18424_/X _18269_/Y _18249_/X _18470_/Y VGND VGND VPWR VPWR _18471_/X sky130_fd_sc_hd__a211o_4
X_15683_ _12240_/X _15748_/B VGND VGND VPWR VPWR _15684_/C sky130_fd_sc_hd__or2_4
XFILLER_45_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15902__B _15902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12895_ _12895_/A _23955_/Q VGND VGND VPWR VPWR _12895_/X sky130_fd_sc_hd__or2_4
XFILLER_79_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17422_ _17422_/A _17422_/B _17422_/C _17422_/D VGND VGND VPWR VPWR _17423_/B sky130_fd_sc_hd__or4_4
XANTENNA__15190__A _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13703__A _15487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14634_ _15036_/A _14706_/B VGND VGND VPWR VPWR _14634_/X sky130_fd_sc_hd__or2_4
X_11846_ _13987_/A VGND VGND VPWR VPWR _11847_/A sky130_fd_sc_hd__buf_2
X_17353_ _16910_/A _17364_/A _17365_/A VGND VGND VPWR VPWR _17354_/B sky130_fd_sc_hd__o21a_4
XFILLER_14_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21920__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11777_ _11691_/X VGND VGND VPWR VPWR _11782_/A sky130_fd_sc_hd__buf_2
X_14565_ _14563_/X VGND VGND VPWR VPWR _14565_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17166__B1 _17165_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12319__A _14322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18902__A1 _15911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16304_ _16185_/A _16240_/B VGND VGND VPWR VPWR _16306_/B sky130_fd_sc_hd__or2_4
X_13516_ _13511_/X _13516_/B _13515_/X VGND VGND VPWR VPWR _13517_/C sky130_fd_sc_hd__and3_4
X_17284_ _17533_/A VGND VGND VPWR VPWR _17287_/A sky130_fd_sc_hd__inv_2
X_14496_ _13845_/A VGND VGND VPWR VPWR _14533_/A sky130_fd_sc_hd__buf_2
XANTENNA__20536__A _22100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19023_ _19016_/X _19022_/X _19016_/X _24335_/Q VGND VGND VPWR VPWR _24335_/D sky130_fd_sc_hd__a2bb2o_4
X_16235_ _16234_/Y VGND VGND VPWR VPWR _16235_/X sky130_fd_sc_hd__buf_2
X_13447_ _12910_/A VGND VGND VPWR VPWR _13447_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13378_ _12829_/A VGND VGND VPWR VPWR _13378_/X sky130_fd_sc_hd__buf_2
X_16166_ _16202_/A _23735_/Q VGND VGND VPWR VPWR _16167_/C sky130_fd_sc_hd__or2_4
X_15117_ _14040_/X _15101_/X _15117_/C VGND VGND VPWR VPWR _15118_/C sky130_fd_sc_hd__or3_4
X_12329_ _12711_/A _12329_/B VGND VGND VPWR VPWR _12330_/C sky130_fd_sc_hd__or2_4
X_16097_ _16097_/A _16171_/B VGND VGND VPWR VPWR _16098_/C sky130_fd_sc_hd__or2_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15048_ _14128_/A _15025_/X _15032_/X _15039_/X _15047_/X VGND VGND VPWR VPWR _15048_/X
+ sky130_fd_sc_hd__a32o_4
X_19925_ _22985_/A VGND VGND VPWR VPWR _19925_/X sky130_fd_sc_hd__buf_2
XANTENNA__12989__A _12989_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11893__A _15023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19856_ _19603_/A _19556_/Y _19562_/X _19855_/X VGND VGND VPWR VPWR _19856_/X sky130_fd_sc_hd__a211o_4
XFILLER_96_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18807_ _15379_/X _18802_/X _24418_/Q _18803_/X VGND VGND VPWR VPWR _24418_/D sky130_fd_sc_hd__o22a_4
X_19787_ _19813_/A VGND VGND VPWR VPWR _19787_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16999_ _17680_/A _16977_/B _16999_/C _16985_/X VGND VGND VPWR VPWR _18013_/B sky130_fd_sc_hd__or4_4
XFILLER_96_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18676__A _18066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18738_ _18735_/X _18737_/X _18486_/X VGND VGND VPWR VPWR _18751_/A sky130_fd_sc_hd__a21o_4
XFILLER_77_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19394__B2 _24205_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18669_ _18653_/X _11625_/X _18668_/Y _24451_/Q _18605_/X VGND VGND VPWR VPWR _24451_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16196__A _16227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20700_ _20342_/B _20754_/B VGND VGND VPWR VPWR _20701_/C sky130_fd_sc_hd__or2_4
XFILLER_97_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21680_ _21574_/X _21676_/X _23681_/Q _21637_/X VGND VGND VPWR VPWR _21680_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22926__A _22968_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20631_ _18407_/X _20447_/X _20492_/X _20630_/Y VGND VGND VPWR VPWR _20631_/X sky130_fd_sc_hd__a211o_4
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12229__A _12691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16924__A _16923_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23350_ _23313_/CLK _23350_/D VGND VGND VPWR VPWR _12222_/B sky130_fd_sc_hd__dfxtp_4
X_20562_ _20301_/A VGND VGND VPWR VPWR _20562_/X sky130_fd_sc_hd__buf_2
XFILLER_109_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22301_ _12146_/B VGND VGND VPWR VPWR _23325_/D sky130_fd_sc_hd__buf_2
X_23281_ _23313_/CLK _23281_/D VGND VGND VPWR VPWR _13149_/B sky130_fd_sc_hd__dfxtp_4
X_20493_ _20493_/A VGND VGND VPWR VPWR _20493_/X sky130_fd_sc_hd__buf_2
XFILLER_69_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14444__A _12862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22232_ _22117_/X _22229_/X _15432_/B _22226_/X VGND VGND VPWR VPWR _22232_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22453__B2 _22447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22163_ _22083_/X _22158_/X _16424_/B _22162_/X VGND VGND VPWR VPWR _22163_/X sky130_fd_sc_hd__o22a_4
X_21114_ _21118_/A VGND VGND VPWR VPWR _21130_/A sky130_fd_sc_hd__inv_2
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22094_ _22093_/X _22089_/X _12276_/B _22084_/X VGND VGND VPWR VPWR _23446_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12899__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21045_ _20779_/X _21044_/X _24041_/Q _21041_/X VGND VGND VPWR VPWR _24041_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15275__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19970__A _19994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17632__A1 _17261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_HCLK_A clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22508__A2 _22507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22996_ _22995_/X VGND VGND VPWR VPWR HADDR[19] sky130_fd_sc_hd__inv_2
XANTENNA__15722__B _15722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21947_ _21831_/X _21945_/X _15802_/B _21942_/X VGND VGND VPWR VPWR _21947_/X sky130_fd_sc_hd__o22a_4
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14619__A _13927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21192__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11700_ _12360_/A VGND VGND VPWR VPWR _11700_/X sky130_fd_sc_hd__buf_2
XFILLER_54_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13523__A _12980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12434_/X _12680_/B VGND VGND VPWR VPWR _13586_/A sky130_fd_sc_hd__or2_4
XFILLER_42_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ _21799_/X _21873_/X _16405_/B _21877_/X VGND VGND VPWR VPWR _21878_/X sky130_fd_sc_hd__o22a_4
XFILLER_58_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A VGND VGND VPWR VPWR _17054_/A sky130_fd_sc_hd__buf_2
XANTENNA__21740__A _21740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _20733_/X _20828_/X _11511_/A _20686_/X VGND VGND VPWR VPWR _20829_/X sky130_fd_sc_hd__o22a_4
X_23617_ _23819_/CLK _21780_/X VGND VGND VPWR VPWR _23617_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19688__A2 _19829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _20558_/A IRQ[18] VGND VGND VPWR VPWR _20156_/A sky130_fd_sc_hd__and2_4
X_14350_ _15616_/A _14350_/B _14350_/C VGND VGND VPWR VPWR _14351_/C sky130_fd_sc_hd__and3_4
XANTENNA__21495__A2 _21491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23548_ _24026_/CLK _21926_/X VGND VGND VPWR VPWR _23548_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22692__B2 _22690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13301_ _13301_/A _23984_/Q VGND VGND VPWR VPWR _13302_/C sky130_fd_sc_hd__or2_4
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14281_ _15558_/A _14277_/X _14280_/X VGND VGND VPWR VPWR _14281_/X sky130_fd_sc_hd__or3_4
XFILLER_17_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11978__A _11977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23479_ _23539_/CLK _22033_/X VGND VGND VPWR VPWR _23479_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13232_ _13256_/A _13157_/B VGND VGND VPWR VPWR _13234_/B sky130_fd_sc_hd__or2_4
X_16020_ _16047_/A _23768_/Q VGND VGND VPWR VPWR _16020_/X sky130_fd_sc_hd__or2_4
XFILLER_109_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19845__C1 _19876_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15169__B _15240_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22571__A _22600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18112__A2 _17922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13163_ _12711_/A _23569_/Q VGND VGND VPWR VPWR _13164_/C sky130_fd_sc_hd__or2_4
XFILLER_87_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22995__A2 _17672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16123__A1 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19860__A2 _19859_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12114_ _11992_/X _12089_/X _12096_/X _12105_/X _12113_/X VGND VGND VPWR VPWR _12114_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20803__B _20556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24357__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21187__A _21180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13094_ _13119_/A _23666_/Q VGND VGND VPWR VPWR _13094_/X sky130_fd_sc_hd__or2_4
X_17971_ _17971_/A VGND VGND VPWR VPWR _17971_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19710_ _19449_/A VGND VGND VPWR VPWR _19710_/X sky130_fd_sc_hd__buf_2
XFILLER_78_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12045_ _11888_/A VGND VGND VPWR VPWR _12083_/A sky130_fd_sc_hd__buf_2
X_16922_ _11585_/A _17285_/A _11580_/Y _16921_/X VGND VGND VPWR VPWR _17105_/A sky130_fd_sc_hd__or4_4
XANTENNA__12602__A _13726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_13_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_13_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19641_ _19624_/A VGND VGND VPWR VPWR _19744_/B sky130_fd_sc_hd__inv_2
XFILLER_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16853_ _15914_/B _16835_/X _15914_/B _16835_/X VGND VGND VPWR VPWR _16853_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15804_ _12876_/A _15800_/X _15804_/C VGND VGND VPWR VPWR _15804_/X sky130_fd_sc_hd__or3_4
XFILLER_24_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19572_ _19744_/A _19572_/B _19572_/C VGND VGND VPWR VPWR _19573_/A sky130_fd_sc_hd__or3_4
XFILLER_65_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16784_ _16803_/A _23611_/Q VGND VGND VPWR VPWR _16784_/X sky130_fd_sc_hd__or2_4
X_13996_ _12568_/A _23498_/Q VGND VGND VPWR VPWR _13997_/C sky130_fd_sc_hd__or2_4
X_18523_ _17103_/X _18213_/Y _17933_/A _18522_/X VGND VGND VPWR VPWR _18523_/X sky130_fd_sc_hd__a211o_4
XANTENNA__19376__B2 _24214_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15735_ _11741_/X _15735_/B _15734_/X VGND VGND VPWR VPWR _15735_/X sky130_fd_sc_hd__or3_4
XFILLER_111_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15632__B _23691_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12947_ _12947_/A _12945_/X _12946_/X VGND VGND VPWR VPWR _12948_/C sky130_fd_sc_hd__and3_4
XANTENNA__23884__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14529__A _13754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22380__B1 _14868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13433__A _11861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18454_ _18314_/X _18439_/Y _18357_/X _18453_/X VGND VGND VPWR VPWR _18454_/X sky130_fd_sc_hd__o22a_4
X_15666_ _15685_/A _15737_/B VGND VGND VPWR VPWR _15668_/B sky130_fd_sc_hd__or2_4
X_12878_ _12878_/A VGND VGND VPWR VPWR _12879_/A sky130_fd_sc_hd__buf_2
X_17405_ _14074_/A _17013_/A _17013_/A _17404_/X VGND VGND VPWR VPWR _17407_/B sky130_fd_sc_hd__a2bb2o_4
X_14617_ _14617_/A VGND VGND VPWR VPWR _14734_/A sky130_fd_sc_hd__buf_2
X_11829_ _11829_/A _24094_/Q VGND VGND VPWR VPWR _11830_/C sky130_fd_sc_hd__or2_4
X_18385_ _18354_/B _18383_/X _18354_/A _18384_/X VGND VGND VPWR VPWR _18385_/X sky130_fd_sc_hd__o22a_4
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17139__B1 _17007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15597_ _15643_/A _15589_/X _15597_/C VGND VGND VPWR VPWR _15613_/B sky130_fd_sc_hd__and3_4
XFILLER_14_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _17618_/C _17336_/B _17307_/Y _17335_/X VGND VGND VPWR VPWR _17337_/A sky130_fd_sc_hd__or4_4
XFILLER_33_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14548_ _14536_/A _14484_/B VGND VGND VPWR VPWR _14549_/C sky130_fd_sc_hd__or2_4
XANTENNA__21486__A2 _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11888__A _11888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17267_ _17266_/X _17781_/B VGND VGND VPWR VPWR _17267_/X sky130_fd_sc_hd__and2_4
X_14479_ _13022_/A _14479_/B VGND VGND VPWR VPWR _14479_/X sky130_fd_sc_hd__or2_4
XANTENNA__14264__A _14174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19006_ _19002_/X _19005_/X _19002_/X _24338_/Q VGND VGND VPWR VPWR _19006_/X sky130_fd_sc_hd__a2bb2o_4
X_16218_ _16206_/A _16216_/X _16217_/X VGND VGND VPWR VPWR _16222_/B sky130_fd_sc_hd__and3_4
XANTENNA__21238__A2 _21235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15079__B _15079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17198_ _17151_/X _17189_/X _17817_/A _17197_/X VGND VGND VPWR VPWR _17198_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__23264__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19300__A1 _23064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12923__A1 _11980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20446__B1 _20284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16149_ _16145_/A _16219_/B VGND VGND VPWR VPWR _16149_/X sky130_fd_sc_hd__or2_4
XFILLER_66_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19908_ _19899_/X _24153_/Q _19903_/X _20358_/B VGND VGND VPWR VPWR _24153_/D sky130_fd_sc_hd__o22a_4
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12512__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20749__A1 _20613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20749__B2 _20724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19839_ _19839_/A _19839_/B VGND VGND VPWR VPWR _19839_/X sky130_fd_sc_hd__or2_4
XFILLER_112_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15823__A _15823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22850_ _17283_/Y _22778_/Y _22794_/A VGND VGND VPWR VPWR _22850_/X sky130_fd_sc_hd__o21a_4
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16638__B _23996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21801_ _21799_/X _21793_/X _23610_/Q _21800_/X VGND VGND VPWR VPWR _23610_/D sky130_fd_sc_hd__o22a_4
XFILLER_65_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22781_ _22781_/A VGND VGND VPWR VPWR _22781_/X sky130_fd_sc_hd__buf_2
XANTENNA__14439__A _12441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21174__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17917__A2 _17913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13343__A _15784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21732_ _21578_/X _21705_/A _23647_/Q _21687_/X VGND VGND VPWR VPWR _21732_/X sky130_fd_sc_hd__o22a_4
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21663_ _21543_/X _21662_/X _15765_/B _21659_/X VGND VGND VPWR VPWR _23694_/D sky130_fd_sc_hd__o22a_4
X_24451_ _24229_/CLK _24451_/D HRESETn VGND VGND VPWR VPWR _24451_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20614_ _20512_/A VGND VGND VPWR VPWR _20614_/X sky130_fd_sc_hd__buf_2
X_23402_ _24011_/CLK _22185_/X VGND VGND VPWR VPWR _13970_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_71_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19030__A _19002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24382_ _24435_/CLK _24382_/D HRESETn VGND VGND VPWR VPWR _24382_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22674__A1 _21795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21594_ _21512_/X _21591_/X _23739_/Q _21588_/X VGND VGND VPWR VPWR _23739_/D sky130_fd_sc_hd__o22a_4
XFILLER_36_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22674__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23333_ _23973_/CLK _23333_/D VGND VGND VPWR VPWR _14501_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__11798__A _11798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20545_ _20493_/X _20544_/X _24306_/Q _20500_/X VGND VGND VPWR VPWR _20546_/B sky130_fd_sc_hd__o22a_4
XFILLER_20_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23264_ _24032_/CLK _23264_/D VGND VGND VPWR VPWR _14868_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20476_ _20468_/X _20475_/Y _24277_/Q _20301_/X VGND VGND VPWR VPWR _20476_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22426__B2 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22391__A _22384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20437__B1 _20288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22215_ _22222_/A VGND VGND VPWR VPWR _22215_/X sky130_fd_sc_hd__buf_2
X_23195_ _23260_/CLK _22525_/X VGND VGND VPWR VPWR _16754_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_69_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14902__A _15146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23757__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22146_ _22145_/X _22137_/X _14883_/B _22071_/X VGND VGND VPWR VPWR _22146_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13518__A _13572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22077_ _22101_/A VGND VGND VPWR VPWR _22077_/X sky130_fd_sc_hd__buf_2
XFILLER_59_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12422__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21028_ _20487_/X _21023_/X _12643_/B _21027_/X VGND VGND VPWR VPWR _24053_/D sky130_fd_sc_hd__o22a_4
XFILLER_87_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15733__A _12795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13850_ _15314_/A VGND VGND VPWR VPWR _13851_/A sky130_fd_sc_hd__buf_2
XFILLER_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12801_ _12754_/X _12799_/X _12801_/C VGND VGND VPWR VPWR _12805_/B sky130_fd_sc_hd__and3_4
X_13781_ _13608_/A _23719_/Q VGND VGND VPWR VPWR _13781_/X sky130_fd_sc_hd__or2_4
XFILLER_90_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22979_ _23003_/A _22979_/B VGND VGND VPWR VPWR _22979_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22362__B1 _15725_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15520_ _15519_/X VGND VGND VPWR VPWR _15520_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13253__A _13260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12732_ _12706_/A _12732_/B _12732_/C VGND VGND VPWR VPWR _12732_/X sky130_fd_sc_hd__or3_4
XFILLER_43_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18046__A1_N _18425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21470__A _21470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15451_ _11977_/X _15428_/X _15435_/X _15442_/X _15450_/X VGND VGND VPWR VPWR _15451_/X
+ sky130_fd_sc_hd__a32o_4
X_12663_ _12955_/A _12663_/B _12662_/X VGND VGND VPWR VPWR _12663_/X sky130_fd_sc_hd__or3_4
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _15637_/A _23398_/Q VGND VGND VPWR VPWR _14402_/X sky130_fd_sc_hd__or2_4
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _15047_/A _14995_/A _12860_/A _13651_/A VGND VGND VPWR VPWR _11614_/X sky130_fd_sc_hd__or4_4
X_18170_ _18129_/X _18169_/X _19995_/A _18129_/X VGND VGND VPWR VPWR _24470_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21468__A2 _21463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_4_0_HCLK clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _15312_/X _15381_/X VGND VGND VPWR VPWR _15382_/X sky130_fd_sc_hd__and2_4
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12937_/A VGND VGND VPWR VPWR _12640_/A sky130_fd_sc_hd__buf_2
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16283__B _16283_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ _22017_/A VGND VGND VPWR VPWR _21007_/A sky130_fd_sc_hd__inv_2
XFILLER_51_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14333_ _15398_/A _14329_/X _14332_/X VGND VGND VPWR VPWR _14333_/X sky130_fd_sc_hd__or3_4
X_11545_ _20520_/A IRQ[20] VGND VGND VPWR VPWR _20158_/A sky130_fd_sc_hd__and2_4
XFILLER_7_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ _17052_/A _16916_/B VGND VGND VPWR VPWR _17052_/X sky130_fd_sc_hd__or2_4
XFILLER_32_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14264_ _14174_/X _14263_/A VGND VGND VPWR VPWR _14265_/A sky130_fd_sc_hd__or2_4
XANTENNA__22417__B2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12316__B _12316_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16003_ _11915_/A _16003_/B _16002_/X VGND VGND VPWR VPWR _16003_/X sky130_fd_sc_hd__and3_4
X_13215_ _13228_/A _24017_/Q VGND VGND VPWR VPWR _13217_/B sky130_fd_sc_hd__or2_4
XANTENNA__15908__A _15907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14195_ _14195_/A _14195_/B _14195_/C VGND VGND VPWR VPWR _14201_/B sky130_fd_sc_hd__and3_4
XANTENNA__14812__A _13690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13146_ _12720_/A _13144_/X _13145_/X VGND VGND VPWR VPWR _13146_/X sky130_fd_sc_hd__and3_4
XFILLER_98_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13428__A _13428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13077_ _13088_/A VGND VGND VPWR VPWR _13119_/A sky130_fd_sc_hd__buf_2
X_17954_ _18062_/A _17627_/A VGND VGND VPWR VPWR _17954_/X sky130_fd_sc_hd__or2_4
XFILLER_65_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12332__A _12315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12028_ _11992_/X _11999_/X _12006_/X _12017_/X _12027_/X VGND VGND VPWR VPWR _12028_/X
+ sky130_fd_sc_hd__a32o_4
X_16905_ _16897_/A _16904_/Y _16897_/A _16904_/Y VGND VGND VPWR VPWR _16905_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21645__A _21637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17885_ _16927_/X _17881_/X _17639_/X _17884_/X VGND VGND VPWR VPWR _17885_/X sky130_fd_sc_hd__o22a_4
XFILLER_26_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16739__A _11966_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15643__A _15643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16836_ _15914_/B _16835_/X _15650_/A VGND VGND VPWR VPWR _16836_/X sky130_fd_sc_hd__o21a_4
X_19624_ _19624_/A _19623_/X VGND VGND VPWR VPWR _19624_/Y sky130_fd_sc_hd__nor2_4
XFILLER_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19555_ _20342_/B _19551_/X _19553_/X _19554_/X VGND VGND VPWR VPWR _19555_/X sky130_fd_sc_hd__a211o_4
X_16767_ _16803_/A _16767_/B VGND VGND VPWR VPWR _16767_/X sky130_fd_sc_hd__or2_4
XFILLER_59_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13979_ _12302_/A _13979_/B _13978_/X VGND VGND VPWR VPWR _13979_/X sky130_fd_sc_hd__or3_4
XANTENNA__14259__A _11669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21156__B2 _21151_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18506_ _18487_/X _18494_/Y _18495_/X _18497_/X _18505_/Y VGND VGND VPWR VPWR _18506_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13163__A _12711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15718_ _15725_/A _15656_/B VGND VGND VPWR VPWR _15719_/C sky130_fd_sc_hd__or2_4
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19486_ _19691_/A VGND VGND VPWR VPWR _19486_/Y sky130_fd_sc_hd__inv_2
X_16698_ _16698_/A _23995_/Q VGND VGND VPWR VPWR _16699_/C sky130_fd_sc_hd__or2_4
XANTENNA__22476__A _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21380__A _21373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18437_ _18344_/X _16974_/B _18414_/Y VGND VGND VPWR VPWR _18437_/Y sky130_fd_sc_hd__a21oi_4
X_15649_ _15582_/X _15649_/B VGND VGND VPWR VPWR _15650_/A sky130_fd_sc_hd__or2_4
XFILLER_72_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18368_ _17864_/X _18144_/X _17823_/X _18116_/X VGND VGND VPWR VPWR _18368_/X sky130_fd_sc_hd__o22a_4
XFILLER_72_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22656__B2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17319_ _17143_/X _17201_/A VGND VGND VPWR VPWR _18658_/A sky130_fd_sc_hd__and2_4
XANTENNA__20667__B1 _20666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18299_ _18298_/X VGND VGND VPWR VPWR _18299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12507__A _13031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20330_ _20500_/A VGND VGND VPWR VPWR _20330_/X sky130_fd_sc_hd__buf_2
XFILLER_116_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20724__A _20488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20261_ _24414_/Q _18814_/X _24446_/Q _20260_/X VGND VGND VPWR VPWR _20261_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18088__B2 _18087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15818__A _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22000_ _21835_/X _21995_/X _23499_/Q _21999_/X VGND VGND VPWR VPWR _22000_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21092__B1 _15465_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22722__A2_N _19303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20192_ _21581_/A _21296_/A _21583_/A _21212_/A VGND VGND VPWR VPWR _20193_/A sky130_fd_sc_hd__or4_4
XFILLER_66_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21631__A2 _21626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15537__B _23979_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24340__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13338__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12242__A _12695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23951_ _24047_/CLK _23951_/D VGND VGND VPWR VPWR _13540_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_69_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16649__A _16616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21395__B2 _21359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22592__B1 _13456_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22902_ _23051_/A _18644_/A _22901_/X VGND VGND VPWR VPWR _22902_/X sky130_fd_sc_hd__or3_4
XFILLER_84_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23882_ _23915_/CLK _23882_/D VGND VGND VPWR VPWR _23882_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_5_4_0_HCLK_A clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16368__B _16368_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22833_ _13350_/Y _22825_/X _22831_/X _22832_/X VGND VGND VPWR VPWR _22834_/A sky130_fd_sc_hd__a211o_4
XFILLER_77_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14169__A _15023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13073__A _12613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22764_ _22763_/A _22763_/B VGND VGND VPWR VPWR _22765_/B sky130_fd_sc_hd__or2_4
XFILLER_25_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22386__A _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21715_ _21548_/X _21712_/X _15406_/B _21709_/X VGND VGND VPWR VPWR _21715_/X sky130_fd_sc_hd__o22a_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22695_ _21831_/A _22693_/X _15835_/B _22690_/X VGND VGND VPWR VPWR _22695_/X sky130_fd_sc_hd__o22a_4
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16384__A _16002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13801__A _13659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21646_ _21514_/X _21641_/X _16437_/B _21645_/X VGND VGND VPWR VPWR _21646_/X sky130_fd_sc_hd__o22a_4
X_24434_ _23326_/CLK _18785_/X HRESETn VGND VGND VPWR VPWR _24434_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21577_ _21576_/X _21568_/X _14864_/B _21515_/A VGND VGND VPWR VPWR _23744_/D sky130_fd_sc_hd__o22a_4
X_24365_ _24365_/CLK _18902_/X HRESETn VGND VGND VPWR VPWR _24365_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__12417__A _15889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20528_ _20517_/X _20526_/X _19128_/A _20527_/X VGND VGND VPWR VPWR _20529_/B sky130_fd_sc_hd__o22a_4
X_23316_ _23316_/CLK _23316_/D VGND VGND VPWR VPWR _23316_/Q sky130_fd_sc_hd__dfxtp_4
X_24296_ _24299_/CLK _24296_/D HRESETn VGND VGND VPWR VPWR _24296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12136__B _23933_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23010__A _18193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15728__A _13133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20459_ _20459_/A VGND VGND VPWR VPWR _20459_/X sky130_fd_sc_hd__buf_2
X_23247_ _23827_/CLK _23247_/D VGND VGND VPWR VPWR _13427_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14632__A _13927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21449__B _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18104__A _18297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13000_ _12890_/A _12998_/X _12999_/X VGND VGND VPWR VPWR _13000_/X sky130_fd_sc_hd__and3_4
X_23178_ _23978_/CLK _23178_/D VGND VGND VPWR VPWR _14011_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21622__A2 _21619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15447__B _23852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22129_ _22129_/A VGND VGND VPWR VPWR _22129_/X sky130_fd_sc_hd__buf_2
XANTENNA__13248__A _13260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12115__A2 _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14951_ _14925_/A _14949_/X _14951_/C VGND VGND VPWR VPWR _14952_/C sky130_fd_sc_hd__and3_4
XANTENNA__17662__B _17662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16559__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21386__B2 _21380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13902_ _13890_/A _23079_/Q VGND VGND VPWR VPWR _13904_/B sky130_fd_sc_hd__or2_4
XANTENNA__15463__A _15487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17670_ _16948_/Y _17497_/X VGND VGND VPWR VPWR _17684_/A sky130_fd_sc_hd__or2_4
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14882_ _14912_/A _14882_/B VGND VGND VPWR VPWR _14882_/X sky130_fd_sc_hd__or2_4
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16621_ _16621_/A _16621_/B _16621_/C VGND VGND VPWR VPWR _16622_/C sky130_fd_sc_hd__and3_4
X_13833_ _13632_/A _13833_/B _13832_/X VGND VGND VPWR VPWR _13833_/X sky130_fd_sc_hd__and3_4
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14079__A _14906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21138__B2 _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18774__A _18781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19340_ _19336_/A VGND VGND VPWR VPWR _19340_/X sky130_fd_sc_hd__buf_2
X_16552_ _16583_/A _23548_/Q VGND VGND VPWR VPWR _16553_/C sky130_fd_sc_hd__or2_4
X_13764_ _12937_/A _24072_/Q VGND VGND VPWR VPWR _13765_/C sky130_fd_sc_hd__or2_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15503_ _15491_/A _15501_/X _15503_/C VGND VGND VPWR VPWR _15503_/X sky130_fd_sc_hd__and3_4
X_12715_ _12682_/X _12689_/X _12696_/X _12706_/X _12714_/X VGND VGND VPWR VPWR _12715_/X
+ sky130_fd_sc_hd__a32o_4
X_19271_ _19218_/B VGND VGND VPWR VPWR _19271_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20897__B1 HRDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16483_ _16465_/A _23962_/Q VGND VGND VPWR VPWR _16484_/C sky130_fd_sc_hd__or2_4
X_13695_ _13890_/A VGND VGND VPWR VPWR _13695_/X sky130_fd_sc_hd__buf_2
XANTENNA__20361__A2 _18814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14807__A _12599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18222_ _18204_/X _18209_/Y _18215_/X _18220_/X _18221_/Y VGND VGND VPWR VPWR _18222_/X
+ sky130_fd_sc_hd__a32o_4
X_15434_ _15411_/A _15434_/B _15433_/X VGND VGND VPWR VPWR _15435_/C sky130_fd_sc_hd__and3_4
X_12646_ _12646_/A VGND VGND VPWR VPWR _12951_/A sky130_fd_sc_hd__buf_2
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23922__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22638__B2 _22633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ _18153_/A VGND VGND VPWR VPWR _18153_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15365_ _15325_/X _15365_/B _15365_/C VGND VGND VPWR VPWR _15365_/X sky130_fd_sc_hd__and3_4
X_12577_ _12638_/A VGND VGND VPWR VPWR _12970_/A sky130_fd_sc_hd__buf_2
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12327__A _12320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21310__B2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17104_ _19823_/A VGND VGND VPWR VPWR _21005_/A sky130_fd_sc_hd__inv_2
X_14316_ _15576_/A VGND VGND VPWR VPWR _14431_/A sky130_fd_sc_hd__buf_2
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _11528_/A _11527_/X VGND VGND VPWR VPWR _11528_/X sky130_fd_sc_hd__or2_4
X_18084_ _17989_/X _17564_/X _18081_/X _18082_/X _18083_/Y VGND VGND VPWR VPWR _18085_/B
+ sky130_fd_sc_hd__a32o_4
X_15296_ _12439_/A _15296_/B VGND VGND VPWR VPWR _15296_/X sky130_fd_sc_hd__or2_4
XANTENNA__12046__B _12123_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17035_ _17034_/Y _17467_/B VGND VGND VPWR VPWR _17342_/A sky130_fd_sc_hd__or2_4
X_14247_ _14247_/A _23689_/Q VGND VGND VPWR VPWR _14249_/B sky130_fd_sc_hd__or2_4
XANTENNA__14542__A _13695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21074__B1 _24025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21613__A2 _21612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14178_ _14178_/A VGND VGND VPWR VPWR _14197_/A sky130_fd_sc_hd__buf_2
XFILLER_28_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13158__A _15707_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13129_ _13129_/A _13045_/B VGND VGND VPWR VPWR _13129_/X sky130_fd_sc_hd__or2_4
XFILLER_119_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12062__A _11924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18986_ _18965_/X _18984_/X _18985_/Y _18968_/X VGND VGND VPWR VPWR _18986_/X sky130_fd_sc_hd__o22a_4
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17937_ _17862_/X _17936_/X _17869_/X VGND VGND VPWR VPWR _17937_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16469__A _16194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21377__B2 _21373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15373__A _14000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17868_ _17868_/A VGND VGND VPWR VPWR _17868_/X sky130_fd_sc_hd__buf_2
XFILLER_66_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20585__C1 _20584_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24129__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19607_ _19521_/X VGND VGND VPWR VPWR _19607_/X sky130_fd_sc_hd__buf_2
XFILLER_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16819_ _16525_/X _16817_/X _16898_/A VGND VGND VPWR VPWR _16819_/X sky130_fd_sc_hd__o21a_4
X_17799_ _17824_/A VGND VGND VPWR VPWR _17800_/A sky130_fd_sc_hd__buf_2
XFILLER_53_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21129__B2 _21123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19538_ _19538_/A VGND VGND VPWR VPWR _19817_/C sky130_fd_sc_hd__buf_2
XANTENNA__22877__A1 _12116_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19469_ _24152_/Q _19433_/Y HRDATA[26] _19433_/A VGND VGND VPWR VPWR _19469_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14717__A _15643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21500_ _21500_/A VGND VGND VPWR VPWR _21556_/A sky130_fd_sc_hd__buf_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13621__A _15424_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22480_ _22403_/X _22479_/X _15992_/B _22476_/X VGND VGND VPWR VPWR _22480_/X sky130_fd_sc_hd__o22a_4
X_21431_ _21265_/X _21426_/X _15560_/B _21430_/X VGND VGND VPWR VPWR _23819_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12237__A _12209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24150_ _24162_/CLK _24150_/D HRESETn VGND VGND VPWR VPWR _24150_/Q sky130_fd_sc_hd__dfrtp_4
X_21362_ _21369_/A VGND VGND VPWR VPWR _21362_/X sky130_fd_sc_hd__buf_2
XANTENNA__16859__A2 _15119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16651__B _24060_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20313_ _24221_/Q _20282_/X _20312_/X VGND VGND VPWR VPWR _20314_/A sky130_fd_sc_hd__o21a_4
X_23101_ _23485_/CLK _23101_/D VGND VGND VPWR VPWR _23101_/Q sky130_fd_sc_hd__dfxtp_4
X_24081_ _24082_/CLK _20575_/X VGND VGND VPWR VPWR _24081_/Q sky130_fd_sc_hd__dfxtp_4
X_21293_ _21293_/A VGND VGND VPWR VPWR _21293_/X sky130_fd_sc_hd__buf_2
XANTENNA__14452__A _12533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23032_ _23027_/A _18018_/X VGND VGND VPWR VPWR _23032_/Y sky130_fd_sc_hd__nand2_4
XFILLER_116_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20244_ _20244_/A _20500_/A VGND VGND VPWR VPWR _20270_/B sky130_fd_sc_hd__or2_4
XANTENNA__21604__A2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13068__A _13097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20175_ _18603_/Y _20133_/Y _20174_/X VGND VGND VPWR VPWR _20175_/X sky130_fd_sc_hd__o21a_4
XFILLER_88_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21368__B2 _21366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23934_ _23320_/CLK _21220_/X VGND VGND VPWR VPWR _23934_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12700__A _12711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13058__B1 _11596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23865_ _23770_/CLK _23865_/D VGND VGND VPWR VPWR _16297_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18594__A _18593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22816_ _15453_/Y _22814_/X _22795_/X _22815_/X VGND VGND VPWR VPWR _22817_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22868__A1 _16444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23945__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23796_ _23315_/CLK _21469_/X VGND VGND VPWR VPWR _23796_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20879__B1 _20490_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15730__B _15674_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22747_ _22747_/A _22732_/X _22735_/X _22746_/X VGND VGND VPWR VPWR _22747_/X sky130_fd_sc_hd__or4_4
XFILLER_73_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21540__B2 _21539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12500_ _13016_/A VGND VGND VPWR VPWR _12500_/X sky130_fd_sc_hd__buf_2
XFILLER_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13480_ _13448_/X _13568_/B VGND VGND VPWR VPWR _13480_/X sky130_fd_sc_hd__or2_4
XFILLER_40_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_66_0_HCLK clkbuf_7_66_0_HCLK/A VGND VGND VPWR VPWR _24299_/CLK sky130_fd_sc_hd__clkbuf_1
X_22678_ _21802_/A _22672_/X _16293_/B _22676_/X VGND VGND VPWR VPWR _22678_/X sky130_fd_sc_hd__o22a_4
XFILLER_13_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12431_ _12338_/Y _12430_/X VGND VGND VPWR VPWR _12434_/A sky130_fd_sc_hd__and2_4
X_24417_ _24320_/CLK _24417_/D HRESETn VGND VGND VPWR VPWR _11541_/A sky130_fd_sc_hd__dfrtp_4
X_21629_ _21572_/X _21626_/X _15256_/B _21623_/X VGND VGND VPWR VPWR _23714_/D sky130_fd_sc_hd__o22a_4
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15150_ _14990_/A _15150_/B VGND VGND VPWR VPWR _15151_/C sky130_fd_sc_hd__or2_4
X_12362_ _12398_/A _12362_/B _12361_/X VGND VGND VPWR VPWR _12362_/X sky130_fd_sc_hd__and3_4
X_24348_ _24344_/CLK _18948_/X HRESETn VGND VGND VPWR VPWR _24348_/Q sky130_fd_sc_hd__dfstp_4
X_14101_ _14101_/A VGND VGND VPWR VPWR _15010_/A sky130_fd_sc_hd__buf_2
X_12293_ _12725_/A _12293_/B VGND VGND VPWR VPWR _12293_/X sky130_fd_sc_hd__or2_4
X_15081_ _15109_/A _15081_/B VGND VGND VPWR VPWR _15083_/B sky130_fd_sc_hd__or2_4
X_24279_ _24435_/CLK _19250_/X HRESETn VGND VGND VPWR VPWR _24279_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23325__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21056__B1 _14892_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14032_ _14045_/A _23978_/Q VGND VGND VPWR VPWR _14033_/C sky130_fd_sc_hd__or2_4
XFILLER_49_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15177__B _15177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18840_ _17194_/X _18834_/X _24400_/Q _18835_/X VGND VGND VPWR VPWR _24400_/D sky130_fd_sc_hd__o22a_4
XFILLER_45_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18771_ _17266_/X _18765_/X _24444_/Q _18768_/X VGND VGND VPWR VPWR _18771_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23475__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15983_ _15994_/A _15981_/X _15983_/C VGND VGND VPWR VPWR _15987_/B sky130_fd_sc_hd__and3_4
XANTENNA__16289__A _15939_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17722_ _17718_/X VGND VGND VPWR VPWR _17723_/A sky130_fd_sc_hd__inv_2
X_14934_ _14658_/A _14934_/B _14934_/C VGND VGND VPWR VPWR _14934_/X sky130_fd_sc_hd__or3_4
XFILLER_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13706__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12610__A _13083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17653_ _16985_/A _17653_/B VGND VGND VPWR VPWR _17653_/X sky130_fd_sc_hd__or2_4
XFILLER_114_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21923__A _21919_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14865_ _12216_/A _14863_/X _14864_/X VGND VGND VPWR VPWR _14865_/X sky130_fd_sc_hd__and3_4
XFILLER_48_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16604_ _16800_/A _23516_/Q VGND VGND VPWR VPWR _16605_/C sky130_fd_sc_hd__or2_4
XFILLER_91_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13816_ _13624_/A _13814_/X _13815_/X VGND VGND VPWR VPWR _13816_/X sky130_fd_sc_hd__and3_4
X_17584_ _17447_/A _17452_/X _17454_/A VGND VGND VPWR VPWR _17584_/Y sky130_fd_sc_hd__o21ai_4
X_14796_ _13710_/A _14796_/B _14795_/X VGND VGND VPWR VPWR _14796_/X sky130_fd_sc_hd__and3_4
XFILLER_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20539__A _20285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19323_ _19321_/X _18126_/X _19321_/X _24247_/Q VGND VGND VPWR VPWR _24247_/D sky130_fd_sc_hd__a2bb2o_4
X_16535_ _16538_/A _16614_/B VGND VGND VPWR VPWR _16537_/B sky130_fd_sc_hd__or2_4
X_13747_ _13747_/A _13743_/X _13747_/C VGND VGND VPWR VPWR _13755_/B sky130_fd_sc_hd__or3_4
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15640__B _15570_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18009__A _18198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14537__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13441__A _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19254_ _24277_/Q _19225_/X _19253_/Y VGND VGND VPWR VPWR _24277_/D sky130_fd_sc_hd__o21a_4
X_16466_ _16506_/A _16464_/X _16466_/C VGND VGND VPWR VPWR _16466_/X sky130_fd_sc_hd__and3_4
X_13678_ _13678_/A _13759_/B VGND VGND VPWR VPWR _13678_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18205_ _18205_/A _17525_/B VGND VGND VPWR VPWR _18205_/X sky130_fd_sc_hd__and2_4
XFILLER_73_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15417_ _13645_/A _15474_/B VGND VGND VPWR VPWR _15418_/C sky130_fd_sc_hd__or2_4
X_12629_ _12963_/A _12629_/B _12629_/C VGND VGND VPWR VPWR _12629_/X sky130_fd_sc_hd__and3_4
X_19185_ _19117_/B VGND VGND VPWR VPWR _19185_/Y sky130_fd_sc_hd__inv_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16397_ _16100_/X VGND VGND VPWR VPWR _16397_/X sky130_fd_sc_hd__buf_2
XANTENNA__16752__A _16747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18136_ _18265_/A _17464_/B VGND VGND VPWR VPWR _18136_/Y sky130_fd_sc_hd__nor2_4
X_15348_ _13871_/A _15282_/B VGND VGND VPWR VPWR _15350_/B sky130_fd_sc_hd__or2_4
XANTENNA__21834__A2 _21829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20274__A _18577_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11896__A _14463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18067_ _18267_/A _18064_/X _18065_/X _18067_/D VGND VGND VPWR VPWR _18068_/A sky130_fd_sc_hd__or4_4
XANTENNA__15368__A _14009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15279_ _14752_/A _15279_/B _15278_/X VGND VGND VPWR VPWR _15279_/X sky130_fd_sc_hd__or3_4
XANTENNA__14272__A _12260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17018_ _17018_/A VGND VGND VPWR VPWR _17018_/X sky130_fd_sc_hd__buf_2
XANTENNA__15087__B _23871_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23818__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15815__B _15815_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18969_ _18965_/X _18966_/Y _18967_/Y _18968_/X VGND VGND VPWR VPWR _18969_/X sky130_fd_sc_hd__o22a_4
XFILLER_45_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16199__A _16215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13616__A _15424_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22011__A2 _22009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21980_ _21802_/X _21974_/X _23513_/Q _21978_/X VGND VGND VPWR VPWR _23513_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23968__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12520__A _13029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20931_ _18679_/X _20332_/A _20731_/X _20930_/Y VGND VGND VPWR VPWR _20931_/X sky130_fd_sc_hd__a211o_4
XFILLER_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21770__B2 _21766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15831__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20862_ _20715_/A _20862_/B VGND VGND VPWR VPWR _20862_/Y sky130_fd_sc_hd__nor2_4
X_23650_ _24066_/CLK _23650_/D VGND VGND VPWR VPWR _15266_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20449__A _20449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19715__A1 _19876_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22601_ _22439_/X _22600_/X _23145_/Q _22597_/X VGND VGND VPWR VPWR _23145_/D sky130_fd_sc_hd__o22a_4
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20793_ _20673_/X _20784_/Y _20791_/X _20792_/Y _20692_/X VGND VGND VPWR VPWR _20793_/X
+ sky130_fd_sc_hd__a32o_4
X_23581_ _23485_/CLK _23581_/D VGND VGND VPWR VPWR _23581_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13351__A _12813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22532_ _22408_/X _22529_/X _12228_/B _22526_/X VGND VGND VPWR VPWR _23190_/D sky130_fd_sc_hd__o22a_4
XFILLER_52_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22463_ _22462_/X _22416_/A _15052_/B _22386_/X VGND VGND VPWR VPWR _23231_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19479__B1 _19481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24202_ _24202_/CLK _19398_/X HRESETn VGND VGND VPWR VPWR _24202_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21414_ _21237_/X _21412_/X _16132_/B _21409_/X VGND VGND VPWR VPWR _21414_/X sky130_fd_sc_hd__o22a_4
X_22394_ _20338_/A VGND VGND VPWR VPWR _22394_/X sky130_fd_sc_hd__buf_2
XFILLER_87_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21825__A2 _21817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21345_ _21291_/X _21340_/X _23872_/Q _21301_/X VGND VGND VPWR VPWR _23872_/D sky130_fd_sc_hd__o22a_4
X_24133_ _24241_/CLK _19993_/Y HRESETn VGND VGND VPWR VPWR _16943_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_11_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21038__B1 _15686_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21276_ _21275_/X _21271_/X _23911_/Q _21266_/X VGND VGND VPWR VPWR _21276_/X sky130_fd_sc_hd__o22a_4
X_24064_ _24032_/CLK _24064_/D VGND VGND VPWR VPWR _14903_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23498__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18589__A _18216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21589__B2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_HCLK clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_20227_ _20226_/X VGND VGND VPWR VPWR _20286_/A sky130_fd_sc_hd__buf_2
X_23015_ _23015_/A VGND VGND VPWR VPWR _23018_/A sky130_fd_sc_hd__buf_2
XANTENNA__18454__B2 _18453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20158_ _20158_/A _20157_/Y VGND VGND VPWR VPWR _20158_/X sky130_fd_sc_hd__or2_4
XANTENNA__15725__B _15725_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12980_ _12980_/A _12980_/B VGND VGND VPWR VPWR _12982_/B sky130_fd_sc_hd__or2_4
X_20089_ _20089_/A _20087_/Y _20089_/C _20089_/D VGND VGND VPWR VPWR _20089_/X sky130_fd_sc_hd__and4_4
XANTENNA__12430__A _12429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21210__B1 _15088_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11931_ _13025_/A VGND VGND VPWR VPWR _13048_/A sky130_fd_sc_hd__buf_2
X_23917_ _23698_/CLK _23917_/D VGND VGND VPWR VPWR _15805_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19954__B2 _19953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15741__A _12792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21761__B2 _21759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14650_ _14197_/A VGND VGND VPWR VPWR _15201_/A sky130_fd_sc_hd__buf_2
XFILLER_22_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11862_ _11861_/X VGND VGND VPWR VPWR _16152_/A sky130_fd_sc_hd__buf_2
X_23848_ _23304_/CLK _21385_/X VGND VGND VPWR VPWR _13760_/B sky130_fd_sc_hd__dfxtp_4
X_13601_ _13955_/A VGND VGND VPWR VPWR _14778_/A sky130_fd_sc_hd__buf_2
XFILLER_72_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16556__B _23580_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14581_ _15144_/A _14579_/X _14581_/C VGND VGND VPWR VPWR _14581_/X sky130_fd_sc_hd__and3_4
X_11793_ _11824_/A _11793_/B _11792_/X VGND VGND VPWR VPWR _11793_/X sky130_fd_sc_hd__or3_4
X_23779_ _23494_/CLK _23779_/D VGND VGND VPWR VPWR _14777_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_92_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14357__A _15592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21513__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16320_ _13422_/A _16316_/X _16320_/C VGND VGND VPWR VPWR _16320_/X sky130_fd_sc_hd__or3_4
XANTENNA__13261__A _13242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13532_ _13529_/X _13532_/B _13532_/C VGND VGND VPWR VPWR _13536_/B sky130_fd_sc_hd__and3_4
XFILLER_57_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16251_ _16243_/X _24025_/Q VGND VGND VPWR VPWR _16251_/X sky130_fd_sc_hd__or2_4
X_13463_ _13463_/A _13540_/B VGND VGND VPWR VPWR _13464_/C sky130_fd_sc_hd__or2_4
XFILLER_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15202_ _15190_/A _23553_/Q VGND VGND VPWR VPWR _15203_/C sky130_fd_sc_hd__or2_4
X_12414_ _12384_/X _12331_/B VGND VGND VPWR VPWR _12414_/X sky130_fd_sc_hd__or2_4
X_16182_ _16202_/A _23575_/Q VGND VGND VPWR VPWR _16183_/C sky130_fd_sc_hd__or2_4
X_13394_ _13357_/X _13394_/B _13394_/C VGND VGND VPWR VPWR _13400_/B sky130_fd_sc_hd__and3_4
X_15133_ _14089_/A _23745_/Q VGND VGND VPWR VPWR _15134_/C sky130_fd_sc_hd__or2_4
X_12345_ _12373_/A VGND VGND VPWR VPWR _12794_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14092__A _14991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12605__A _12605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15064_ _15069_/A _23999_/Q VGND VGND VPWR VPWR _15064_/X sky130_fd_sc_hd__or2_4
X_19941_ _18241_/A _19941_/B VGND VGND VPWR VPWR _19944_/B sky130_fd_sc_hd__nor2_4
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12276_ _12711_/A _12276_/B VGND VGND VPWR VPWR _12276_/X sky130_fd_sc_hd__or2_4
XFILLER_68_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20822__A _20445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14015_ _14026_/A VGND VGND VPWR VPWR _14045_/A sky130_fd_sc_hd__buf_2
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19872_ _19485_/A _19872_/B _19872_/C _19881_/B VGND VGND VPWR VPWR _19872_/X sky130_fd_sc_hd__and4_4
XFILLER_116_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22241__A2 _22236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24403__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18823_ _12184_/X _18818_/X _20296_/A _18821_/X VGND VGND VPWR VPWR _24413_/D sky130_fd_sc_hd__o22a_4
XFILLER_96_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13436__A _11913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15966_ _15937_/X _15964_/X _15965_/X VGND VGND VPWR VPWR _15966_/X sky130_fd_sc_hd__and3_4
X_18754_ _17736_/A _17126_/X _17738_/X VGND VGND VPWR VPWR _18754_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_114_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14917_ _14128_/A _14894_/X _14901_/X _14908_/X _14916_/X VGND VGND VPWR VPWR _14917_/X
+ sky130_fd_sc_hd__a32o_4
X_17705_ _16956_/A _17404_/X VGND VGND VPWR VPWR _17705_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15897_ _13494_/X _15893_/X _15897_/C VGND VGND VPWR VPWR _15905_/B sky130_fd_sc_hd__or3_4
X_18685_ _17734_/X VGND VGND VPWR VPWR _18685_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20555__A2 _20939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14848_ _11669_/A _14840_/X _14848_/C VGND VGND VPWR VPWR _14848_/X sky130_fd_sc_hd__and3_4
X_17636_ _17077_/X _17097_/Y _17260_/X _17633_/Y _17635_/X VGND VGND VPWR VPWR _17636_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17567_ _17565_/Y _18081_/A VGND VGND VPWR VPWR _17567_/X sky130_fd_sc_hd__or2_4
X_14779_ _13966_/A _14779_/B VGND VGND VPWR VPWR _14781_/B sky130_fd_sc_hd__or2_4
XFILLER_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13171__A _15689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16518_ _16515_/X _16517_/Y VGND VGND VPWR VPWR _16518_/X sky130_fd_sc_hd__or2_4
X_19306_ _24140_/Q VGND VGND VPWR VPWR _19306_/Y sky130_fd_sc_hd__inv_2
X_17498_ _13059_/Y _17014_/X _17022_/X _17497_/X VGND VGND VPWR VPWR _17498_/X sky130_fd_sc_hd__o22a_4
XFILLER_17_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18920__A2 _18891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16449_ _11700_/X VGND VGND VPWR VPWR _16464_/A sky130_fd_sc_hd__buf_2
X_19237_ _19235_/A _19236_/A _19235_/Y _19236_/Y VGND VGND VPWR VPWR _19237_/X sky130_fd_sc_hd__o22a_4
X_19168_ _24304_/Q _19169_/A _19167_/Y VGND VGND VPWR VPWR _19168_/X sky130_fd_sc_hd__o21a_4
XFILLER_69_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18119_ _17874_/A _18118_/X VGND VGND VPWR VPWR _18119_/Y sky130_fd_sc_hd__nor2_4
X_19099_ _18965_/A _19097_/X _19098_/Y _19084_/X VGND VGND VPWR VPWR _19099_/X sky130_fd_sc_hd__o22a_4
XFILLER_69_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22480__A2 _22479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12515__A _13048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21130_ _21130_/A VGND VGND VPWR VPWR _21130_/X sky130_fd_sc_hd__buf_2
XANTENNA__20491__A1 _20229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21061_ _21112_/A _21348_/B _21162_/C _21784_/D VGND VGND VPWR VPWR _21061_/X sky130_fd_sc_hd__or4_4
XANTENNA__15826__A _12522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22232__A2 _22229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24144__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18202__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20012_ _19994_/X _17667_/A _20000_/X _20011_/X VGND VGND VPWR VPWR _20013_/A sky130_fd_sc_hd__o22a_4
XFILLER_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13346__A _15695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21991__B2 _21985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21563__A _21527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21963_ _21859_/X _21959_/X _15213_/B _21920_/X VGND VGND VPWR VPWR _23521_/D sky130_fd_sc_hd__o22a_4
XFILLER_67_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21743__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23702_ _23473_/CLK _23702_/D VGND VGND VPWR VPWR _12331_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_76_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20914_ _24195_/Q _20873_/X _20913_/X VGND VGND VPWR VPWR _20915_/A sky130_fd_sc_hd__o21a_4
XFILLER_82_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21894_ _21887_/A VGND VGND VPWR VPWR _21894_/X sky130_fd_sc_hd__buf_2
XFILLER_55_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23633_ _23122_/CLK _23633_/D VGND VGND VPWR VPWR _13190_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20849_/B _20650_/A VGND VGND VPWR VPWR _20845_/X sky130_fd_sc_hd__or2_4
XANTENNA__22299__A2 _22272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14177__A _14177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18872__A _18762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23170__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24296__CLK _24299_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23564_ _23564_/CLK _23564_/D VGND VGND VPWR VPWR _15471_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20776_ _20913_/A _20775_/X VGND VGND VPWR VPWR _20776_/X sky130_fd_sc_hd__or2_4
XANTENNA__22394__A _20338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18372__B1 _17259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22515_ _22068_/A _21582_/A _21297_/A _21213_/A VGND VGND VPWR VPWR _22516_/A sky130_fd_sc_hd__or4_4
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23495_ _23079_/CLK _23495_/D VGND VGND VPWR VPWR _23495_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16392__A _15948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14905__A _15146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22446_ _22446_/A VGND VGND VPWR VPWR _22446_/X sky130_fd_sc_hd__buf_2
XFILLER_6_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18675__A1 _18499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22377_ _22139_/X _22375_/X _14798_/B _22372_/X VGND VGND VPWR VPWR _23267_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12425__A _13550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12130_ _11748_/X _12128_/X _12129_/X VGND VGND VPWR VPWR _12130_/X sky130_fd_sc_hd__and3_4
X_24116_ _24203_/CLK _20081_/X HRESETn VGND VGND VPWR VPWR _16960_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_11_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21328_ _21261_/X _21326_/X _23885_/Q _21323_/X VGND VGND VPWR VPWR _23885_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21738__A _21737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12061_ _12051_/X _12061_/B _12061_/C VGND VGND VPWR VPWR _12061_/X sky130_fd_sc_hd__or3_4
X_21259_ _21247_/A VGND VGND VPWR VPWR _21259_/X sky130_fd_sc_hd__buf_2
X_24047_ _24047_/CLK _24047_/D VGND VGND VPWR VPWR _13466_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_81_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22223__A2 _22222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21431__B1 _15560_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15455__B _15455_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15820_ _15820_/A _15816_/X _15820_/C VGND VGND VPWR VPWR _15820_/X sky130_fd_sc_hd__or3_4
XANTENNA__13256__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21982__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17650__A2 _17544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12160__A _11717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22569__A _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15751_ _15751_/A _15686_/B VGND VGND VPWR VPWR _15751_/X sky130_fd_sc_hd__or2_4
X_12963_ _12963_/A _12963_/B _12963_/C VGND VGND VPWR VPWR _12963_/X sky130_fd_sc_hd__and3_4
XFILLER_45_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17670__B _17497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14702_ _14055_/A _14694_/X _14701_/X VGND VGND VPWR VPWR _14702_/X sky130_fd_sc_hd__and3_4
XANTENNA__15471__A _12585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11914_ _11913_/X VGND VGND VPWR VPWR _11915_/A sky130_fd_sc_hd__buf_2
X_18470_ _17874_/A _18271_/X VGND VGND VPWR VPWR _18470_/Y sky130_fd_sc_hd__nor2_4
X_15682_ _12693_/A _15747_/B VGND VGND VPWR VPWR _15684_/B sky130_fd_sc_hd__or2_4
X_12894_ _12462_/A _23891_/Q VGND VGND VPWR VPWR _12894_/X sky130_fd_sc_hd__or2_4
XFILLER_73_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17421_ _17421_/A VGND VGND VPWR VPWR _17422_/D sky130_fd_sc_hd__inv_2
X_14633_ _14603_/A _14631_/X _14632_/X VGND VGND VPWR VPWR _14633_/X sky130_fd_sc_hd__and3_4
XFILLER_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11845_ _15047_/A VGND VGND VPWR VPWR _13987_/A sky130_fd_sc_hd__buf_2
XFILLER_60_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18782__A _18782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17352_ _18395_/A VGND VGND VPWR VPWR _17382_/A sky130_fd_sc_hd__inv_2
X_14564_ _14563_/X VGND VGND VPWR VPWR _14564_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11776_ _11773_/X _11776_/B _11775_/X VGND VGND VPWR VPWR _11776_/X sky130_fd_sc_hd__and3_4
XANTENNA__17166__A1 _14565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16303_ _12837_/A VGND VGND VPWR VPWR _16303_/X sky130_fd_sc_hd__buf_2
X_13515_ _13559_/A _23279_/Q VGND VGND VPWR VPWR _13515_/X sky130_fd_sc_hd__or2_4
X_17283_ _14336_/X VGND VGND VPWR VPWR _17283_/Y sky130_fd_sc_hd__inv_2
X_14495_ _12383_/A _14431_/B VGND VGND VPWR VPWR _14495_/X sky130_fd_sc_hd__or2_4
XFILLER_105_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14815__A _14815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_36_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19022_ _18994_/X _19020_/X _19021_/Y _18999_/X VGND VGND VPWR VPWR _19022_/X sky130_fd_sc_hd__o22a_4
X_16234_ _16233_/X VGND VGND VPWR VPWR _16234_/Y sky130_fd_sc_hd__inv_2
X_13446_ _13442_/X _13443_/X _13446_/C VGND VGND VPWR VPWR _13452_/B sky130_fd_sc_hd__and3_4
X_16165_ _13397_/X VGND VGND VPWR VPWR _16202_/A sky130_fd_sc_hd__buf_2
XFILLER_86_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18666__A1 _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13377_ _13376_/X _13311_/B VGND VGND VPWR VPWR _13377_/X sky130_fd_sc_hd__or2_4
X_15116_ _14071_/A _15108_/X _15115_/X VGND VGND VPWR VPWR _15117_/C sky130_fd_sc_hd__and3_4
X_12328_ _12710_/A _12328_/B VGND VGND VPWR VPWR _12328_/X sky130_fd_sc_hd__or2_4
XANTENNA__21648__A _21662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16096_ _16096_/A _16096_/B VGND VGND VPWR VPWR _16098_/B sky130_fd_sc_hd__or2_4
XANTENNA__20552__A _20552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15047_ _15047_/A _15047_/B VGND VGND VPWR VPWR _15047_/X sky130_fd_sc_hd__and2_4
X_19924_ _20190_/A VGND VGND VPWR VPWR _22985_/A sky130_fd_sc_hd__buf_2
XANTENNA__15646__A _15645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12259_ _12728_/A _12259_/B VGND VGND VPWR VPWR _12259_/X sky130_fd_sc_hd__or2_4
XANTENNA__18022__A _18202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14550__A _13695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19855_ _19603_/A _19689_/A _19622_/A VGND VGND VPWR VPWR _19855_/X sky130_fd_sc_hd__o21a_4
XFILLER_116_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18806_ _14851_/X _18802_/X _20901_/A _18803_/X VGND VGND VPWR VPWR _24419_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13166__A _12315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19786_ _19718_/B VGND VGND VPWR VPWR _19786_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16998_ _16998_/A _16969_/B _16997_/X _18642_/A VGND VGND VPWR VPWR _16999_/C sky130_fd_sc_hd__or4_4
XFILLER_83_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19918__B2 _20490_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18737_ _18656_/A _17612_/X _17090_/X _18736_/X VGND VGND VPWR VPWR _18737_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15949_ _13437_/X VGND VGND VPWR VPWR _15959_/A sky130_fd_sc_hd__buf_2
XANTENNA__16477__A _16159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20528__A2 _20526_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21725__B2 _21723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22922__B1 _22924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18668_ _18668_/A VGND VGND VPWR VPWR _18668_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17944__A3 _17939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17619_ _17619_/A _17619_/B _17619_/C VGND VGND VPWR VPWR _18537_/B sky130_fd_sc_hd__or3_4
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_118_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR _23315_/CLK sky130_fd_sc_hd__clkbuf_1
X_18599_ _16919_/Y _18577_/Y _18594_/Y _17006_/A _18598_/X VGND VGND VPWR VPWR _18599_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_75_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20630_ _20630_/A _20630_/B VGND VGND VPWR VPWR _20630_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__20727__A HRDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20561_ _20561_/A VGND VGND VPWR VPWR _20561_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14725__A _14725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22300_ _11790_/B VGND VGND VPWR VPWR _23326_/D sky130_fd_sc_hd__buf_2
X_20492_ _20492_/A VGND VGND VPWR VPWR _20492_/X sky130_fd_sc_hd__buf_2
X_23280_ _24047_/CLK _23280_/D VGND VGND VPWR VPWR _13296_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24396__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22231_ _22115_/X _22229_/X _15824_/B _22226_/X VGND VGND VPWR VPWR _22231_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22453__A2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12245__A _12235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22162_ _22162_/A VGND VGND VPWR VPWR _22162_/X sky130_fd_sc_hd__buf_2
XFILLER_69_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21113_ _21113_/A VGND VGND VPWR VPWR _21118_/A sky130_fd_sc_hd__buf_2
XFILLER_47_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15556__A _15556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22093_ _20463_/A VGND VGND VPWR VPWR _22093_/X sky130_fd_sc_hd__buf_2
XFILLER_114_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14460__A _12269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21044_ _21015_/A VGND VGND VPWR VPWR _21044_/X sky130_fd_sc_hd__buf_2
XFILLER_99_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18867__A _12098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21964__B2 _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22995_ _22985_/X _17672_/A _22967_/X _22994_/X VGND VGND VPWR VPWR _22995_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16387__A _15999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15291__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13804__A _13647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21946_ _21828_/X _21945_/X _15670_/B _21942_/X VGND VGND VPWR VPWR _21946_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18593__B1 _17998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21192__A2 _21190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21877_ _21869_/X VGND VGND VPWR VPWR _21877_/X sky130_fd_sc_hd__buf_2
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _17069_/A VGND VGND VPWR VPWR _11631_/A sky130_fd_sc_hd__inv_2
X_23616_ _23073_/CLK _21781_/X VGND VGND VPWR VPWR _23616_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ _20622_/X _20827_/X _19211_/A _20736_/X VGND VGND VPWR VPWR _20828_/X sky130_fd_sc_hd__o22a_4
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _24432_/Q IRQ[17] _11560_/X VGND VGND VPWR VPWR _20086_/A sky130_fd_sc_hd__a21o_4
X_23547_ _24026_/CLK _23547_/D VGND VGND VPWR VPWR _23547_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18896__A1 _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20759_ _20517_/A VGND VGND VPWR VPWR _20759_/X sky130_fd_sc_hd__buf_2
XANTENNA__22692__A2 _22686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18107__A _18107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14635__A _15037_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13300_/A _23664_/Q VGND VGND VPWR VPWR _13300_/X sky130_fd_sc_hd__or2_4
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ _12320_/A _14278_/X _14279_/X VGND VGND VPWR VPWR _14280_/X sky130_fd_sc_hd__and3_4
XFILLER_6_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23478_ _23539_/CLK _22034_/X VGND VGND VPWR VPWR _12312_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13231_ _13231_/A _13231_/B _13231_/C VGND VGND VPWR VPWR _13235_/B sky130_fd_sc_hd__and3_4
X_22429_ _22427_/X _22428_/X _15652_/B _22423_/X VGND VGND VPWR VPWR _23246_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19845__B1 _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13162_ _12710_/A _13162_/B VGND VGND VPWR VPWR _13162_/X sky130_fd_sc_hd__or2_4
XANTENNA__20372__A _20372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24311__CLK _24299_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12113_ _16741_/A _12113_/B VGND VGND VPWR VPWR _12113_/X sky130_fd_sc_hd__and2_4
XANTENNA__11994__A _11994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15466__A _12585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13093_ _13082_/A _13086_/X _13092_/X VGND VGND VPWR VPWR _13093_/X sky130_fd_sc_hd__or3_4
X_17970_ _17818_/X _17828_/X _17813_/X _17816_/X VGND VGND VPWR VPWR _17971_/A sky130_fd_sc_hd__o22a_4
XFILLER_46_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12044_ _11995_/A VGND VGND VPWR VPWR _12044_/X sky130_fd_sc_hd__buf_2
X_16921_ _16919_/Y _17079_/A VGND VGND VPWR VPWR _16921_/X sky130_fd_sc_hd__or2_4
XFILLER_46_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21955__B2 _21949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19640_ _19637_/Y _19640_/B VGND VGND VPWR VPWR _19640_/X sky130_fd_sc_hd__and2_4
XFILLER_77_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17681__A _17681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16852_ _12996_/B _16899_/B _12996_/B _16899_/B VGND VGND VPWR VPWR _16876_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15803_ _12522_/A _15803_/B _15803_/C VGND VGND VPWR VPWR _15804_/C sky130_fd_sc_hd__and3_4
XFILLER_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16783_ _11823_/A _16783_/B _16782_/X VGND VGND VPWR VPWR _16783_/X sky130_fd_sc_hd__and3_4
X_19571_ _19566_/X VGND VGND VPWR VPWR _19659_/A sky130_fd_sc_hd__inv_2
X_13995_ _14841_/A _13995_/B VGND VGND VPWR VPWR _13995_/X sky130_fd_sc_hd__or2_4
XFILLER_20_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21707__A1 _21534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16297__A _15956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21707__B2 _21702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15734_ _15774_/A _15732_/X _15733_/X VGND VGND VPWR VPWR _15734_/X sky130_fd_sc_hd__and3_4
X_18522_ _18216_/A _18212_/Y VGND VGND VPWR VPWR _18522_/X sky130_fd_sc_hd__and2_4
XANTENNA__13714__A _13711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12946_ _12953_/A _23443_/Q VGND VGND VPWR VPWR _12946_/X sky130_fd_sc_hd__or2_4
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22380__B2 _22344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21931__A _21938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15665_ _15688_/A _15665_/B _15665_/C VGND VGND VPWR VPWR _15665_/X sky130_fd_sc_hd__or3_4
X_18453_ _18440_/X _18445_/Y _18447_/X _18451_/X _18452_/Y VGND VGND VPWR VPWR _18453_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_73_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12877_ _15392_/A VGND VGND VPWR VPWR _12878_/A sky130_fd_sc_hd__buf_2
X_14616_ _14727_/A _14614_/X _14615_/X VGND VGND VPWR VPWR _14616_/X sky130_fd_sc_hd__and3_4
X_17404_ _17042_/A _17404_/B VGND VGND VPWR VPWR _17404_/X sky130_fd_sc_hd__and2_4
X_11828_ _11758_/X VGND VGND VPWR VPWR _11829_/A sky130_fd_sc_hd__buf_2
X_18384_ _18383_/A _16976_/B VGND VGND VPWR VPWR _18384_/X sky130_fd_sc_hd__and2_4
X_15596_ _15604_/A _15592_/X _15596_/C VGND VGND VPWR VPWR _15597_/C sky130_fd_sc_hd__or3_4
XANTENNA__17139__A1 _14988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17321_/Y _17334_/X VGND VGND VPWR VPWR _17335_/X sky130_fd_sc_hd__or2_4
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14554_/A _14547_/B VGND VGND VPWR VPWR _14547_/X sky130_fd_sc_hd__or2_4
XANTENNA__18887__A1 _17164_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11759_ _11758_/X VGND VGND VPWR VPWR _11819_/A sky130_fd_sc_hd__buf_2
XFILLER_105_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14545__A _13754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17266_ _16678_/X VGND VGND VPWR VPWR _17266_/X sky130_fd_sc_hd__buf_2
X_14478_ _13054_/A _14476_/X _14477_/X VGND VGND VPWR VPWR _14482_/B sky130_fd_sc_hd__and3_4
X_16217_ _16193_/A _16217_/B VGND VGND VPWR VPWR _16217_/X sky130_fd_sc_hd__or2_4
X_19005_ _18994_/X _19003_/Y _19004_/Y _18999_/X VGND VGND VPWR VPWR _19005_/X sky130_fd_sc_hd__o22a_4
X_13429_ _13467_/A _13427_/X _13428_/X VGND VGND VPWR VPWR _13433_/B sky130_fd_sc_hd__and3_4
XANTENNA__18639__A1 _18697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17197_ _17130_/X _17193_/X _17163_/X _17196_/X VGND VGND VPWR VPWR _17197_/X sky130_fd_sc_hd__o22a_4
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12065__A _11994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20446__A1 _20229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16148_ _15937_/X VGND VGND VPWR VPWR _16151_/A sky130_fd_sc_hd__buf_2
XFILLER_118_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16079_ _16008_/Y _16077_/X VGND VGND VPWR VPWR _16080_/A sky130_fd_sc_hd__or2_4
XANTENNA__14280__A _12320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22199__B2 _22162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19907_ _19899_/X _24154_/Q _19903_/X _20342_/B VGND VGND VPWR VPWR _19907_/X sky130_fd_sc_hd__o22a_4
XFILLER_64_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15095__B _23807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21946__B2 _21942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19838_ _19573_/Y _19723_/B _19486_/Y VGND VGND VPWR VPWR _19839_/B sky130_fd_sc_hd__o21a_4
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19769_ HRDATA[0] VGND VGND VPWR VPWR _19769_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22002__A _22002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21800_ _21787_/X VGND VGND VPWR VPWR _21800_/X sky130_fd_sc_hd__buf_2
XFILLER_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22780_ _22777_/X _22779_/X VGND VGND VPWR VPWR _22781_/A sky130_fd_sc_hd__or2_4
XANTENNA__16000__A _15999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22371__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21174__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22937__A _22967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22371__B2 _22365_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21731_ _21576_/X _21726_/X _14872_/B _21687_/X VGND VGND VPWR VPWR _23648_/D sky130_fd_sc_hd__o22a_4
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24450_ _24203_/CLK _24450_/D HRESETn VGND VGND VPWR VPWR _24450_/Q sky130_fd_sc_hd__dfrtp_4
X_21662_ _21662_/A VGND VGND VPWR VPWR _21662_/X sky130_fd_sc_hd__buf_2
XFILLER_80_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22123__B2 _22120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23401_ _23910_/CLK _23401_/D VGND VGND VPWR VPWR _23401_/Q sky130_fd_sc_hd__dfxtp_4
X_20613_ _20511_/A VGND VGND VPWR VPWR _20613_/X sky130_fd_sc_hd__buf_2
XFILLER_51_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24363__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24381_ _24435_/CLK _24381_/D HRESETn VGND VGND VPWR VPWR _18930_/A sky130_fd_sc_hd__dfstp_4
X_21593_ _21510_/X _21591_/X _23740_/Q _21588_/X VGND VGND VPWR VPWR _23740_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14455__A _12450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22674__A2 _22672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20685__A1 _20622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23332_ _23812_/CLK _23332_/D VGND VGND VPWR VPWR _14652_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_71_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20544_ _20494_/X _20543_/X _24338_/Q _20453_/X VGND VGND VPWR VPWR _20544_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23089__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20685__B2 _20497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22672__A _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23263_ _23487_/CLK _23263_/D VGND VGND VPWR VPWR _23263_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17766__A _17766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22426__A2 _22416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20475_ _20475_/A VGND VGND VPWR VPWR _20475_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22214_ _22086_/X _22208_/X _16282_/B _22212_/X VGND VGND VPWR VPWR _23385_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23194_ _23130_/CLK _23194_/D VGND VGND VPWR VPWR _16387_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_105_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14902__B _23456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15286__A _14152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22145_ _22460_/A VGND VGND VPWR VPWR _22145_/X sky130_fd_sc_hd__buf_2
XANTENNA__12703__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22076_ _22125_/A VGND VGND VPWR VPWR _22101_/A sky130_fd_sc_hd__buf_2
XANTENNA__21937__B2 _21935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21027_ _21027_/A VGND VGND VPWR VPWR _21027_/X sky130_fd_sc_hd__buf_2
XFILLER_101_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12800_ _12800_/A _23988_/Q VGND VGND VPWR VPWR _12801_/C sky130_fd_sc_hd__or2_4
XFILLER_95_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13780_ _15399_/A _23335_/Q VGND VGND VPWR VPWR _13782_/B sky130_fd_sc_hd__or2_4
X_22978_ _22978_/A VGND VGND VPWR VPWR _23003_/A sky130_fd_sc_hd__buf_2
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18566__B1 _17782_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22362__B2 _22358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14349__B _14272_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12731_ _12705_/A _12728_/X _12730_/X VGND VGND VPWR VPWR _12732_/C sky130_fd_sc_hd__and3_4
X_21929_ _21799_/X _21924_/X _16401_/B _21928_/X VGND VGND VPWR VPWR _21929_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20912__A2 _20444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15450_ _15450_/A _15449_/X VGND VGND VPWR VPWR _15450_/X sky130_fd_sc_hd__and2_4
XFILLER_54_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12662_ _12954_/A _12662_/B _12662_/C VGND VGND VPWR VPWR _12662_/X sky130_fd_sc_hd__and3_4
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_101_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR _23770_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _15601_/A _14311_/B VGND VGND VPWR VPWR _14401_/X sky130_fd_sc_hd__or2_4
XANTENNA__22114__B2 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _15413_/A VGND VGND VPWR VPWR _13651_/A sky130_fd_sc_hd__buf_2
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11989__A _11936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15380_/Y VGND VGND VPWR VPWR _15381_/X sky130_fd_sc_hd__buf_2
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _13718_/A VGND VGND VPWR VPWR _12937_/A sky130_fd_sc_hd__buf_2
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14365__A _15643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ _17120_/A VGND VGND VPWR VPWR _17227_/A sky130_fd_sc_hd__buf_2
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _15578_/A _14332_/B _14331_/X VGND VGND VPWR VPWR _14332_/X sky130_fd_sc_hd__and3_4
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ _24438_/Q IRQ[23] _20160_/A VGND VGND VPWR VPWR _11544_/X sky130_fd_sc_hd__a21o_4
XANTENNA_clkbuf_5_21_0_HCLK_A clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17051_ _17054_/A _16916_/A _16909_/B _11632_/X VGND VGND VPWR VPWR _17051_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _14263_/A VGND VGND VPWR VPWR _14263_/X sky130_fd_sc_hd__buf_2
XFILLER_51_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22417__A2 _22416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16002_ _16002_/A _23864_/Q VGND VGND VPWR VPWR _16002_/X sky130_fd_sc_hd__or2_4
XFILLER_109_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13214_ _13214_/A _13214_/B _13214_/C VGND VGND VPWR VPWR _13214_/X sky130_fd_sc_hd__and3_4
X_14194_ _14182_/A _23753_/Q VGND VGND VPWR VPWR _14195_/C sky130_fd_sc_hd__or2_4
XANTENNA__15196__A _15201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13145_ _12240_/X _13145_/B VGND VGND VPWR VPWR _13145_/X sky130_fd_sc_hd__or2_4
XANTENNA__12613__A _12613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13076_ _13128_/A _13074_/X _13075_/X VGND VGND VPWR VPWR _13082_/B sky130_fd_sc_hd__and3_4
X_17953_ _17895_/Y _17951_/X _17896_/A _17952_/X VGND VGND VPWR VPWR _17953_/X sky130_fd_sc_hd__o22a_4
XFILLER_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12027_ _11853_/X _12027_/B VGND VGND VPWR VPWR _12027_/X sky130_fd_sc_hd__and2_4
X_16904_ _16903_/X VGND VGND VPWR VPWR _16904_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22050__B1 _23467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17884_ _17767_/X _17883_/X _17767_/X _17883_/X VGND VGND VPWR VPWR _17884_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20600__A1 _20468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19623_ _19600_/X _19808_/A _19622_/Y _19822_/A VGND VGND VPWR VPWR _19623_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20600__B2 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16835_ _15391_/X _15919_/Y VGND VGND VPWR VPWR _16835_/X sky130_fd_sc_hd__and2_4
XFILLER_4_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13444__A _12520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19554_ _19793_/A VGND VGND VPWR VPWR _19554_/X sky130_fd_sc_hd__buf_2
X_13978_ _12196_/A _13978_/B _13977_/X VGND VGND VPWR VPWR _13978_/X sky130_fd_sc_hd__and3_4
X_16766_ _12152_/A VGND VGND VPWR VPWR _16803_/A sky130_fd_sc_hd__buf_2
XFILLER_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21156__A2 _21154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22353__B2 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18505_ _18505_/A VGND VGND VPWR VPWR _18505_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12929_ _12640_/A _12929_/B VGND VGND VPWR VPWR _12929_/X sky130_fd_sc_hd__or2_4
X_15717_ _15724_/A _15655_/B VGND VGND VPWR VPWR _15719_/B sky130_fd_sc_hd__or2_4
XANTENNA__13163__B _23569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16697_ _12083_/A _23675_/Q VGND VGND VPWR VPWR _16697_/X sky130_fd_sc_hd__or2_4
X_19485_ _19485_/A _19872_/B VGND VGND VPWR VPWR _19691_/A sky130_fd_sc_hd__or2_4
XFILLER_94_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18436_ _18344_/X _18351_/B VGND VGND VPWR VPWR _18436_/Y sky130_fd_sc_hd__nand2_4
X_15648_ _15649_/B VGND VGND VPWR VPWR _15648_/X sky130_fd_sc_hd__buf_2
XANTENNA__16474__B _16398_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11899__A _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15579_ _15398_/A _15575_/X _15579_/C VGND VGND VPWR VPWR _15579_/X sky130_fd_sc_hd__or3_4
X_18367_ _18367_/A VGND VGND VPWR VPWR _18367_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22656__A2 _22650_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14275__A _12257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17318_ _18656_/B VGND VGND VPWR VPWR _18655_/B sky130_fd_sc_hd__inv_2
X_18298_ _18244_/A _18298_/B _18298_/C _18298_/D VGND VGND VPWR VPWR _18298_/X sky130_fd_sc_hd__or4_4
XANTENNA__12507__B _12620_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17249_ _17249_/A _17817_/A VGND VGND VPWR VPWR _17249_/X sky130_fd_sc_hd__or2_4
X_20260_ _20449_/A VGND VGND VPWR VPWR _20260_/X sky130_fd_sc_hd__buf_2
XFILLER_116_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18088__A2 _18061_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15818__B _15818_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13619__A _12883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20191_ _22017_/A _22017_/B VGND VGND VPWR VPWR _21212_/A sky130_fd_sc_hd__or2_4
XANTENNA__21092__B2 _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12523__A _13019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21836__A _21812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23950_ _24044_/CLK _23950_/D VGND VGND VPWR VPWR _15748_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_44_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15834__A _12914_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21395__A2 _21390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22901_ _18610_/A _18701_/X _18607_/X VGND VGND VPWR VPWR _22901_/X sky130_fd_sc_hd__o21a_4
XFILLER_69_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22592__B2 _22590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15553__B _23947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23881_ _23561_/CLK _23881_/D VGND VGND VPWR VPWR _23881_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16271__A1 _11852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13354__A _12803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22832_ _15120_/Y _22826_/X _22827_/X VGND VGND VPWR VPWR _22832_/X sky130_fd_sc_hd__o21a_4
XFILLER_99_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19373__A2_N _18061_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22667__A _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22763_ _22763_/A _22763_/B VGND VGND VPWR VPWR _22763_/Y sky130_fd_sc_hd__nand2_4
XFILLER_112_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16665__A _16630_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21714_ _21546_/X _21712_/X _15798_/B _21709_/X VGND VGND VPWR VPWR _21714_/X sky130_fd_sc_hd__o22a_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22694_ _21543_/A _22693_/X _15762_/B _22690_/X VGND VGND VPWR VPWR _22694_/X sky130_fd_sc_hd__o22a_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24433_ _23326_/CLK _18786_/X HRESETn VGND VGND VPWR VPWR _20558_/A sky130_fd_sc_hd__dfrtp_4
X_21645_ _21637_/X VGND VGND VPWR VPWR _21645_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19976__A _20000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11602__A _11599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20658__B2 _20473_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24364_ _24365_/CLK _24364_/D HRESETn VGND VGND VPWR VPWR _24364_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_16_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21576_ _21291_/A VGND VGND VPWR VPWR _21576_/X sky130_fd_sc_hd__buf_2
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18720__B1 _18048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20915__A _20915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23315_ _23315_/CLK _23315_/D VGND VGND VPWR VPWR _22311_/A sky130_fd_sc_hd__dfxtp_4
X_20527_ _20242_/X VGND VGND VPWR VPWR _20527_/X sky130_fd_sc_hd__buf_2
X_24295_ _24299_/CLK _24295_/D HRESETn VGND VGND VPWR VPWR _24295_/Q sky130_fd_sc_hd__dfrtp_4
X_23246_ _23564_/CLK _23246_/D VGND VGND VPWR VPWR _15652_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20458_ _24246_/Q VGND VGND VPWR VPWR _20458_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23874__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21083__A1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13529__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21083__B2 _21079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23177_ _23978_/CLK _22551_/X VGND VGND VPWR VPWR _23177_/Q sky130_fd_sc_hd__dfxtp_4
X_20389_ _20376_/X _20377_/X _20288_/X _20388_/Y VGND VGND VPWR VPWR _20389_/X sky130_fd_sc_hd__a211o_4
XFILLER_97_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22128_ _22127_/X _22125_/X _13729_/B _22120_/X VGND VGND VPWR VPWR _22128_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20650__A _20650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12152__B _23901_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_26_0_HCLK clkbuf_6_13_0_HCLK/X VGND VGND VPWR VPWR _23145_/CLK sky130_fd_sc_hd__clkbuf_1
X_14950_ _15074_/A _23520_/Q VGND VGND VPWR VPWR _14951_/C sky130_fd_sc_hd__or2_4
XANTENNA__15744__A _11680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22059_ _22052_/A VGND VGND VPWR VPWR _22059_/X sky130_fd_sc_hd__buf_2
XFILLER_102_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_89_0_HCLK clkbuf_6_44_0_HCLK/X VGND VGND VPWR VPWR _24092_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21386__A2 _21383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18787__B1 _24432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13901_ _13901_/A _13893_/X _13900_/X VGND VGND VPWR VPWR _13901_/X sky130_fd_sc_hd__and3_4
X_14881_ _12250_/A _14881_/B _14880_/X VGND VGND VPWR VPWR _14885_/B sky130_fd_sc_hd__and3_4
XFILLER_97_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15463__B _15463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13264__A _13257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13832_ _13635_/A _13906_/B VGND VGND VPWR VPWR _13832_/X sky130_fd_sc_hd__or2_4
X_16620_ _16651_/A _16620_/B VGND VGND VPWR VPWR _16621_/C sky130_fd_sc_hd__or2_4
XFILLER_1_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18539__B1 _18398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21138__A2 _21133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16551_ _11903_/A VGND VGND VPWR VPWR _16583_/A sky130_fd_sc_hd__buf_2
XANTENNA__21481__A _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13763_ _12935_/A _23464_/Q VGND VGND VPWR VPWR _13765_/B sky130_fd_sc_hd__or2_4
XFILLER_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12714_ _15812_/A _12713_/X VGND VGND VPWR VPWR _12714_/X sky130_fd_sc_hd__and2_4
X_15502_ _15497_/A _23788_/Q VGND VGND VPWR VPWR _15503_/C sky130_fd_sc_hd__or2_4
XFILLER_91_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16482_ _16464_/A _16413_/B VGND VGND VPWR VPWR _16482_/X sky130_fd_sc_hd__or2_4
X_19270_ _19218_/A _19218_/B _19269_/Y VGND VGND VPWR VPWR _24269_/D sky130_fd_sc_hd__o21a_4
XFILLER_95_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13694_ _13694_/A VGND VGND VPWR VPWR _13890_/A sky130_fd_sc_hd__buf_2
X_15433_ _12211_/A _23404_/Q VGND VGND VPWR VPWR _15433_/X sky130_fd_sc_hd__or2_4
X_18221_ _17456_/Y _18219_/X _18160_/X VGND VGND VPWR VPWR _18221_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__22099__B1 _12711_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12645_ _12964_/A _12641_/X _12645_/C VGND VGND VPWR VPWR _12656_/B sky130_fd_sc_hd__or3_4
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22638__A2 _22636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12608__A _12963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ _15333_/A _15304_/B VGND VGND VPWR VPWR _15365_/C sky130_fd_sc_hd__or2_4
X_18152_ _18152_/A _18151_/X VGND VGND VPWR VPWR _18152_/X sky130_fd_sc_hd__or2_4
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12576_ _13700_/A VGND VGND VPWR VPWR _12638_/A sky130_fd_sc_hd__buf_2
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21310__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14315_ _14315_/A VGND VGND VPWR VPWR _15576_/A sky130_fd_sc_hd__buf_2
X_17103_ _18713_/A VGND VGND VPWR VPWR _17103_/X sky130_fd_sc_hd__buf_2
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _11527_/A _11526_/X VGND VGND VPWR VPWR _11527_/X sky130_fd_sc_hd__or2_4
X_18083_ _18083_/A VGND VGND VPWR VPWR _18083_/Y sky130_fd_sc_hd__inv_2
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15295_ _12531_/A _15291_/X _15294_/X VGND VGND VPWR VPWR _15295_/X sky130_fd_sc_hd__or3_4
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17034_ _17105_/A VGND VGND VPWR VPWR _17034_/Y sky130_fd_sc_hd__inv_2
X_14246_ _14246_/A _14244_/X _14246_/C VGND VGND VPWR VPWR _14250_/B sky130_fd_sc_hd__and3_4
XANTENNA__13439__A _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21074__B2 _21072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14177_ _14177_/A VGND VGND VPWR VPWR _14183_/A sky130_fd_sc_hd__buf_2
XFILLER_113_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13128_ _13128_/A _13126_/X _13128_/C VGND VGND VPWR VPWR _13132_/B sky130_fd_sc_hd__and3_4
X_18985_ _24373_/Q VGND VGND VPWR VPWR _18985_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15654__A _15654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13059_ _13059_/A VGND VGND VPWR VPWR _13059_/Y sky130_fd_sc_hd__inv_2
X_17936_ _17798_/X _17935_/X _17866_/X VGND VGND VPWR VPWR _17936_/X sky130_fd_sc_hd__o21a_4
XFILLER_39_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18030__A _18137_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21377__A2 _21376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22574__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17867_ _17864_/X _17865_/X _17866_/X VGND VGND VPWR VPWR _17867_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18965__A _18965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19606_ _19624_/A _19605_/X VGND VGND VPWR VPWR _19606_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13174__A _12728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16818_ _16682_/A _16815_/Y _16681_/A VGND VGND VPWR VPWR _16898_/A sky130_fd_sc_hd__o21ai_4
XFILLER_113_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17798_ _17797_/X VGND VGND VPWR VPWR _17798_/X sky130_fd_sc_hd__buf_2
X_19537_ _19537_/A _19537_/B VGND VGND VPWR VPWR _19537_/Y sky130_fd_sc_hd__nand2_4
X_16749_ _16772_/A _16749_/B VGND VGND VPWR VPWR _16752_/B sky130_fd_sc_hd__or2_4
XFILLER_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13902__A _13890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19468_ _19464_/Y _19523_/A VGND VGND VPWR VPWR _19468_/X sky130_fd_sc_hd__or2_4
XFILLER_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18419_ _18295_/A _17377_/B VGND VGND VPWR VPWR _18419_/Y sky130_fd_sc_hd__nor2_4
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14567__A1 _14493_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19399_ _19385_/A VGND VGND VPWR VPWR _19399_/X sky130_fd_sc_hd__buf_2
XANTENNA__12518__A _12518_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21430_ _21416_/A VGND VGND VPWR VPWR _21430_/X sky130_fd_sc_hd__buf_2
XANTENNA__21837__B1 _23595_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17505__A1 _16624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21361_ _21232_/X _21355_/X _16297_/B _21359_/X VGND VGND VPWR VPWR _23865_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15829__A _12477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18205__A _18205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23100_ _23100_/CLK _23100_/D VGND VGND VPWR VPWR _23100_/Q sky130_fd_sc_hd__dfxtp_4
X_20312_ _20484_/A _20312_/B VGND VGND VPWR VPWR _20312_/X sky130_fd_sc_hd__or2_4
X_24080_ _23157_/CLK _24080_/D VGND VGND VPWR VPWR _24080_/Q sky130_fd_sc_hd__dfxtp_4
X_21292_ _21291_/X _21283_/X _14879_/B _21230_/A VGND VGND VPWR VPWR _21292_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23031_ _23031_/A VGND VGND VPWR VPWR HADDR[25] sky130_fd_sc_hd__inv_2
X_20243_ _20242_/X VGND VGND VPWR VPWR _20500_/A sky130_fd_sc_hd__buf_2
XFILLER_104_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12253__A _15448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20812__A1 _18570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20174_ _20077_/D _20173_/X VGND VGND VPWR VPWR _20174_/X sky130_fd_sc_hd__or2_4
XFILLER_27_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15564__A _11911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22014__B1 _14857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21368__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23277__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23933_ _23931_/CLK _23933_/D VGND VGND VPWR VPWR _23933_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18875__A _18891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23864_ _24088_/CLK _23864_/D VGND VGND VPWR VPWR _23864_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13058__A1 _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22815_ _22821_/A _17298_/Y VGND VGND VPWR VPWR _22815_/X sky130_fd_sc_hd__or2_4
X_23795_ _23859_/CLK _21471_/X VGND VGND VPWR VPWR _12974_/B sky130_fd_sc_hd__dfxtp_4
X_22746_ _22737_/X _22746_/B _22746_/C _22746_/D VGND VGND VPWR VPWR _22746_/X sky130_fd_sc_hd__or4_4
XFILLER_77_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21540__A2 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22677_ _21799_/A _22672_/X _16434_/B _22676_/X VGND VGND VPWR VPWR _23098_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12428__A _12672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12430_ _12429_/X VGND VGND VPWR VPWR _12430_/X sky130_fd_sc_hd__buf_2
X_24416_ _24425_/CLK _24416_/D HRESETn VGND VGND VPWR VPWR _20966_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21628_ _21570_/X _21626_/X _14791_/B _21623_/X VGND VGND VPWR VPWR _23715_/D sky130_fd_sc_hd__o22a_4
XFILLER_103_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12361_ _12381_/A _12241_/B VGND VGND VPWR VPWR _12361_/X sky130_fd_sc_hd__or2_4
X_24347_ _24344_/CLK _24347_/D HRESETn VGND VGND VPWR VPWR _11532_/A sky130_fd_sc_hd__dfstp_4
XFILLER_16_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21559_ _21558_/X _21556_/X _13713_/B _21551_/X VGND VGND VPWR VPWR _23752_/D sky130_fd_sc_hd__o22a_4
X_14100_ _14991_/A VGND VGND VPWR VPWR _14108_/A sky130_fd_sc_hd__buf_2
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15080_ _15104_/A _15080_/B _15079_/X VGND VGND VPWR VPWR _15080_/X sky130_fd_sc_hd__and3_4
XFILLER_10_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12292_ _15688_/A _12292_/B _12291_/X VGND VGND VPWR VPWR _12292_/X sky130_fd_sc_hd__or3_4
X_24278_ _24435_/CLK _19252_/X HRESETn VGND VGND VPWR VPWR _24278_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15458__B _15458_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14362__B _14279_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14031_ _14031_/A _23658_/Q VGND VGND VPWR VPWR _14033_/B sky130_fd_sc_hd__or2_4
X_23229_ _24092_/CLK _22473_/X VGND VGND VPWR VPWR _12177_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17954__A _18062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13259__A _13211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21056__B2 _21012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19872__C _19872_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18770_ _12184_/X _18765_/X _20297_/A _18768_/X VGND VGND VPWR VPWR _24445_/D sky130_fd_sc_hd__o22a_4
X_15982_ _15957_/A _23832_/Q VGND VGND VPWR VPWR _15983_/C sky130_fd_sc_hd__or2_4
XFILLER_118_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22556__B2 _22554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16289__B _16289_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17721_ _17723_/B _17720_/X VGND VGND VPWR VPWR _17721_/X sky130_fd_sc_hd__or2_4
XFILLER_23_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14933_ _15063_/A _14930_/X _14932_/X VGND VGND VPWR VPWR _14934_/C sky130_fd_sc_hd__and3_4
XFILLER_94_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20031__A2 _17893_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17652_ _17652_/A _17652_/B VGND VGND VPWR VPWR _17659_/A sky130_fd_sc_hd__and2_4
XFILLER_36_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14864_ _13984_/A _14864_/B VGND VGND VPWR VPWR _14864_/X sky130_fd_sc_hd__or2_4
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17983__B2 _17982_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16603_ _12153_/A VGND VGND VPWR VPWR _16800_/A sky130_fd_sc_hd__buf_2
X_13815_ _13623_/A _13815_/B VGND VGND VPWR VPWR _13815_/X sky130_fd_sc_hd__or2_4
X_14795_ _13851_/A _14733_/B VGND VGND VPWR VPWR _14795_/X sky130_fd_sc_hd__or2_4
X_17583_ _17559_/A _17567_/X VGND VGND VPWR VPWR _17583_/X sky130_fd_sc_hd__or2_4
XFILLER_21_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14818__A _14039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22100__A _22100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19322_ _19318_/X _18090_/X _19321_/X _20414_/A VGND VGND VPWR VPWR _24248_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13722__A _13770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20539__B _20539_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13746_ _12646_/A _13746_/B _13746_/C VGND VGND VPWR VPWR _13747_/C sky130_fd_sc_hd__and3_4
X_16534_ _11936_/X VGND VGND VPWR VPWR _16542_/A sky130_fd_sc_hd__buf_2
XFILLER_1_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19253_ _19226_/X VGND VGND VPWR VPWR _19253_/Y sky130_fd_sc_hd__inv_2
X_13677_ _13677_/A _13675_/X _13676_/X VGND VGND VPWR VPWR _13681_/B sky130_fd_sc_hd__and3_4
X_16465_ _16465_/A _16405_/B VGND VGND VPWR VPWR _16466_/C sky130_fd_sc_hd__or2_4
XFILLER_108_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18204_ _18204_/A _17455_/X VGND VGND VPWR VPWR _18204_/X sky130_fd_sc_hd__or2_4
X_12628_ _12643_/A _12628_/B VGND VGND VPWR VPWR _12629_/C sky130_fd_sc_hd__or2_4
X_15416_ _15443_/A _15473_/B VGND VGND VPWR VPWR _15418_/B sky130_fd_sc_hd__or2_4
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16396_ _16400_/A _16472_/B VGND VGND VPWR VPWR _16396_/X sky130_fd_sc_hd__or2_4
X_19184_ _24296_/Q _19117_/B _19183_/Y VGND VGND VPWR VPWR _24296_/D sky130_fd_sc_hd__o21a_4
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15347_ _11661_/A _15347_/B _15346_/X VGND VGND VPWR VPWR _15347_/X sky130_fd_sc_hd__or3_4
X_18135_ _18205_/A _17523_/Y VGND VGND VPWR VPWR _18135_/X sky130_fd_sc_hd__and2_4
XANTENNA__15649__A _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12559_ _11842_/X _11618_/X _12517_/X _11596_/X _12558_/X VGND VGND VPWR VPWR _12559_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22492__B1 _13568_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14553__A _13754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15278_ _14603_/A _15276_/X _15277_/X VGND VGND VPWR VPWR _15278_/X sky130_fd_sc_hd__and3_4
X_18066_ _18066_/A _18066_/B VGND VGND VPWR VPWR _18067_/D sky130_fd_sc_hd__and2_4
XFILLER_7_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14272__B _14272_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14229_ _14204_/A _23593_/Q VGND VGND VPWR VPWR _14232_/B sky130_fd_sc_hd__or2_4
X_17017_ _17010_/A VGND VGND VPWR VPWR _17018_/A sky130_fd_sc_hd__inv_2
XANTENNA__13169__A _15812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21047__B2 _21041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22244__B1 _14698_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12073__A _12096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18968_ _18999_/A VGND VGND VPWR VPWR _18968_/X sky130_fd_sc_hd__buf_2
XANTENNA__12801__A _12754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17919_ _17911_/X _17214_/X _17912_/X _17204_/X VGND VGND VPWR VPWR _17919_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_39_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18899_ _18877_/A VGND VGND VPWR VPWR _18899_/X sky130_fd_sc_hd__buf_2
XANTENNA__19412__B2 _24192_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_72_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR _23293_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20022__A2 _17674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20930_ _20825_/X _20930_/B VGND VGND VPWR VPWR _20930_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19963__A2 _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21770__A2 _21769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20861_ _20759_/X _20860_/X _19114_/A _20769_/X VGND VGND VPWR VPWR _20862_/B sky130_fd_sc_hd__o22a_4
XANTENNA__15831__B _15831_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14728__A _14158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22600_ _22600_/A VGND VGND VPWR VPWR _22600_/X sky130_fd_sc_hd__buf_2
XANTENNA__13632__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23580_ _23485_/CLK _23580_/D VGND VGND VPWR VPWR _23580_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20792_ _20792_/A VGND VGND VPWR VPWR _20792_/Y sky130_fd_sc_hd__inv_2
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22945__A _18506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22531_ _22406_/X _22529_/X _16096_/B _22526_/X VGND VGND VPWR VPWR _22531_/X sky130_fd_sc_hd__o22a_4
XFILLER_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12248__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22462_ _21001_/A VGND VGND VPWR VPWR _22462_/X sky130_fd_sc_hd__buf_2
XFILLER_33_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24201_ _24473_/CLK _19400_/X HRESETn VGND VGND VPWR VPWR _24201_/Q sky130_fd_sc_hd__dfrtp_4
X_21413_ _21234_/X _21412_/X _23832_/Q _21409_/X VGND VGND VPWR VPWR _23832_/D sky130_fd_sc_hd__o22a_4
XFILLER_13_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15559__A _14283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21286__B2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22393_ _22390_/X _22392_/X _12118_/B _22387_/X VGND VGND VPWR VPWR _23261_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14463__A _14463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24132_ _24241_/CLK _19999_/Y HRESETn VGND VGND VPWR VPWR _24132_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21344_ _21289_/X _21340_/X _23873_/Q _21301_/X VGND VGND VPWR VPWR _21344_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24063_ _23313_/CLK _24063_/D VGND VGND VPWR VPWR _24063_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21038__B2 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21275_ _20819_/A VGND VGND VPWR VPWR _21275_/X sky130_fd_sc_hd__buf_2
XFILLER_11_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19100__B1 _18971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23014_ _22985_/A VGND VGND VPWR VPWR _23014_/X sky130_fd_sc_hd__buf_2
X_20226_ _20226_/A _20226_/B VGND VGND VPWR VPWR _20226_/X sky130_fd_sc_hd__or2_4
XANTENNA__19651__A1 _19554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13807__A _13614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20261__A2 _18814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20157_ _24434_/Q IRQ[19] _20156_/X VGND VGND VPWR VPWR _20157_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__13279__A1 _13202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12711__A _12711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23912__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22538__B2 _22533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20549__B1 _20548_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20088_ _20071_/B VGND VGND VPWR VPWR _20089_/C sky130_fd_sc_hd__inv_2
XFILLER_58_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17414__B1 _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11930_ _13813_/A VGND VGND VPWR VPWR _13025_/A sky130_fd_sc_hd__buf_2
XFILLER_85_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21210__B2 _21165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19954__A2 _19364_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23916_ _23698_/CLK _23916_/D VGND VGND VPWR VPWR _23916_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21761__A2 _21755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11861_ _12458_/A VGND VGND VPWR VPWR _11861_/X sky130_fd_sc_hd__buf_2
X_23847_ _23847_/CLK _21386_/X VGND VGND VPWR VPWR _13906_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14638__A _14172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13600_ _13600_/A VGND VGND VPWR VPWR _15435_/A sky130_fd_sc_hd__buf_2
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14580_ _14575_/X _14662_/B VGND VGND VPWR VPWR _14581_/C sky130_fd_sc_hd__or2_4
X_11792_ _11823_/A _11790_/X _11791_/X VGND VGND VPWR VPWR _11792_/X sky130_fd_sc_hd__and3_4
X_23778_ _23907_/CLK _23778_/D VGND VGND VPWR VPWR _15304_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21513__A2 _21508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13531_ _13559_/A _13531_/B VGND VGND VPWR VPWR _13532_/C sky130_fd_sc_hd__or2_4
XANTENNA__22710__B2 _22704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22729_ _22728_/Y _22772_/A _22728_/Y _22772_/A VGND VGND VPWR VPWR _22747_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13261__B _24081_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12158__A _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16250_ _16151_/A _16248_/X _16249_/X VGND VGND VPWR VPWR _16250_/X sky130_fd_sc_hd__and3_4
X_13462_ _13427_/A _23887_/Q VGND VGND VPWR VPWR _13462_/X sky130_fd_sc_hd__or2_4
XFILLER_16_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15201_ _15201_/A _15146_/B VGND VGND VPWR VPWR _15201_/X sky130_fd_sc_hd__or2_4
X_12413_ _12596_/A VGND VGND VPWR VPWR _12413_/X sky130_fd_sc_hd__buf_2
XANTENNA__11997__A _11997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16181_ _16201_/A _16181_/B VGND VGND VPWR VPWR _16183_/B sky130_fd_sc_hd__or2_4
XANTENNA__15469__A _13770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13393_ _13354_/X _23952_/Q VGND VGND VPWR VPWR _13394_/C sky130_fd_sc_hd__or2_4
XFILLER_51_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15132_ _14083_/A _15132_/B VGND VGND VPWR VPWR _15132_/X sky130_fd_sc_hd__or2_4
X_12344_ _12826_/A _12206_/B VGND VGND VPWR VPWR _12344_/X sky130_fd_sc_hd__or2_4
XFILLER_86_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22590__A _22583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23442__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15063_ _15063_/A VGND VGND VPWR VPWR _15104_/A sky130_fd_sc_hd__buf_2
X_19940_ _18062_/A _18744_/X VGND VGND VPWR VPWR _19940_/X sky130_fd_sc_hd__or2_4
XANTENNA__21029__B2 _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12275_ _12238_/X VGND VGND VPWR VPWR _12711_/A sky130_fd_sc_hd__buf_2
X_14014_ _14021_/A _24010_/Q VGND VGND VPWR VPWR _14017_/B sky130_fd_sc_hd__or2_4
XFILLER_107_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19871_ _19730_/A _19730_/D _19742_/B VGND VGND VPWR VPWR _19881_/B sky130_fd_sc_hd__o21ai_4
XFILLER_49_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18822_ _11837_/X _18818_/X _24414_/Q _18821_/X VGND VGND VPWR VPWR _24414_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12621__A _12605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18753_ _17006_/A _18752_/X _17737_/A _16935_/X VGND VGND VPWR VPWR _18753_/X sky130_fd_sc_hd__o22a_4
X_15965_ _15956_/A _23576_/Q VGND VGND VPWR VPWR _15965_/X sky130_fd_sc_hd__or2_4
XFILLER_49_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17704_ _16956_/A _17404_/X VGND VGND VPWR VPWR _17704_/X sky130_fd_sc_hd__and2_4
XFILLER_114_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17405__B1 _17013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15932__A _11884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_59_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14916_ _15047_/A _14916_/B VGND VGND VPWR VPWR _14916_/X sky130_fd_sc_hd__and2_4
X_18684_ _17741_/X VGND VGND VPWR VPWR _18684_/Y sky130_fd_sc_hd__inv_2
X_15896_ _13500_/X _15894_/X _15895_/X VGND VGND VPWR VPWR _15897_/C sky130_fd_sc_hd__and3_4
X_17635_ _17077_/A _17633_/B _17634_/X VGND VGND VPWR VPWR _17635_/X sky130_fd_sc_hd__o21a_4
X_14847_ _14847_/A _14843_/X _14846_/X VGND VGND VPWR VPWR _14848_/C sky130_fd_sc_hd__or3_4
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13452__A _11861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17566_ _16235_/X _17564_/B VGND VGND VPWR VPWR _18081_/A sky130_fd_sc_hd__and2_4
X_14778_ _14778_/A _14778_/B _14778_/C VGND VGND VPWR VPWR _14778_/X sky130_fd_sc_hd__and3_4
XFILLER_56_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19305_ _19304_/X VGND VGND VPWR VPWR _19305_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22701__B2 _22697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16517_ _16516_/X VGND VGND VPWR VPWR _16517_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13729_ _15497_/A _13729_/B VGND VGND VPWR VPWR _13729_/X sky130_fd_sc_hd__or2_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17497_ _17506_/A _17497_/B VGND VGND VPWR VPWR _17497_/X sky130_fd_sc_hd__or2_4
XFILLER_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12068__A _11966_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19236_ _19236_/A VGND VGND VPWR VPWR _19236_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16448_ _12830_/A VGND VGND VPWR VPWR _16506_/A sky130_fd_sc_hd__buf_2
XFILLER_20_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15379__A _11652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19167_ _19167_/A VGND VGND VPWR VPWR _19167_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16379_ _16302_/X _16376_/X _16378_/Y VGND VGND VPWR VPWR _16519_/A sky130_fd_sc_hd__a21o_4
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14283__A _14283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18118_ _18040_/X _18117_/X _17868_/A VGND VGND VPWR VPWR _18118_/X sky130_fd_sc_hd__o21a_4
X_19098_ _19098_/A VGND VGND VPWR VPWR _19098_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22217__B1 _16211_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18049_ _18047_/A _18046_/X _18048_/X VGND VGND VPWR VPWR _18049_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_99_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21060_ _21060_/A VGND VGND VPWR VPWR _21784_/D sky130_fd_sc_hd__buf_2
XFILLER_67_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20011_ _18259_/X _20009_/X _20010_/Y _19996_/X VGND VGND VPWR VPWR _20011_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13627__A _13794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12531__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16003__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21991__A2 _21988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15842__A _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21962_ _21857_/X _21959_/X _15343_/B _21956_/X VGND VGND VPWR VPWR _23522_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23701_ _24021_/CLK _21653_/X VGND VGND VPWR VPWR _12660_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_66_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21743__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20913_ _20913_/A _20912_/X VGND VGND VPWR VPWR _20913_/X sky130_fd_sc_hd__or2_4
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21893_ _21826_/X _21887_/X _13521_/B _21891_/X VGND VGND VPWR VPWR _21893_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14458__A _15404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23632_ _23632_/CLK _23632_/D VGND VGND VPWR VPWR _13337_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ _20844_/A _20844_/B VGND VGND VPWR VPWR _20844_/X sky130_fd_sc_hd__or2_4
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_2_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR _24126_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23563_ _23915_/CLK _23563_/D VGND VGND VPWR VPWR _23563_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17769__A _17769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20775_ _24233_/Q _20639_/X _20774_/X VGND VGND VPWR VPWR _20775_/X sky130_fd_sc_hd__o21a_4
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18372__A1 _17792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18372__B2 _18153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22514_ _11749_/B VGND VGND VPWR VPWR _22514_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23494_ _23494_/CLK _23494_/D VGND VGND VPWR VPWR _14269_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20195__A _16929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22445_ _22444_/X _22440_/X _13841_/B _22435_/X VGND VGND VPWR VPWR _22445_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15289__A _14149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12706__A _12706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22376_ _22136_/X _22375_/X _14667_/B _22372_/X VGND VGND VPWR VPWR _23268_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24115_ _24203_/CLK _24115_/D HRESETn VGND VGND VPWR VPWR _16966_/A sky130_fd_sc_hd__dfrtp_4
X_21327_ _21258_/X _21326_/X _15747_/B _21323_/X VGND VGND VPWR VPWR _23886_/D sky130_fd_sc_hd__o22a_4
XFILLER_46_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12060_ _12088_/A _12060_/B _12060_/C VGND VGND VPWR VPWR _12061_/C sky130_fd_sc_hd__and3_4
X_24046_ _23692_/CLK _24046_/D VGND VGND VPWR VPWR _15686_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21258_ _21543_/A VGND VGND VPWR VPWR _21258_/X sky130_fd_sc_hd__buf_2
XFILLER_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20209_ _20444_/A VGND VGND VPWR VPWR _20209_/X sky130_fd_sc_hd__buf_2
XFILLER_81_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17635__B1 _17634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13537__A _13557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21431__B2 _21430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21189_ _20611_/X _21183_/X _13540_/B _21187_/X VGND VGND VPWR VPWR _23951_/D sky130_fd_sc_hd__o22a_4
XFILLER_49_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12441__A _12441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12160__B _23837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19865__A1_N _19531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15752__A _12777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12962_ _12974_/A _24051_/Q VGND VGND VPWR VPWR _12963_/C sky130_fd_sc_hd__or2_4
X_15750_ _15750_/A _15685_/B VGND VGND VPWR VPWR _15752_/B sky130_fd_sc_hd__or2_4
XFILLER_46_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21195__B1 _23947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16567__B _23612_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11913_ _12464_/A VGND VGND VPWR VPWR _11913_/X sky130_fd_sc_hd__buf_2
X_14701_ _15108_/A _14697_/X _14700_/X VGND VGND VPWR VPWR _14701_/X sky130_fd_sc_hd__or3_4
XFILLER_79_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18060__B1 _18016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15471__B _15471_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12893_ _13491_/A _12855_/X _12867_/X _12876_/X _12892_/X VGND VGND VPWR VPWR _12893_/X
+ sky130_fd_sc_hd__a32o_4
X_15681_ _12682_/X _15658_/X _15665_/X _15672_/X _15680_/X VGND VGND VPWR VPWR _15681_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_46_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17420_ _18525_/B _17419_/Y VGND VGND VPWR VPWR _17421_/A sky130_fd_sc_hd__or2_4
XANTENNA__13272__A _13202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11844_ _11843_/X VGND VGND VPWR VPWR _11844_/X sky130_fd_sc_hd__buf_2
X_14632_ _13927_/A _14632_/B VGND VGND VPWR VPWR _14632_/X sky130_fd_sc_hd__or2_4
XFILLER_73_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14563_ _11656_/A _14531_/X _14563_/C VGND VGND VPWR VPWR _14563_/X sky130_fd_sc_hd__and3_4
X_17351_ _17349_/Y _18466_/B VGND VGND VPWR VPWR _18395_/A sky130_fd_sc_hd__or2_4
XFILLER_18_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23808__CLK _23840_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17679__A _17681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11775_ _11734_/A _23582_/Q VGND VGND VPWR VPWR _11775_/X sky130_fd_sc_hd__or2_4
XANTENNA__22695__B1 _15835_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16302_ _11843_/X _11619_/X _16271_/X _11597_/X _16301_/X VGND VGND VPWR VPWR _16302_/X
+ sky130_fd_sc_hd__a32o_4
X_13514_ _12640_/A VGND VGND VPWR VPWR _13559_/A sky130_fd_sc_hd__buf_2
X_14494_ _13896_/A VGND VGND VPWR VPWR _14494_/X sky130_fd_sc_hd__buf_2
X_17282_ _17282_/A VGND VGND VPWR VPWR _17282_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19021_ _24367_/Q VGND VGND VPWR VPWR _19021_/Y sky130_fd_sc_hd__inv_2
X_13445_ _13450_/A _13531_/B VGND VGND VPWR VPWR _13446_/C sky130_fd_sc_hd__or2_4
X_16233_ _16233_/A VGND VGND VPWR VPWR _16233_/X sky130_fd_sc_hd__buf_2
XANTENNA__19894__A _19933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12616__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13376_ _12827_/A VGND VGND VPWR VPWR _13376_/X sky130_fd_sc_hd__buf_2
X_16164_ _16201_/A _16092_/B VGND VGND VPWR VPWR _16164_/X sky130_fd_sc_hd__or2_4
XANTENNA__18666__A2 _18664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20833__A _20833_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12327_ _12320_/A VGND VGND VPWR VPWR _12744_/A sky130_fd_sc_hd__buf_2
X_15115_ _15115_/A _15115_/B _15115_/C VGND VGND VPWR VPWR _15115_/X sky130_fd_sc_hd__or3_4
X_16095_ _16095_/A _16086_/X _16095_/C VGND VGND VPWR VPWR _16095_/X sky130_fd_sc_hd__or3_4
XANTENNA__14831__A _12575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21670__B2 _21666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15046_ _13986_/A _15042_/X _15046_/C VGND VGND VPWR VPWR _15047_/B sky130_fd_sc_hd__or3_4
X_19923_ _19909_/A _24142_/Q _22723_/A _19770_/X VGND VGND VPWR VPWR _24142_/D sky130_fd_sc_hd__o22a_4
X_12258_ _12742_/A VGND VGND VPWR VPWR _12728_/A sky130_fd_sc_hd__buf_2
XANTENNA__14550__B _14486_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19854_ _19643_/A _19853_/X VGND VGND VPWR VPWR _19854_/X sky130_fd_sc_hd__and2_4
XFILLER_29_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21422__B2 _21416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12189_ _11842_/A VGND VGND VPWR VPWR _12189_/X sky130_fd_sc_hd__buf_2
X_18805_ _17297_/X _18802_/X _24420_/Q _18803_/X VGND VGND VPWR VPWR _24420_/D sky130_fd_sc_hd__o22a_4
X_19785_ _19766_/B VGND VGND VPWR VPWR _19785_/Y sky130_fd_sc_hd__inv_2
X_16997_ _16997_/A VGND VGND VPWR VPWR _16997_/X sky130_fd_sc_hd__buf_2
XANTENNA__15662__A _12725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18736_ _17221_/Y _17808_/X VGND VGND VPWR VPWR _18736_/X sky130_fd_sc_hd__and2_4
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15948_ _15948_/A VGND VGND VPWR VPWR _15994_/A sky130_fd_sc_hd__buf_2
XANTENNA__21186__B1 _23953_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21725__A2 _21719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22922__A1 _18593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18667_ _18224_/A _18654_/X _18198_/A _18666_/X VGND VGND VPWR VPWR _18668_/A sky130_fd_sc_hd__o22a_4
X_15879_ _15879_/A _15879_/B VGND VGND VPWR VPWR _15881_/B sky130_fd_sc_hd__or2_4
XANTENNA__14278__A _15552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20933__B1 _20932_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13182__A _15697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17618_ _17605_/A _17295_/X _17618_/C _18578_/A VGND VGND VPWR VPWR _17619_/C sky130_fd_sc_hd__and4_4
XFILLER_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18598_ _18595_/Y _22921_/B _18595_/Y _22921_/B VGND VGND VPWR VPWR _18598_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21489__A1 _21277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17549_ _16376_/X _17549_/B VGND VGND VPWR VPWR _17550_/B sky130_fd_sc_hd__and2_4
XANTENNA__21489__B2 _21488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13910__A _13910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20560_ _20425_/X _20557_/Y _20559_/X _19010_/Y _20473_/X VGND VGND VPWR VPWR _20561_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_14_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19219_ _19219_/A _19219_/B VGND VGND VPWR VPWR _19220_/B sky130_fd_sc_hd__and2_4
XFILLER_34_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20491_ _20229_/A _20490_/X _20284_/X VGND VGND VPWR VPWR _20491_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__12526__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22230_ _22112_/X _22229_/X _15757_/B _22226_/X VGND VGND VPWR VPWR _22230_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20743__A _20743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22161_ _22081_/X _22158_/X _16792_/B _22155_/X VGND VGND VPWR VPWR _23419_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15837__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21661__B2 _21659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21112_ _21112_/A _21112_/B _21348_/C _21734_/B VGND VGND VPWR VPWR _21113_/A sky130_fd_sc_hd__or4_4
X_22092_ _22091_/X _22089_/X _16189_/B _22084_/X VGND VGND VPWR VPWR _23447_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15556__B _15556_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17880__A3 _17872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21043_ _20748_/X _21037_/X _24042_/Q _21041_/X VGND VGND VPWR VPWR _24042_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13357__A _12769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21413__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12261__A _12260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24323__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21964__A2 _21959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18867__B _20248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21574__A _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16668__A _16599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15572__A _12460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22994_ _22989_/A _22994_/B _22994_/C VGND VGND VPWR VPWR _22994_/X sky130_fd_sc_hd__and3_4
XFILLER_55_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16387__B _16387_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_42_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_42_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21945_ _21938_/A VGND VGND VPWR VPWR _21945_/X sky130_fd_sc_hd__buf_2
XFILLER_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18593__A1 _17878_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _21797_/X _21873_/X _23579_/Q _21870_/X VGND VGND VPWR VPWR _23579_/D sky130_fd_sc_hd__o22a_4
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ _23217_/CLK _21782_/X VGND VGND VPWR VPWR _23615_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _20681_/X _20826_/X _19072_/A _20625_/X VGND VGND VPWR VPWR _20827_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19542__B1 _19582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13820__A _15435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _24431_/Q IRQ[16] VGND VGND VPWR VPWR _11560_/X sky130_fd_sc_hd__and2_4
X_23546_ _23472_/CLK _21929_/X VGND VGND VPWR VPWR _16401_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20758_ _20516_/A VGND VGND VPWR VPWR _20758_/X sky130_fd_sc_hd__buf_2
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22429__B1 _15652_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23477_ _23315_/CLK _23477_/D VGND VGND VPWR VPWR _12542_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_52_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20689_ _20630_/A _20689_/B VGND VGND VPWR VPWR _20689_/Y sky130_fd_sc_hd__nor2_4
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13242_/A _23985_/Q VGND VGND VPWR VPWR _13231_/C sky130_fd_sc_hd__or2_4
X_22428_ _22416_/A VGND VGND VPWR VPWR _22428_/X sky130_fd_sc_hd__buf_2
XANTENNA__21101__B1 _14278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13161_ _15695_/A _13155_/X _13160_/X VGND VGND VPWR VPWR _13161_/X sky130_fd_sc_hd__or3_4
XANTENNA__15747__A _13129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20455__A2 _20454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22359_ _22107_/X _22354_/X _13296_/B _22358_/X VGND VGND VPWR VPWR _23280_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14651__A _15201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12112_ _12112_/A _12108_/X _12112_/C VGND VGND VPWR VPWR _12113_/B sky130_fd_sc_hd__or3_4
X_13092_ _13109_/A _13089_/X _13092_/C VGND VGND VPWR VPWR _13092_/X sky130_fd_sc_hd__and3_4
XANTENNA__15466__B _15403_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12043_ _16718_/A _12040_/X _12043_/C VGND VGND VPWR VPWR _12050_/B sky130_fd_sc_hd__and3_4
X_16920_ _17030_/B VGND VGND VPWR VPWR _17079_/A sky130_fd_sc_hd__inv_2
X_24029_ _24026_/CLK _24029_/D VGND VGND VPWR VPWR _24029_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13267__A _11671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_124_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR _23632_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21955__A2 _21952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16851_ _16851_/A _16847_/X _16850_/X VGND VGND VPWR VPWR _16851_/X sky130_fd_sc_hd__and3_4
XANTENNA__17681__B _17487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15802_ _12477_/X _15802_/B VGND VGND VPWR VPWR _15803_/C sky130_fd_sc_hd__or2_4
XANTENNA__15482__A _13097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19570_ _19570_/A VGND VGND VPWR VPWR _19706_/A sky130_fd_sc_hd__buf_2
X_16782_ _16618_/X _23963_/Q VGND VGND VPWR VPWR _16782_/X sky130_fd_sc_hd__or2_4
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13994_ _14010_/A VGND VGND VPWR VPWR _14841_/A sky130_fd_sc_hd__buf_2
XFILLER_24_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21707__A2 _21705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18521_ _17422_/D _18519_/X VGND VGND VPWR VPWR _18521_/X sky130_fd_sc_hd__or2_4
XFILLER_98_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15733_ _12795_/A _15677_/B VGND VGND VPWR VPWR _15733_/X sky130_fd_sc_hd__or2_4
X_12945_ _12976_/A _12945_/B VGND VGND VPWR VPWR _12945_/X sky130_fd_sc_hd__or2_4
XFILLER_4_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14098__A _14098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22380__A2 _22375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18452_ _17382_/B _18450_/X _18160_/A VGND VGND VPWR VPWR _18452_/Y sky130_fd_sc_hd__a21oi_4
X_15664_ _15664_/A _15662_/X _15663_/X VGND VGND VPWR VPWR _15665_/C sky130_fd_sc_hd__and3_4
XANTENNA__16595__B1 _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ _12876_/A _12870_/X _12876_/C VGND VGND VPWR VPWR _12876_/X sky130_fd_sc_hd__or3_4
X_17403_ _11634_/A _17344_/B _17402_/X _17125_/Y VGND VGND VPWR VPWR _17404_/B sky130_fd_sc_hd__a211o_4
X_14615_ _11894_/A _14696_/B VGND VGND VPWR VPWR _14615_/X sky130_fd_sc_hd__or2_4
X_11827_ _11827_/A _23486_/Q VGND VGND VPWR VPWR _11830_/B sky130_fd_sc_hd__or2_4
X_18383_ _18383_/A _18383_/B VGND VGND VPWR VPWR _18383_/X sky130_fd_sc_hd__and2_4
X_15595_ _15631_/A _15595_/B _15594_/X VGND VGND VPWR VPWR _15596_/C sky130_fd_sc_hd__and3_4
XFILLER_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14826__A _13872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13730__A _15491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _15381_/X _17863_/A _17324_/X _17333_/X VGND VGND VPWR VPWR _17334_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _16069_/A VGND VGND VPWR VPWR _11758_/X sky130_fd_sc_hd__buf_2
X_14546_ _13901_/A _14538_/X _14546_/C VGND VGND VPWR VPWR _14546_/X sky130_fd_sc_hd__and3_4
XFILLER_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17265_ _17264_/X VGND VGND VPWR VPWR _17781_/B sky130_fd_sc_hd__inv_2
X_11689_ _12837_/A VGND VGND VPWR VPWR _16447_/A sky130_fd_sc_hd__buf_2
X_14477_ _12512_/A _14477_/B VGND VGND VPWR VPWR _14477_/X sky130_fd_sc_hd__or2_4
XFILLER_35_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12346__A _12794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19004_ _24370_/Q VGND VGND VPWR VPWR _19004_/Y sky130_fd_sc_hd__inv_2
X_16216_ _16223_/A _23095_/Q VGND VGND VPWR VPWR _16216_/X sky130_fd_sc_hd__or2_4
X_13428_ _13428_/A _23503_/Q VGND VGND VPWR VPWR _13428_/X sky130_fd_sc_hd__or2_4
XANTENNA__21659__A _21659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17196_ _15909_/B _17100_/X _17195_/Y _17065_/X VGND VGND VPWR VPWR _17196_/X sky130_fd_sc_hd__o22a_4
XFILLER_31_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13359_ _13358_/X _13287_/B VGND VGND VPWR VPWR _13362_/B sky130_fd_sc_hd__or2_4
X_16147_ _16147_/A _16147_/B _16147_/C VGND VGND VPWR VPWR _16147_/X sky130_fd_sc_hd__and3_4
XANTENNA__15657__A _12720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21643__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14561__A _13770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16078_ _16008_/Y _16077_/X VGND VGND VPWR VPWR _16081_/A sky130_fd_sc_hd__and2_4
XFILLER_5_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22199__A2 _22172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18968__A _18999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13177__A _13317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15029_ _15006_/A _15097_/B VGND VGND VPWR VPWR _15029_/X sky130_fd_sc_hd__or2_4
X_19906_ _19899_/X _24155_/Q _19903_/X _20317_/B VGND VGND VPWR VPWR _19906_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12081__A _11992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21946__A2 _21945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19837_ _19445_/A _19836_/X VGND VGND VPWR VPWR _19837_/X sky130_fd_sc_hd__or2_4
XFILLER_116_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13905__A _13909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19768_ _19710_/X _19763_/X _19767_/X _16599_/X _19697_/X VGND VGND VPWR VPWR _24175_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_68_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21159__B1 _14873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18719_ _18443_/A _17611_/Y _18715_/X _18718_/Y VGND VGND VPWR VPWR _18719_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_5_29_0_HCLK clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19699_ HRDATA[6] VGND VGND VPWR VPWR _19699_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16000__B _23704_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17405__A2_N _17013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22371__A2 _22368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21730_ _21574_/X _21726_/X _23649_/Q _21687_/X VGND VGND VPWR VPWR _23649_/D sky130_fd_sc_hd__o22a_4
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21661_ _21541_/X _21655_/X _13487_/B _21659_/X VGND VGND VPWR VPWR _21661_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23400_ _23368_/CLK _22188_/X VGND VGND VPWR VPWR _23400_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18208__A _18267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22123__A2 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20612_ _20511_/X _20611_/X _13566_/B _20592_/X VGND VGND VPWR VPWR _20612_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13640__A _13659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24380_ _24435_/CLK _18881_/X HRESETn VGND VGND VPWR VPWR _24380_/Q sky130_fd_sc_hd__dfstp_4
X_21592_ _21506_/X _21591_/X _23741_/Q _21588_/X VGND VGND VPWR VPWR _23741_/D sky130_fd_sc_hd__o22a_4
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21331__B1 _23883_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23331_ _23907_/CLK _23331_/D VGND VGND VPWR VPWR _14790_/B sky130_fd_sc_hd__dfxtp_4
X_20543_ _20403_/X _20542_/X _19223_/A _20497_/X VGND VGND VPWR VPWR _20543_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21882__B2 _21877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23262_ _23358_/CLK _22389_/X VGND VGND VPWR VPWR _11705_/B sky130_fd_sc_hd__dfxtp_4
X_20474_ _20425_/X _20469_/Y _20472_/X _18985_/Y _20473_/X VGND VGND VPWR VPWR _20475_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__17766__B _17274_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16670__B _24092_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22213_ _22083_/X _22208_/X _16423_/B _22212_/X VGND VGND VPWR VPWR _22213_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23193_ _23130_/CLK _23193_/D VGND VGND VPWR VPWR _16248_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14471__A _12862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23503__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22144_ _22143_/X _22137_/X _15150_/B _22071_/X VGND VGND VPWR VPWR _23425_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18878__A _18892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13087__A _13087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22075_ _20314_/A VGND VGND VPWR VPWR _22075_/X sky130_fd_sc_hd__buf_2
XFILLER_0_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21026_ _20464_/X _21023_/X _24054_/Q _21020_/X VGND VGND VPWR VPWR _21026_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13815__A _13623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22977_ _22977_/A VGND VGND VPWR VPWR HADDR[16] sky130_fd_sc_hd__inv_2
XANTENNA__22362__A2 _22361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24009__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12730_ _12730_/A _12819_/B VGND VGND VPWR VPWR _12730_/X sky130_fd_sc_hd__or2_4
XFILLER_83_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21928_ _21920_/X VGND VGND VPWR VPWR _21928_/X sky130_fd_sc_hd__buf_2
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12661_ _12622_/X _12661_/B VGND VGND VPWR VPWR _12662_/C sky130_fd_sc_hd__or2_4
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21859_ _21574_/A VGND VGND VPWR VPWR _21859_/X sky130_fd_sc_hd__buf_2
XFILLER_43_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14646__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22114__A2 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _13966_/A VGND VGND VPWR VPWR _15413_/A sky130_fd_sc_hd__buf_2
X_14400_ _15623_/A _14400_/B _14400_/C VGND VGND VPWR VPWR _14404_/B sky130_fd_sc_hd__and3_4
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13550__A _13550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12591_/X _12462_/B VGND VGND VPWR VPWR _12592_/X sky130_fd_sc_hd__or2_4
X_15380_ _15379_/X VGND VGND VPWR VPWR _15380_/Y sky130_fd_sc_hd__inv_2
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24159__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _20470_/A IRQ[22] VGND VGND VPWR VPWR _20160_/A sky130_fd_sc_hd__and2_4
X_14331_ _15574_/A _14410_/B VGND VGND VPWR VPWR _14331_/X sky130_fd_sc_hd__or2_4
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_49_0_HCLK clkbuf_6_24_0_HCLK/X VGND VGND VPWR VPWR _24011_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23529_ _23910_/CLK _23529_/D VGND VGND VPWR VPWR _23529_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17957__A _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12166__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _14261_/X VGND VGND VPWR VPWR _14263_/A sky130_fd_sc_hd__inv_2
X_17050_ _17072_/A VGND VGND VPWR VPWR _17083_/B sky130_fd_sc_hd__inv_2
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16580__B _24092_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13213_ _12794_/A _13145_/B VGND VGND VPWR VPWR _13214_/C sky130_fd_sc_hd__or2_4
X_16001_ _13477_/X VGND VGND VPWR VPWR _16002_/A sky130_fd_sc_hd__buf_2
X_14193_ _14225_/A _23177_/Q VGND VGND VPWR VPWR _14195_/B sky130_fd_sc_hd__or2_4
XANTENNA__21625__B2 _21623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14381__A _13710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13144_ _12693_/A _13144_/B VGND VGND VPWR VPWR _13144_/X sky130_fd_sc_hd__or2_4
XFILLER_48_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18197__A2_N _18196_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13075_ _13112_/A _13075_/B VGND VGND VPWR VPWR _13075_/X sky130_fd_sc_hd__or2_4
X_17952_ _17951_/A _17894_/D VGND VGND VPWR VPWR _17952_/X sky130_fd_sc_hd__and2_4
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12026_ _16113_/A _12026_/B _12026_/C VGND VGND VPWR VPWR _12027_/B sky130_fd_sc_hd__or3_4
X_16903_ _12034_/A _16903_/B _16903_/C _16903_/D VGND VGND VPWR VPWR _16903_/X sky130_fd_sc_hd__or4_4
XFILLER_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17883_ _17769_/X _17882_/Y VGND VGND VPWR VPWR _17883_/X sky130_fd_sc_hd__and2_4
XFILLER_117_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22050__B2 _22049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22103__A _20552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19622_ _19622_/A VGND VGND VPWR VPWR _19622_/Y sky130_fd_sc_hd__inv_2
X_16834_ _13277_/X _16833_/Y VGND VGND VPWR VPWR _16834_/X sky130_fd_sc_hd__or2_4
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19553_ _19553_/A HRDATA[12] VGND VGND VPWR VPWR _19553_/X sky130_fd_sc_hd__and2_4
XANTENNA__21942__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16765_ _16747_/X _16763_/X _16765_/C VGND VGND VPWR VPWR _16771_/B sky130_fd_sc_hd__and3_4
XFILLER_98_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13977_ _12209_/A _23626_/Q VGND VGND VPWR VPWR _13977_/X sky130_fd_sc_hd__or2_4
XFILLER_0_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18504_ _17407_/X _18501_/X _17878_/X _18503_/X VGND VGND VPWR VPWR _18505_/A sky130_fd_sc_hd__a211o_4
XFILLER_62_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22353__A2 _22347_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15716_ _13109_/A _15714_/X _15715_/X VGND VGND VPWR VPWR _15716_/X sky130_fd_sc_hd__and3_4
X_12928_ _12591_/X _12928_/B VGND VGND VPWR VPWR _12930_/B sky130_fd_sc_hd__or2_4
X_19484_ _19441_/A VGND VGND VPWR VPWR _19872_/B sky130_fd_sc_hd__inv_2
X_16696_ _16542_/A _16696_/B _16696_/C VGND VGND VPWR VPWR _16696_/X sky130_fd_sc_hd__or3_4
XANTENNA__21561__B1 _23751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20558__A _20558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18435_ _18381_/A VGND VGND VPWR VPWR _18435_/X sky130_fd_sc_hd__buf_2
XFILLER_92_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15647_ _15646_/X VGND VGND VPWR VPWR _15649_/B sky130_fd_sc_hd__inv_2
XFILLER_62_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12859_ _12859_/A _12857_/X _12859_/C VGND VGND VPWR VPWR _12859_/X sky130_fd_sc_hd__and3_4
XANTENNA__18028__A _17090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13460__A _11980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18366_ _17962_/A _18364_/X _18183_/X _18365_/X VGND VGND VPWR VPWR _18367_/A sky130_fd_sc_hd__o22a_4
X_15578_ _15578_/A _15576_/X _15578_/C VGND VGND VPWR VPWR _15579_/C sky130_fd_sc_hd__and3_4
XFILLER_37_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14275__B _14275_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17317_ _17143_/X _17201_/A VGND VGND VPWR VPWR _18656_/B sky130_fd_sc_hd__or2_4
X_14529_ _13754_/A _14525_/X _14529_/C VGND VGND VPWR VPWR _14529_/X sky130_fd_sc_hd__or3_4
XFILLER_50_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18297_ _18297_/A _18297_/B VGND VGND VPWR VPWR _18298_/D sky130_fd_sc_hd__and2_4
XANTENNA__21864__B2 _21787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16771__A _11834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17248_ _17224_/X VGND VGND VPWR VPWR _17249_/A sky130_fd_sc_hd__inv_2
Xclkbuf_6_6_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17179_ _17178_/X VGND VGND VPWR VPWR _17179_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12804__A _12769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18493__B1 _18398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21092__A2 _21089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20190_ _20190_/A VGND VGND VPWR VPWR _20196_/A sky130_fd_sc_hd__inv_2
XFILLER_69_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22041__B2 _22035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22592__A2 _22586_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22900_ _22968_/A VGND VGND VPWR VPWR _23051_/A sky130_fd_sc_hd__buf_2
X_23880_ _23816_/CLK _23880_/D VGND VGND VPWR VPWR _13651_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_99_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22831_ _22777_/X VGND VGND VPWR VPWR _22831_/X sky130_fd_sc_hd__buf_2
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18864__C _18864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15850__A _13522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22762_ _24100_/Q VGND VGND VPWR VPWR _22763_/A sky130_fd_sc_hd__inv_2
XFILLER_65_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21552__B1 _15530_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21713_ _21543_/X _21712_/X _15737_/B _21709_/X VGND VGND VPWR VPWR _23662_/D sky130_fd_sc_hd__o22a_4
XFILLER_80_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _22686_/A VGND VGND VPWR VPWR _22693_/X sky130_fd_sc_hd__buf_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21644_ _21512_/X _21641_/X _23707_/Q _21638_/X VGND VGND VPWR VPWR _23707_/D sky130_fd_sc_hd__o22a_4
X_24432_ _23326_/CLK _24432_/D HRESETn VGND VGND VPWR VPWR _24432_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22683__A _22683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24363_ _24365_/CLK _24363_/D HRESETn VGND VGND VPWR VPWR _24363_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__17777__A _18062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11602__B _18866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ _21574_/X _21568_/X _23745_/Q _21515_/A VGND VGND VPWR VPWR _21575_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18720__A1 _18390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23314_ _23314_/CLK _22312_/X VGND VGND VPWR VPWR _23314_/Q sky130_fd_sc_hd__dfxtp_4
X_20526_ _20518_/X _20524_/X _11524_/A _20525_/X VGND VGND VPWR VPWR _20526_/X sky130_fd_sc_hd__o22a_4
X_24294_ _24299_/CLK _24294_/D HRESETn VGND VGND VPWR VPWR _24294_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14913__B _23840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21607__A1 _21534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23245_ _23564_/CLK _23245_/D VGND VGND VPWR VPWR _15845_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_101_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20457_ _18162_/X _20447_/X _20319_/X _20456_/Y VGND VGND VPWR VPWR _20457_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21607__B2 _21602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12714__A _15812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21083__A2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23176_ _23079_/CLK _23176_/D VGND VGND VPWR VPWR _13712_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20388_ _20387_/X VGND VGND VPWR VPWR _20388_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22280__B2 _22276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22127_ _22127_/A VGND VGND VPWR VPWR _22127_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22058_ _21850_/X _22052_/X _14476_/B _22056_/X VGND VGND VPWR VPWR _23461_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22032__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18787__A1 _17194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13900_ _13884_/A _13896_/X _13900_/C VGND VGND VPWR VPWR _13900_/X sky130_fd_sc_hd__or3_4
X_21009_ _21348_/A _21112_/B _21162_/C _21734_/B VGND VGND VPWR VPWR _21009_/X sky130_fd_sc_hd__or4_4
XANTENNA__13545__A _13507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14880_ _14880_/A _23552_/Q VGND VGND VPWR VPWR _14880_/X sky130_fd_sc_hd__or2_4
XFILLER_87_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21762__A _21755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13831_ _12203_/A _13831_/B VGND VGND VPWR VPWR _13833_/B sky130_fd_sc_hd__or2_4
XFILLER_29_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18539__A1 _18142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19736__B1 _20895_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15760__A _11680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16550_ _16567_/A _16550_/B VGND VGND VPWR VPWR _16550_/X sky130_fd_sc_hd__or2_4
XFILLER_112_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13762_ _13738_/A _13762_/B _13761_/X VGND VGND VPWR VPWR _13762_/X sky130_fd_sc_hd__or3_4
Xclkbuf_5_12_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_15501_ _15477_/A _23084_/Q VGND VGND VPWR VPWR _15501_/X sky130_fd_sc_hd__or2_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12713_ _12713_/A _12709_/X _12712_/X VGND VGND VPWR VPWR _12713_/X sky130_fd_sc_hd__or3_4
X_16481_ _11666_/X _16463_/X _16481_/C VGND VGND VPWR VPWR _16513_/B sky130_fd_sc_hd__or3_4
X_13693_ _14010_/A VGND VGND VPWR VPWR _13694_/A sky130_fd_sc_hd__buf_2
X_18220_ _17456_/Y _18219_/X VGND VGND VPWR VPWR _18220_/X sky130_fd_sc_hd__or2_4
XFILLER_43_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23549__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15432_ _15432_/A _15432_/B VGND VGND VPWR VPWR _15434_/B sky130_fd_sc_hd__or2_4
X_12644_ _12963_/A _12642_/X _12644_/C VGND VGND VPWR VPWR _12645_/C sky130_fd_sc_hd__and3_4
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22099__B2 _22096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22593__A _22586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18151_ _17584_/Y _18151_/B VGND VGND VPWR VPWR _18151_/X sky130_fd_sc_hd__and2_4
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12575_ _12575_/A VGND VGND VPWR VPWR _13700_/A sky130_fd_sc_hd__buf_2
X_15363_ _15332_/A _15303_/B VGND VGND VPWR VPWR _15365_/B sky130_fd_sc_hd__or2_4
XANTENNA__21846__B2 _21836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16591__A _12025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17102_ _17101_/X VGND VGND VPWR VPWR _18713_/A sky130_fd_sc_hd__buf_2
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ _11859_/A _14310_/X _14313_/X VGND VGND VPWR VPWR _14314_/X sky130_fd_sc_hd__or3_4
XFILLER_89_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11526_ _18982_/A _11525_/X VGND VGND VPWR VPWR _11526_/X sky130_fd_sc_hd__or2_4
X_18082_ _18082_/A VGND VGND VPWR VPWR _18082_/X sky130_fd_sc_hd__buf_2
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15294_ _14734_/A _15292_/X _15293_/X VGND VGND VPWR VPWR _15294_/X sky130_fd_sc_hd__and3_4
XFILLER_32_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23699__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17033_ _17033_/A VGND VGND VPWR VPWR _17036_/A sky130_fd_sc_hd__inv_2
X_14245_ _14205_/A _23785_/Q VGND VGND VPWR VPWR _14246_/C sky130_fd_sc_hd__or2_4
XFILLER_67_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12624__A _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15000__A _14151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14176_ _11638_/A VGND VGND VPWR VPWR _14190_/A sky130_fd_sc_hd__buf_2
XANTENNA__22271__B2 _22269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13127_ _13115_/A _24082_/Q VGND VGND VPWR VPWR _13128_/C sky130_fd_sc_hd__or2_4
X_18984_ _18982_/Y _18983_/Y _11526_/X VGND VGND VPWR VPWR _18984_/X sky130_fd_sc_hd__o21a_4
XFILLER_3_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13058_ _11842_/A _11618_/A _13027_/X _11596_/A _13057_/X VGND VGND VPWR VPWR _13059_/A
+ sky130_fd_sc_hd__a32o_4
X_17935_ _17800_/X _17934_/Y _17252_/X VGND VGND VPWR VPWR _17935_/X sky130_fd_sc_hd__o21a_4
XFILLER_41_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18778__A1 _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12009_ _11962_/X VGND VGND VPWR VPWR _16536_/A sky130_fd_sc_hd__buf_2
XANTENNA__13455__A _12464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22574__A2 _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17866_ _17254_/X VGND VGND VPWR VPWR _17866_/X sky130_fd_sc_hd__buf_2
XFILLER_94_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20585__A1 _18334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23079__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21782__B1 _23615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16817_ _16682_/X _16816_/X VGND VGND VPWR VPWR _16817_/X sky130_fd_sc_hd__or2_4
X_19605_ _19876_/B _19600_/X _19511_/B _19822_/A VGND VGND VPWR VPWR _19605_/X sky130_fd_sc_hd__o22a_4
X_17797_ _17837_/A VGND VGND VPWR VPWR _17797_/X sky130_fd_sc_hd__buf_2
XFILLER_19_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19536_ _19536_/A _19536_/B VGND VGND VPWR VPWR _19537_/B sky130_fd_sc_hd__or2_4
XANTENNA__15670__A _15693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16748_ _11754_/X VGND VGND VPWR VPWR _16772_/A sky130_fd_sc_hd__buf_2
XFILLER_81_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16485__B _23610_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19467_ _19517_/A VGND VGND VPWR VPWR _19523_/A sky130_fd_sc_hd__inv_2
X_16679_ _16596_/Y _16678_/X VGND VGND VPWR VPWR _16682_/A sky130_fd_sc_hd__and2_4
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13190__A _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18418_ _18418_/A _18418_/B VGND VGND VPWR VPWR _18418_/X sky130_fd_sc_hd__or2_4
XANTENNA__14567__A2 _14564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19398_ _19396_/X _18484_/Y _19396_/X _24202_/Q VGND VGND VPWR VPWR _19398_/X sky130_fd_sc_hd__a2bb2o_4
X_18349_ _18349_/A _18349_/B VGND VGND VPWR VPWR _18350_/B sky130_fd_sc_hd__or2_4
XANTENNA__21837__B2 _21836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24138__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21360_ _21229_/X _21355_/X _16438_/B _21359_/X VGND VGND VPWR VPWR _21360_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_32_0_HCLK clkbuf_7_33_0_HCLK/A VGND VGND VPWR VPWR _23270_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15829__B _15829_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20311_ _24253_/Q _20283_/X _20310_/X VGND VGND VPWR VPWR _20312_/B sky130_fd_sc_hd__o21a_4
XFILLER_102_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_95_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR _23514_/CLK sky130_fd_sc_hd__clkbuf_1
X_21291_ _21291_/A VGND VGND VPWR VPWR _21291_/X sky130_fd_sc_hd__buf_2
XANTENNA__12534__A _13041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23030_ _23014_/X _18012_/X _23026_/X _23029_/X VGND VGND VPWR VPWR _23031_/A sky130_fd_sc_hd__a211o_4
X_20242_ _11621_/X _20248_/A VGND VGND VPWR VPWR _20242_/X sky130_fd_sc_hd__or2_4
XANTENNA__20751__A _20512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12750__A1 _12716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20173_ _11622_/X _20173_/B VGND VGND VPWR VPWR _20173_/X sky130_fd_sc_hd__and2_4
XANTENNA__19317__A _19317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_HCLK clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22014__B2 _21970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18769__A1 _11837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23932_ _23931_/CLK _21226_/X VGND VGND VPWR VPWR _23932_/Q sky130_fd_sc_hd__dfxtp_4
X_23863_ _23632_/CLK _23863_/D VGND VGND VPWR VPWR _16220_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13058__A2 _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16676__A _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17992__A2 _17568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15580__A _13682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19052__A _18994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22814_ _22779_/X VGND VGND VPWR VPWR _22814_/X sky130_fd_sc_hd__buf_2
XFILLER_57_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23794_ _23794_/CLK _21472_/X VGND VGND VPWR VPWR _13120_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_37_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22745_ SYSTICKCLKDIV[5] _24101_/Q _22743_/Y _22744_/Y VGND VGND VPWR VPWR _22746_/D
+ sky130_fd_sc_hd__o22a_4
XFILLER_73_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14196__A _14207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12709__A _12709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18891__A _18891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11613__A _15413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22676_ _22668_/X VGND VGND VPWR VPWR _22676_/X sky130_fd_sc_hd__buf_2
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21627_ _21567_/X _21626_/X _14654_/B _21623_/X VGND VGND VPWR VPWR _23716_/D sky130_fd_sc_hd__o22a_4
X_24415_ _24425_/CLK _24415_/D HRESETn VGND VGND VPWR VPWR _11540_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12360_ _12360_/A _12236_/B VGND VGND VPWR VPWR _12362_/B sky130_fd_sc_hd__or2_4
X_21558_ _21843_/A VGND VGND VPWR VPWR _21558_/X sky130_fd_sc_hd__buf_2
X_24346_ _24344_/CLK _18957_/X HRESETn VGND VGND VPWR VPWR _24346_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__15739__B _15667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20509_ _20509_/A VGND VGND VPWR VPWR _20509_/X sky130_fd_sc_hd__buf_2
X_12291_ _12695_/A _12289_/X _12290_/X VGND VGND VPWR VPWR _12291_/X sky130_fd_sc_hd__and3_4
X_24277_ _24277_/CLK _24277_/D HRESETn VGND VGND VPWR VPWR _24277_/Q sky130_fd_sc_hd__dfrtp_4
X_21489_ _21277_/X _21484_/X _14328_/B _21488_/X VGND VGND VPWR VPWR _21489_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12444__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14030_ _11646_/A VGND VGND VPWR VPWR _14031_/A sky130_fd_sc_hd__buf_2
XFILLER_107_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23228_ _23324_/CLK _23228_/D VGND VGND VPWR VPWR _16672_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21056__A2 _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12163__B _23421_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11544__A2 IRQ[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23159_ _23313_/CLK _23159_/D VGND VGND VPWR VPWR _16186_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15755__A _15725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22005__B2 _21999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15981_ _15984_/A _15981_/B VGND VGND VPWR VPWR _15981_/X sky130_fd_sc_hd__or2_4
XFILLER_114_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17720_ _17720_/A _17290_/X VGND VGND VPWR VPWR _17720_/X sky130_fd_sc_hd__or2_4
XANTENNA__13275__A _13059_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22556__A2 _22550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14932_ _14937_/A _14868_/B VGND VGND VPWR VPWR _14932_/X sky130_fd_sc_hd__or2_4
XANTENNA__20567__A1 _18309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21764__B1 _15902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17651_ _17651_/A _17651_/B VGND VGND VPWR VPWR _17651_/X sky130_fd_sc_hd__or2_4
X_14863_ _13953_/A _14863_/B VGND VGND VPWR VPWR _14863_/X sky130_fd_sc_hd__or2_4
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19709__B1 _12096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16602_ _16799_/A _16602_/B VGND VGND VPWR VPWR _16602_/X sky130_fd_sc_hd__or2_4
XANTENNA__15490__A _15497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13814_ _13622_/A _13814_/B VGND VGND VPWR VPWR _13814_/X sky130_fd_sc_hd__or2_4
XFILLER_29_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17582_ _17547_/X _17581_/Y _17957_/B _17550_/B VGND VGND VPWR VPWR _17582_/X sky130_fd_sc_hd__a211o_4
XFILLER_63_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14794_ _13872_/A _14794_/B VGND VGND VPWR VPWR _14796_/B sky130_fd_sc_hd__or2_4
X_19321_ _19328_/A VGND VGND VPWR VPWR _19321_/X sky130_fd_sc_hd__buf_2
XFILLER_17_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16533_ _12112_/A _16533_/B _16533_/C VGND VGND VPWR VPWR _16533_/X sky130_fd_sc_hd__or3_4
X_13745_ _12937_/A _13745_/B VGND VGND VPWR VPWR _13746_/C sky130_fd_sc_hd__or2_4
XANTENNA__19897__A _23027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12619__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19252_ _24278_/Q _19226_/X _19251_/Y VGND VGND VPWR VPWR _19252_/X sky130_fd_sc_hd__o21a_4
X_16464_ _16464_/A _16404_/B VGND VGND VPWR VPWR _16464_/X sky130_fd_sc_hd__or2_4
X_13676_ _13635_/A _13757_/B VGND VGND VPWR VPWR _13676_/X sky130_fd_sc_hd__or2_4
X_18203_ _18203_/A VGND VGND VPWR VPWR _18204_/A sky130_fd_sc_hd__buf_2
X_15415_ _13632_/A _15415_/B _15415_/C VGND VGND VPWR VPWR _15419_/B sky130_fd_sc_hd__and3_4
XFILLER_31_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12627_ _12604_/A _12627_/B VGND VGND VPWR VPWR _12629_/B sky130_fd_sc_hd__or2_4
X_19183_ _19118_/B VGND VGND VPWR VPWR _19183_/Y sky130_fd_sc_hd__inv_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16395_ _16394_/X VGND VGND VPWR VPWR _16400_/A sky130_fd_sc_hd__buf_2
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14834__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18134_ _18062_/A _17586_/C VGND VGND VPWR VPWR _18134_/X sky130_fd_sc_hd__or2_4
X_15346_ _14020_/A _15346_/B _15345_/X VGND VGND VPWR VPWR _15346_/X sky130_fd_sc_hd__and3_4
XFILLER_106_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18696__B1 _18500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12558_ _11980_/A _12528_/X _12541_/X _12549_/X _12557_/X VGND VGND VPWR VPWR _12558_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22492__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_19_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11509_ _11509_/A _11508_/X VGND VGND VPWR VPWR _11510_/B sky130_fd_sc_hd__or2_4
X_18065_ _18206_/A _17556_/X VGND VGND VPWR VPWR _18065_/X sky130_fd_sc_hd__and2_4
X_15277_ _15023_/A _15277_/B VGND VGND VPWR VPWR _15277_/X sky130_fd_sc_hd__or2_4
XANTENNA__12354__A _11680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12489_ _12872_/A _12627_/B VGND VGND VPWR VPWR _12489_/X sky130_fd_sc_hd__or2_4
X_17016_ _17015_/X VGND VGND VPWR VPWR _17016_/X sky130_fd_sc_hd__buf_2
XANTENNA__19372__A2_N _18020_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14228_ _14207_/A VGND VGND VPWR VPWR _14246_/A sky130_fd_sc_hd__buf_2
XFILLER_67_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21047__A2 _21044_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22244__B2 _22240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20571__A _20534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11535__A2 IRQ[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15665__A _15688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14159_ _15041_/A VGND VGND VPWR VPWR _15030_/A sky130_fd_sc_hd__buf_2
XFILLER_86_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18967_ _24376_/Q VGND VGND VPWR VPWR _18967_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13185__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17918_ _17798_/X _17909_/X _17823_/X _17917_/X VGND VGND VPWR VPWR _17918_/X sky130_fd_sc_hd__o22a_4
X_18898_ _18898_/A VGND VGND VPWR VPWR _18898_/X sky130_fd_sc_hd__buf_2
X_17849_ _17813_/X _17847_/X _17818_/X _17848_/X VGND VGND VPWR VPWR _17849_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__18620__B1 _17782_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16496__A _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20860_ _20760_/X _20859_/X _24325_/Q _20767_/X VGND VGND VPWR VPWR _20860_/X sky130_fd_sc_hd__o22a_4
X_19519_ _19458_/X _19518_/X HRDATA[5] _19462_/X VGND VGND VPWR VPWR _19866_/B sky130_fd_sc_hd__o22a_4
X_20791_ _18548_/X _20680_/X _20731_/X _20790_/Y VGND VGND VPWR VPWR _20791_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17187__B1 _13591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22530_ _22403_/X _22529_/X _16019_/B _22526_/X VGND VGND VPWR VPWR _23192_/D sky130_fd_sc_hd__o22a_4
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19600__A _19800_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12248__B _12248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22461_ _22460_/X _22452_/X _14856_/B _22386_/X VGND VGND VPWR VPWR _22461_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14744__A _13800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18216__A _18216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21412_ _21419_/A VGND VGND VPWR VPWR _21412_/X sky130_fd_sc_hd__buf_2
X_24200_ _24473_/CLK _19401_/X HRESETn VGND VGND VPWR VPWR _24200_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21286__A2 _21283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22392_ _22416_/A VGND VGND VPWR VPWR _22392_/X sky130_fd_sc_hd__buf_2
XANTENNA__15559__B _23115_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24131_ _23522_/CLK _20004_/Y HRESETn VGND VGND VPWR VPWR _24131_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21343_ _21287_/X _21340_/X _15282_/B _21337_/X VGND VGND VPWR VPWR _23874_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12264__A _12255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24062_ _23774_/CLK _21014_/X VGND VGND VPWR VPWR _24062_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21038__A2 _21037_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21274_ _21273_/X _21271_/X _13723_/B _21266_/X VGND VGND VPWR VPWR _21274_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22235__B2 _22233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23013_ _23013_/A VGND VGND VPWR VPWR HADDR[22] sky130_fd_sc_hd__inv_2
X_20225_ _16910_/X _16913_/X _20223_/X _20224_/X VGND VGND VPWR VPWR _20226_/B sky130_fd_sc_hd__and4_4
XFILLER_104_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17111__B1 _12892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20156_ _20156_/A _20155_/X VGND VGND VPWR VPWR _20156_/X sky130_fd_sc_hd__or2_4
XFILLER_44_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13279__A2 _13278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12711__B _12711_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22538__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20087_ _20098_/B VGND VGND VPWR VPWR _20087_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17414__A1 _17411_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23915_ _23915_/CLK _21267_/X VGND VGND VPWR VPWR _23915_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17414__B2 _17413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21210__A2 _21183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14919__A _14177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13823__A _15411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11860_ _13004_/A VGND VGND VPWR VPWR _12458_/A sky130_fd_sc_hd__buf_2
X_23846_ _23781_/CLK _21388_/X VGND VGND VPWR VPWR _14410_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11791_ _11780_/X _23550_/Q VGND VGND VPWR VPWR _11791_/X sky130_fd_sc_hd__or2_4
XFILLER_92_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20989_ _20987_/X _20988_/X _20240_/X VGND VGND VPWR VPWR _20989_/Y sky130_fd_sc_hd__o21ai_4
X_23777_ _23487_/CLK _23777_/D VGND VGND VPWR VPWR _15177_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12439__A _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17717__A2 _17385_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18914__A1 _14564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22710__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13530_ _13558_/A _13530_/B VGND VGND VPWR VPWR _13532_/B sky130_fd_sc_hd__or2_4
XFILLER_25_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22728_ SYSTICKCLKDIV[7] VGND VGND VPWR VPWR _22728_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20721__A1 _24203_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23032__A _23027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13461_ _11851_/X _13433_/X _13441_/X _13452_/X _13460_/X VGND VGND VPWR VPWR _13461_/X
+ sky130_fd_sc_hd__a32o_4
X_22659_ _22454_/X _22657_/X _14762_/B _22654_/X VGND VGND VPWR VPWR _23107_/D sky130_fd_sc_hd__o22a_4
X_15200_ _14202_/A _15200_/B _15199_/X VGND VGND VPWR VPWR _15217_/B sky130_fd_sc_hd__and3_4
X_12412_ _12412_/A VGND VGND VPWR VPWR _12596_/A sky130_fd_sc_hd__buf_2
X_16180_ _16180_/A _16168_/X _16180_/C VGND VGND VPWR VPWR _16200_/B sky130_fd_sc_hd__and3_4
X_13392_ _13352_/X _13318_/B VGND VGND VPWR VPWR _13394_/B sky130_fd_sc_hd__or2_4
XANTENNA__22474__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15131_ _13972_/A _15127_/X _15130_/X VGND VGND VPWR VPWR _15131_/X sky130_fd_sc_hd__or3_4
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12343_ _12791_/A VGND VGND VPWR VPWR _12826_/A sky130_fd_sc_hd__buf_2
X_24329_ _24330_/CLK _24329_/D HRESETn VGND VGND VPWR VPWR _24329_/Q sky130_fd_sc_hd__dfstp_4
X_12274_ _12710_/A _12274_/B VGND VGND VPWR VPWR _12274_/X sky130_fd_sc_hd__or2_4
X_15062_ _11723_/A _15062_/B _15062_/C VGND VGND VPWR VPWR _15062_/X sky130_fd_sc_hd__and3_4
XANTENNA__20391__A _20484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14013_ _14815_/A _14011_/X _14013_/C VGND VGND VPWR VPWR _14013_/X sky130_fd_sc_hd__and3_4
XFILLER_5_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15485__A _11664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19870_ _19449_/X _19866_/X _19869_/Y _20206_/A _19490_/X VGND VGND VPWR VPWR _19870_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_9_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12902__A _12520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20788__B2 _20686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18821_ _18835_/A VGND VGND VPWR VPWR _18821_/X sky130_fd_sc_hd__buf_2
XANTENNA__13717__B _24008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18752_ _18752_/A VGND VGND VPWR VPWR _18752_/X sky130_fd_sc_hd__buf_2
XFILLER_27_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15964_ _11884_/X _23928_/Q VGND VGND VPWR VPWR _15964_/X sky130_fd_sc_hd__or2_4
XFILLER_62_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17703_ _16973_/A _17346_/X _16973_/A _17346_/X VGND VGND VPWR VPWR _17703_/X sky130_fd_sc_hd__a2bb2o_4
X_14915_ _12529_/A _14911_/X _14914_/X VGND VGND VPWR VPWR _14916_/B sky130_fd_sc_hd__or3_4
XFILLER_7_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17405__B2 _17404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18683_ _16931_/X _18680_/Y _16933_/A _18682_/X VGND VGND VPWR VPWR _18683_/X sky130_fd_sc_hd__o22a_4
XFILLER_76_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15895_ _13554_/A _15839_/B VGND VGND VPWR VPWR _15895_/X sky130_fd_sc_hd__or2_4
XFILLER_110_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14829__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17634_ _18240_/A VGND VGND VPWR VPWR _17634_/X sky130_fd_sc_hd__buf_2
XANTENNA__13733__A _15494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14846_ _12599_/A _14846_/B _14846_/C VGND VGND VPWR VPWR _14846_/X sky130_fd_sc_hd__and3_4
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17565_ _17564_/X VGND VGND VPWR VPWR _17565_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14777_ _13960_/A _14777_/B VGND VGND VPWR VPWR _14778_/C sky130_fd_sc_hd__or2_4
X_11989_ _11936_/X _11989_/B _11989_/C VGND VGND VPWR VPWR _11990_/B sky130_fd_sc_hd__or3_4
XFILLER_75_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23117__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12349__A _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19304_ _16937_/X _17044_/Y _17640_/X _17770_/X VGND VGND VPWR VPWR _19304_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22701__A2 _22700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16516_ _16444_/Y _16513_/X VGND VGND VPWR VPWR _16516_/X sky130_fd_sc_hd__or2_4
XANTENNA__19420__A _16996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13728_ _12605_/A VGND VGND VPWR VPWR _15497_/A sky130_fd_sc_hd__buf_2
X_17496_ _16231_/A _17364_/X _17365_/X VGND VGND VPWR VPWR _17497_/B sky130_fd_sc_hd__o21a_4
XANTENNA__20712__B2 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16763__B _23931_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19235_ _19235_/A VGND VGND VPWR VPWR _19235_/Y sky130_fd_sc_hd__inv_2
X_16447_ _16447_/A _16445_/X _16447_/C VGND VGND VPWR VPWR _16447_/X sky130_fd_sc_hd__and3_4
X_13659_ _13659_/A VGND VGND VPWR VPWR _15429_/A sky130_fd_sc_hd__buf_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14564__A _14563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19166_ _24305_/Q _19167_/A _19165_/Y VGND VGND VPWR VPWR _24305_/D sky130_fd_sc_hd__o21a_4
X_16378_ _16377_/X VGND VGND VPWR VPWR _16378_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14283__B _14283_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18117_ _17969_/X _18116_/X _17254_/X VGND VGND VPWR VPWR _18117_/X sky130_fd_sc_hd__o21a_4
X_15329_ _15325_/X _15329_/B _15329_/C VGND VGND VPWR VPWR _15329_/X sky130_fd_sc_hd__and3_4
X_19097_ _11505_/A _11504_/Y _11506_/Y VGND VGND VPWR VPWR _19097_/X sky130_fd_sc_hd__o21a_4
X_18048_ _18048_/A VGND VGND VPWR VPWR _18048_/X sky130_fd_sc_hd__buf_2
XFILLER_82_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15395__A _13614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13908__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20010_ _20010_/A VGND VGND VPWR VPWR _20010_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19999_ _19999_/A VGND VGND VPWR VPWR _19999_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19397__B2 _24203_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21961_ _21855_/X _21959_/X _14743_/B _21956_/X VGND VGND VPWR VPWR _23523_/D sky130_fd_sc_hd__o22a_4
XFILLER_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22021__A _22020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23700_ _24084_/CLK _23700_/D VGND VGND VPWR VPWR _12827_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13643__A _13643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20912_ _24227_/Q _20444_/A _20911_/X VGND VGND VPWR VPWR _20912_/X sky130_fd_sc_hd__o21a_4
XFILLER_27_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17115__A _15185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21892_ _21823_/X _21887_/X _23568_/Q _21891_/X VGND VGND VPWR VPWR _21892_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22956__A _23015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _20846_/B VGND VGND VPWR VPWR _20844_/A sky130_fd_sc_hd__buf_2
X_23631_ _23987_/CLK _23631_/D VGND VGND VPWR VPWR _13569_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12259__A _12728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20774_ _20640_/X _20756_/X _20757_/X _20773_/Y VGND VGND VPWR VPWR _20774_/X sky130_fd_sc_hd__a211o_4
X_23562_ _23819_/CLK _23562_/D VGND VGND VPWR VPWR _23562_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17769__B _17263_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18372__A2 _18274_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22513_ _22462_/X _22486_/A _23199_/Q _22476_/A VGND VGND VPWR VPWR _22513_/X sky130_fd_sc_hd__o22a_4
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23493_ _23557_/CLK _23493_/D VGND VGND VPWR VPWR _14497_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14474__A _12494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24346__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22444_ _22129_/A VGND VGND VPWR VPWR _22444_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24192__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17785__A _18206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22375_ _22368_/A VGND VGND VPWR VPWR _22375_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21326_ _21319_/A VGND VGND VPWR VPWR _21326_/X sky130_fd_sc_hd__buf_2
X_24114_ _24202_/CLK _24114_/D HRESETn VGND VGND VPWR VPWR _22907_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__14921__B _14857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21100__A _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21257_ _21256_/X _21247_/X _13453_/B _21254_/X VGND VGND VPWR VPWR _23919_/D sky130_fd_sc_hd__o22a_4
X_24045_ _23922_/CLK _21039_/X VGND VGND VPWR VPWR _15818_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13818__A _13630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12722__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20208_ _20421_/A VGND VGND VPWR VPWR _20444_/A sky130_fd_sc_hd__buf_2
XANTENNA__21431__A2 _21426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21188_ _20591_/X _21183_/X _23952_/Q _21187_/X VGND VGND VPWR VPWR _21188_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20139_ _24428_/Q VGND VGND VPWR VPWR _20139_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19505__A _19598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23027__A _23027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12961_ _12949_/A _23603_/Q VGND VGND VPWR VPWR _12963_/B sky130_fd_sc_hd__or2_4
XFILLER_115_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14649__A _15203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21195__B2 _21194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14700_ _14673_/A _14700_/B _14699_/X VGND VGND VPWR VPWR _14700_/X sky130_fd_sc_hd__and3_4
XANTENNA__13553__A _12981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11912_ _11912_/A VGND VGND VPWR VPWR _12464_/A sky130_fd_sc_hd__buf_2
XFILLER_18_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18060__A1 _18011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15680_ _15812_/A _15679_/X VGND VGND VPWR VPWR _15680_/X sky130_fd_sc_hd__and2_4
XFILLER_59_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_15_0_HCLK_A clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12892_ _12892_/A _12892_/B VGND VGND VPWR VPWR _12892_/X sky130_fd_sc_hd__and2_4
XFILLER_79_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14368__B _14292_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14631_ _15006_/A _14703_/B VGND VGND VPWR VPWR _14631_/X sky130_fd_sc_hd__or2_4
X_11843_ _11842_/X VGND VGND VPWR VPWR _11843_/X sky130_fd_sc_hd__buf_2
X_23829_ _23315_/CLK _21417_/X VGND VGND VPWR VPWR _12648_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12169__A _12169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17350_ _15648_/X _17348_/B VGND VGND VPWR VPWR _18466_/B sky130_fd_sc_hd__and2_4
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14562_ _11799_/A _14546_/X _14561_/X VGND VGND VPWR VPWR _14563_/C sky130_fd_sc_hd__or3_4
X_11774_ _11774_/A _23934_/Q VGND VGND VPWR VPWR _11776_/B sky130_fd_sc_hd__or2_4
XANTENNA__17679__B _17487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22695__B2 _22690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16301_ _11982_/A _16278_/X _16285_/X _16292_/X _16300_/X VGND VGND VPWR VPWR _16301_/X
+ sky130_fd_sc_hd__a32o_4
X_13513_ _13558_/A _13513_/B VGND VGND VPWR VPWR _13516_/B sky130_fd_sc_hd__or2_4
X_17281_ _17278_/X _17280_/Y VGND VGND VPWR VPWR _17282_/A sky130_fd_sc_hd__or2_4
XFILLER_35_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14493_ _14492_/X VGND VGND VPWR VPWR _14493_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19020_ _19018_/Y _19019_/Y _11521_/B VGND VGND VPWR VPWR _19020_/X sky130_fd_sc_hd__o21a_4
X_16232_ _11658_/X _16232_/B _16232_/C VGND VGND VPWR VPWR _16233_/A sky130_fd_sc_hd__and3_4
XANTENNA__11801__A _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13444_ _12520_/X VGND VGND VPWR VPWR _13450_/A sky130_fd_sc_hd__buf_2
XFILLER_70_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16163_ _13395_/X VGND VGND VPWR VPWR _16201_/A sky130_fd_sc_hd__buf_2
X_13375_ _12837_/A VGND VGND VPWR VPWR _13399_/A sky130_fd_sc_hd__buf_2
X_15114_ _15114_/A _15112_/X _15113_/X VGND VGND VPWR VPWR _15115_/C sky130_fd_sc_hd__and3_4
X_12326_ _13317_/A _12317_/X _12325_/X VGND VGND VPWR VPWR _12326_/X sky130_fd_sc_hd__or3_4
XFILLER_86_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16094_ _16140_/A _16094_/B _16094_/C VGND VGND VPWR VPWR _16095_/C sky130_fd_sc_hd__and3_4
XFILLER_5_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21670__A2 _21669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15045_ _15045_/A _15045_/B _15045_/C VGND VGND VPWR VPWR _15046_/C sky130_fd_sc_hd__and3_4
X_19922_ _19916_/X _24143_/Q _19917_/X _20576_/B VGND VGND VPWR VPWR _24143_/D sky130_fd_sc_hd__o22a_4
XFILLER_79_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13728__A _12605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12257_ _12257_/A VGND VGND VPWR VPWR _12742_/A sky130_fd_sc_hd__buf_2
XANTENNA__16104__A _16109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21945__A _21938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12188_ _12116_/Y _12184_/X _12187_/X VGND VGND VPWR VPWR _12188_/Y sky130_fd_sc_hd__o21ai_4
X_19853_ _19872_/C _19851_/X _19852_/X _19672_/C _19622_/A VGND VGND VPWR VPWR _19853_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21422__A2 _21419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18804_ _14564_/X _18802_/X _20855_/A _18803_/X VGND VGND VPWR VPWR _24421_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15943__A _11933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16996_ _16996_/A VGND VGND VPWR VPWR _16997_/A sky130_fd_sc_hd__inv_2
X_19784_ _19454_/A _19784_/B VGND VGND VPWR VPWR _19784_/X sky130_fd_sc_hd__or2_4
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15947_ _13442_/X VGND VGND VPWR VPWR _15948_/A sky130_fd_sc_hd__buf_2
X_18735_ _18424_/X _18726_/Y _17854_/X _18734_/Y VGND VGND VPWR VPWR _18735_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15662__B _15724_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14559__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21186__B2 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24065__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13463__A _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18666_ _18202_/A _18664_/X _16935_/A _18665_/X VGND VGND VPWR VPWR _18666_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18051__B2 _18050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15878_ _12413_/X _15876_/X _15877_/X VGND VGND VPWR VPWR _15878_/X sky130_fd_sc_hd__and3_4
XFILLER_37_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14278__B _14278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14829_ _14841_/A _14765_/B VGND VGND VPWR VPWR _14829_/X sky130_fd_sc_hd__or2_4
X_17617_ _17321_/Y _17616_/X _17307_/Y VGND VGND VPWR VPWR _18578_/A sky130_fd_sc_hd__and3_4
X_18597_ _16960_/A _22913_/B _16969_/B VGND VGND VPWR VPWR _22921_/B sky130_fd_sc_hd__o21a_4
XFILLER_75_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17548_ _17547_/X VGND VGND VPWR VPWR _17550_/A sky130_fd_sc_hd__inv_2
XANTENNA__21489__A2 _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16493__B _16424_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17479_ _17506_/A _17479_/B VGND VGND VPWR VPWR _17479_/X sky130_fd_sc_hd__or2_4
XANTENNA__14294__A _15448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12807__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20161__A2 IRQ[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19218_ _19218_/A _19218_/B VGND VGND VPWR VPWR _19219_/B sky130_fd_sc_hd__and2_4
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20490_ _20342_/A _20490_/B VGND VGND VPWR VPWR _20490_/X sky130_fd_sc_hd__and2_4
XANTENNA__22438__B2 _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19149_ _19134_/X VGND VGND VPWR VPWR _19149_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22160_ _22079_/X _22158_/X _16658_/B _22155_/X VGND VGND VPWR VPWR _23420_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21661__A2 _21655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21111_ _21583_/A VGND VGND VPWR VPWR _21348_/C sky130_fd_sc_hd__buf_2
XANTENNA__13638__A _15412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22091_ _20441_/A VGND VGND VPWR VPWR _22091_/X sky130_fd_sc_hd__buf_2
XANTENNA__12542__A _12497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21042_ _20723_/X _21037_/X _15556_/B _21041_/X VGND VGND VPWR VPWR _21042_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21413__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22610__B2 _22604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15853__A _12386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19325__A _19328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22993_ _18283_/X _23004_/B VGND VGND VPWR VPWR _22994_/C sky130_fd_sc_hd__or2_4
XANTENNA__21177__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21944_ _21826_/X _21938_/X _23535_/Q _21942_/X VGND VGND VPWR VPWR _23535_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22686__A _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21590__A _21590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23432__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21875_ _21795_/X _21873_/X _23580_/Q _21870_/X VGND VGND VPWR VPWR _23580_/D sky130_fd_sc_hd__o22a_4
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20918__B _20539_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23320_/CLK _21790_/X VGND VGND VPWR VPWR _23614_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _24390_/Q _20623_/X _24422_/Q _20682_/X VGND VGND VPWR VPWR _20826_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22677__A1 _21799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22677__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23545_ _23514_/CLK _21930_/X VGND VGND VPWR VPWR _16260_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20757_ _20515_/A VGND VGND VPWR VPWR _20757_/X sky130_fd_sc_hd__buf_2
XFILLER_51_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12717__A _12709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22429__B2 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20688_ _20493_/X _20687_/X _19121_/A _20500_/X VGND VGND VPWR VPWR _20689_/B sky130_fd_sc_hd__o22a_4
X_23476_ _23539_/CLK _23476_/D VGND VGND VPWR VPWR _12735_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22427_ _22112_/A VGND VGND VPWR VPWR _22427_/X sky130_fd_sc_hd__buf_2
XFILLER_87_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21101__B2 _21100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13160_ _12737_/A _13157_/X _13159_/X VGND VGND VPWR VPWR _13160_/X sky130_fd_sc_hd__and3_4
XFILLER_100_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22358_ _22351_/A VGND VGND VPWR VPWR _22358_/X sky130_fd_sc_hd__buf_2
X_12111_ _11966_/X _12111_/B _12110_/X VGND VGND VPWR VPWR _12112_/C sky130_fd_sc_hd__and3_4
XANTENNA__19771__A2_N _19769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13091_ _13115_/A _13091_/B VGND VGND VPWR VPWR _13092_/C sky130_fd_sc_hd__or2_4
X_21309_ _21301_/X VGND VGND VPWR VPWR _21309_/X sky130_fd_sc_hd__buf_2
XFILLER_108_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13548__A _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22289_ _22129_/X _22286_/X _23335_/Q _22283_/X VGND VGND VPWR VPWR _23335_/D sky130_fd_sc_hd__o22a_4
XFILLER_46_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12042_ _16714_/A _23517_/Q VGND VGND VPWR VPWR _12043_/C sky130_fd_sc_hd__or2_4
X_24028_ _23515_/CLK _24028_/D VGND VGND VPWR VPWR _24028_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22601__B2 _22597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12171__B _23869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16850_ _16850_/A _16850_/B VGND VGND VPWR VPWR _16850_/X sky130_fd_sc_hd__or2_4
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15801_ _12868_/A _23309_/Q VGND VGND VPWR VPWR _15803_/B sky130_fd_sc_hd__or2_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16781_ _16629_/X _23899_/Q VGND VGND VPWR VPWR _16783_/B sky130_fd_sc_hd__or2_4
X_13993_ _12598_/A VGND VGND VPWR VPWR _14050_/A sky130_fd_sc_hd__buf_2
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18520_ _17422_/D _18519_/X VGND VGND VPWR VPWR _18520_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__13283__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15732_ _12792_/A _15732_/B VGND VGND VPWR VPWR _15732_/X sky130_fd_sc_hd__or2_4
X_12944_ _12982_/A _12942_/X _12943_/X VGND VGND VPWR VPWR _12948_/B sky130_fd_sc_hd__and3_4
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18451_ _17382_/B _18450_/X VGND VGND VPWR VPWR _18451_/X sky130_fd_sc_hd__or2_4
X_15663_ _12726_/A _15725_/B VGND VGND VPWR VPWR _15663_/X sky130_fd_sc_hd__or2_4
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12875_ _12910_/A _12875_/B _12875_/C VGND VGND VPWR VPWR _12876_/C sky130_fd_sc_hd__and3_4
XANTENNA__16595__A1 _11844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17402_ _20197_/B _11634_/X _11886_/X _17034_/Y VGND VGND VPWR VPWR _17402_/X sky130_fd_sc_hd__a2bb2o_4
X_14614_ _14725_/A _14695_/B VGND VGND VPWR VPWR _14614_/X sky130_fd_sc_hd__or2_4
X_11826_ _11754_/X VGND VGND VPWR VPWR _11827_/A sky130_fd_sc_hd__buf_2
X_18382_ _18291_/X _18379_/X _20029_/A _18381_/X VGND VGND VPWR VPWR _24463_/D sky130_fd_sc_hd__a2bb2o_4
X_15594_ _15618_/A _23275_/Q VGND VGND VPWR VPWR _15594_/X sky130_fd_sc_hd__or2_4
XFILLER_72_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17333_ _15251_/X _17227_/A _17327_/X _17332_/X VGND VGND VPWR VPWR _17333_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _13754_/A _14541_/X _14544_/X VGND VGND VPWR VPWR _14546_/C sky130_fd_sc_hd__or3_4
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _16025_/A VGND VGND VPWR VPWR _16069_/A sky130_fd_sc_hd__buf_2
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15003__A _14588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17264_ _16596_/Y _17016_/X _17023_/X _17263_/Y VGND VGND VPWR VPWR _17264_/X sky130_fd_sc_hd__o22a_4
X_14476_ _13022_/A _14476_/B VGND VGND VPWR VPWR _14476_/X sky130_fd_sc_hd__or2_4
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11688_ _15774_/A VGND VGND VPWR VPWR _12837_/A sky130_fd_sc_hd__buf_2
X_19003_ _24338_/Q _11522_/X _18996_/Y VGND VGND VPWR VPWR _19003_/Y sky130_fd_sc_hd__a21oi_4
X_16215_ _16215_/A _16215_/B _16215_/C VGND VGND VPWR VPWR _16231_/B sky130_fd_sc_hd__and3_4
X_13427_ _13427_/A _13427_/B VGND VGND VPWR VPWR _13427_/X sky130_fd_sc_hd__or2_4
XANTENNA__15938__A _15937_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17195_ _17194_/X VGND VGND VPWR VPWR _17195_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18314__A _18171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16146_ _16146_/A _16217_/B VGND VGND VPWR VPWR _16147_/C sky130_fd_sc_hd__or2_4
X_13358_ _12827_/A VGND VGND VPWR VPWR _13358_/X sky130_fd_sc_hd__buf_2
XANTENNA__21643__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12309_ _13678_/A VGND VGND VPWR VPWR _15552_/A sky130_fd_sc_hd__buf_2
XANTENNA__13458__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16077_ _16077_/A _16077_/B _16077_/C VGND VGND VPWR VPWR _16077_/X sky130_fd_sc_hd__and3_4
X_13289_ _12540_/A _13287_/X _13289_/C VGND VGND VPWR VPWR _13289_/X sky130_fd_sc_hd__and3_4
XANTENNA__23305__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15028_ _15028_/A _15028_/B _15028_/C VGND VGND VPWR VPWR _15032_/B sky130_fd_sc_hd__and3_4
X_19905_ _19899_/X _24156_/Q _19903_/X _20650_/A VGND VGND VPWR VPWR _24156_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15673__A _12235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19836_ _19637_/A _19834_/X _19703_/A _19835_/X VGND VGND VPWR VPWR _19836_/X sky130_fd_sc_hd__o22a_4
XFILLER_96_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15392__B _15454_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19767_ _19429_/A _19764_/X _19612_/A _19766_/X VGND VGND VPWR VPWR _19767_/X sky130_fd_sc_hd__a211o_4
XFILLER_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16979_ _17673_/A _16979_/B VGND VGND VPWR VPWR _16980_/B sky130_fd_sc_hd__or2_4
XANTENNA__14289__A _15556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21159__B2 _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13193__A _12745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18718_ _18718_/A VGND VGND VPWR VPWR _18718_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20367__C1 _20366_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19698_ _19549_/X _19682_/X _19696_/X _12036_/X _19697_/X VGND VGND VPWR VPWR _24181_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19772__A1 _19873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18649_ _16927_/A _18646_/X _17639_/A _18648_/X VGND VGND VPWR VPWR _18649_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13921__A _13837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21660_ _21538_/X _21655_/X _23696_/Q _21659_/X VGND VGND VPWR VPWR _23696_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22659__B2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20611_ _21256_/A VGND VGND VPWR VPWR _20611_/X sky130_fd_sc_hd__buf_2
X_21591_ _21605_/A VGND VGND VPWR VPWR _21591_/X sky130_fd_sc_hd__buf_2
XANTENNA__12537__A _12466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21331__B2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20542_ _20448_/X _20541_/X _24370_/Q _20407_/X VGND VGND VPWR VPWR _20542_/X sky130_fd_sc_hd__o22a_4
X_23330_ _23522_/CLK _23330_/D VGND VGND VPWR VPWR _15255_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20754__A _20754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20473_ _20473_/A VGND VGND VPWR VPWR _20473_/X sky130_fd_sc_hd__buf_2
X_23261_ _24059_/CLK _23261_/D VGND VGND VPWR VPWR _12118_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15848__A _13546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14752__A _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18224__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22212_ _22212_/A VGND VGND VPWR VPWR _22212_/X sky130_fd_sc_hd__buf_2
X_23192_ _23130_/CLK _23192_/D VGND VGND VPWR VPWR _16019_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_88_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15567__B _24075_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20192__C _21583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22143_ _22458_/A VGND VGND VPWR VPWR _22143_/X sky130_fd_sc_hd__buf_2
XANTENNA__12272__A _13054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22074_ _22066_/Y _22072_/X _22073_/X _22072_/X VGND VGND VPWR VPWR _23454_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16679__A _16596_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22595__B1 _15863_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21025_ _20442_/X _21023_/X _24055_/Q _21020_/X VGND VGND VPWR VPWR _24055_/D sky130_fd_sc_hd__o22a_4
XFILLER_113_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_1_0_HCLK_A clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16398__B _16398_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22976_ _22955_/X _17893_/X _22967_/X _22975_/X VGND VGND VPWR VPWR _22977_/A sky130_fd_sc_hd__a211o_4
XFILLER_28_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19763__A1 _20576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21927_ _21797_/X _21924_/X _23547_/Q _21921_/X VGND VGND VPWR VPWR _23547_/D sky130_fd_sc_hd__o22a_4
XFILLER_76_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17303__A _17297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12660_ _12660_/A _12660_/B VGND VGND VPWR VPWR _12662_/B sky130_fd_sc_hd__or2_4
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _21857_/X _21853_/X _15285_/B _21848_/X VGND VGND VPWR VPWR _23586_/D sky130_fd_sc_hd__o22a_4
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11611_/A VGND VGND VPWR VPWR _13966_/A sky130_fd_sc_hd__buf_2
XFILLER_19_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20760_/X _20808_/X _19065_/A _20767_/X VGND VGND VPWR VPWR _20809_/X sky130_fd_sc_hd__o22a_4
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12935_/A VGND VGND VPWR VPWR _12591_/X sky130_fd_sc_hd__buf_2
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21789_ _21789_/A VGND VGND VPWR VPWR _21789_/X sky130_fd_sc_hd__buf_2
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21322__B2 _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _15576_/A _14330_/B VGND VGND VPWR VPWR _14332_/B sky130_fd_sc_hd__or2_4
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _24418_/Q IRQ[3] _11541_/Y VGND VGND VPWR VPWR _11542_/X sky130_fd_sc_hd__a21bo_4
X_23528_ _23304_/CLK _21954_/X VGND VGND VPWR VPWR _13636_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_11_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _14073_/A _14261_/B _14260_/X VGND VGND VPWR VPWR _14261_/X sky130_fd_sc_hd__and3_4
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23459_ _23270_/CLK _22061_/X VGND VGND VPWR VPWR _14769_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18134__A _18062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16000_ _15999_/X _23704_/Q VGND VGND VPWR VPWR _16003_/B sky130_fd_sc_hd__or2_4
XFILLER_32_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13212_ _12791_/A _13144_/B VGND VGND VPWR VPWR _13214_/B sky130_fd_sc_hd__or2_4
XANTENNA__22822__A1 _15713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21625__A2 _21619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14192_ _13709_/A VGND VGND VPWR VPWR _14195_/A sky130_fd_sc_hd__buf_2
XFILLER_67_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17829__B2 _17828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13143_ _12706_/A _13139_/X _13142_/X VGND VGND VPWR VPWR _13143_/X sky130_fd_sc_hd__or3_4
XFILLER_83_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12182__A _16677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13074_ _13104_/A _13005_/B VGND VGND VPWR VPWR _13074_/X sky130_fd_sc_hd__or2_4
X_17951_ _17951_/A _17894_/X VGND VGND VPWR VPWR _17951_/X sky130_fd_sc_hd__and2_4
XANTENNA__23478__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21389__B2 _21387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12025_ _12025_/A _12025_/B _12025_/C VGND VGND VPWR VPWR _12026_/C sky130_fd_sc_hd__and3_4
X_16902_ _16902_/A VGND VGND VPWR VPWR _16903_/D sky130_fd_sc_hd__inv_2
X_17882_ _17641_/X VGND VGND VPWR VPWR _17882_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22050__A2 _22045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_30_0_HCLK_A clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19621_ _19621_/A VGND VGND VPWR VPWR _19622_/A sky130_fd_sc_hd__buf_2
XFILLER_4_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16833_ _13280_/B _16832_/X _13272_/X VGND VGND VPWR VPWR _16833_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_111_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16764_ _16773_/A _23579_/Q VGND VGND VPWR VPWR _16765_/C sky130_fd_sc_hd__or2_4
X_19552_ _19416_/B VGND VGND VPWR VPWR _19553_/A sky130_fd_sc_hd__buf_2
X_13976_ _12202_/A _14066_/B VGND VGND VPWR VPWR _13978_/B sky130_fd_sc_hd__or2_4
XFILLER_59_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20839__A _20488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15715_ _13130_/A _15715_/B VGND VGND VPWR VPWR _15715_/X sky130_fd_sc_hd__or2_4
X_18503_ _18697_/A _17409_/A VGND VGND VPWR VPWR _18503_/X sky130_fd_sc_hd__and2_4
X_12927_ _12967_/A _12925_/X _12926_/X VGND VGND VPWR VPWR _12927_/X sky130_fd_sc_hd__and3_4
X_16695_ _16718_/A _16695_/B _16695_/C VGND VGND VPWR VPWR _16696_/C sky130_fd_sc_hd__and3_4
X_19483_ _19538_/A _19541_/A VGND VGND VPWR VPWR _19483_/X sky130_fd_sc_hd__or2_4
XANTENNA__14837__A _14021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21561__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13741__A _11648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15646_ _15645_/X VGND VGND VPWR VPWR _15646_/X sky130_fd_sc_hd__buf_2
X_18434_ _18381_/X _18433_/X _24461_/Q _18381_/X VGND VGND VPWR VPWR _18434_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12858_ _12895_/A _12858_/B VGND VGND VPWR VPWR _12859_/C sky130_fd_sc_hd__or2_4
X_11809_ _11747_/X _11805_/X _11809_/C VGND VGND VPWR VPWR _11817_/B sky130_fd_sc_hd__or3_4
X_18365_ _17969_/X _18111_/X _17866_/X VGND VGND VPWR VPWR _18365_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15577_ _15393_/A _15577_/B VGND VGND VPWR VPWR _15578_/C sky130_fd_sc_hd__or2_4
X_12789_ _12800_/A _23572_/Q VGND VGND VPWR VPWR _12790_/C sky130_fd_sc_hd__or2_4
XANTENNA__12357__A _15743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21313__B2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17316_ _18583_/B _17311_/X _17618_/C VGND VGND VPWR VPWR _17316_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_33_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14528_ _13711_/X _14528_/B _14527_/X VGND VGND VPWR VPWR _14529_/C sky130_fd_sc_hd__and3_4
X_18296_ _18242_/A _17510_/X VGND VGND VPWR VPWR _18298_/C sky130_fd_sc_hd__nor2_4
XANTENNA__21864__A2 _21817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20574__A _20574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18190__B1 _18189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17247_ _17246_/X VGND VGND VPWR VPWR _17247_/Y sky130_fd_sc_hd__inv_2
X_14459_ _12459_/A _14455_/X _14459_/C VGND VGND VPWR VPWR _14460_/B sky130_fd_sc_hd__or3_4
XANTENNA__14572__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17178_ _13772_/X VGND VGND VPWR VPWR _17178_/X sky130_fd_sc_hd__buf_2
X_16129_ _16109_/A _16129_/B _16129_/C VGND VGND VPWR VPWR _16130_/C sky130_fd_sc_hd__and3_4
XANTENNA__13188__A _15784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18493__A1 _18142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22577__B1 _16407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13916__A _11670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22041__A2 _22038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12820__A _12769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19819_ _19640_/B _19846_/B _19669_/Y VGND VGND VPWR VPWR _19819_/X sky130_fd_sc_hd__o21a_4
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22830_ _22830_/A VGND VGND VPWR VPWR HWDATA[16] sky130_fd_sc_hd__inv_2
XFILLER_42_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19603__A _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_55_0_HCLK clkbuf_7_54_0_HCLK/A VGND VGND VPWR VPWR _24044_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22761_ _22759_/Y _22763_/B _22754_/X VGND VGND VPWR VPWR _24099_/D sky130_fd_sc_hd__and3_4
XFILLER_53_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14747__A _15037_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21552__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13651__A _13651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21712_ _21705_/A VGND VGND VPWR VPWR _21712_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22692_ _21256_/A _22686_/X _13484_/B _22690_/X VGND VGND VPWR VPWR _22692_/X sky130_fd_sc_hd__o22a_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ _24334_/CLK _24431_/D HRESETn VGND VGND VPWR VPWR _24431_/Q sky130_fd_sc_hd__dfrtp_4
X_21643_ _21510_/X _21641_/X _23708_/Q _21638_/X VGND VGND VPWR VPWR _23708_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20107__A2 _20106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24362_ _24330_/CLK _18907_/X HRESETn VGND VGND VPWR VPWR _24362_/Q sky130_fd_sc_hd__dfstp_4
X_21574_ _21574_/A VGND VGND VPWR VPWR _21574_/X sky130_fd_sc_hd__buf_2
XANTENNA__20484__A _20484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23313_ _23313_/CLK _22313_/X VGND VGND VPWR VPWR _13157_/B sky130_fd_sc_hd__dfxtp_4
X_20525_ _20525_/A VGND VGND VPWR VPWR _20525_/X sky130_fd_sc_hd__buf_2
X_24293_ _24293_/CLK _24293_/D HRESETn VGND VGND VPWR VPWR _19114_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14482__A _13025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20456_ _20502_/A _20455_/X VGND VGND VPWR VPWR _20456_/Y sky130_fd_sc_hd__nor2_4
X_23244_ _23404_/CLK _23244_/D VGND VGND VPWR VPWR _15454_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_107_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21607__A2 _21605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20815__B1 _20814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17793__A _18082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20387_ _18050_/X _20578_/A _20290_/X _20386_/Y VGND VGND VPWR VPWR _20387_/X sky130_fd_sc_hd__a211o_4
X_23175_ _23557_/CLK _23175_/D VGND VGND VPWR VPWR _13784_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22280__A2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22126_ _22124_/X _22125_/X _23433_/Q _22120_/X VGND VGND VPWR VPWR _23433_/D sky130_fd_sc_hd__o22a_4
XFILLER_0_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22204__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13826__A _13631_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22057_ _21847_/X _22052_/X _14317_/B _22056_/X VGND VGND VPWR VPWR _22057_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12730__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21008_ _21008_/A VGND VGND VPWR VPWR _21734_/B sky130_fd_sc_hd__buf_2
XFILLER_101_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17995__B1 _17874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20594__A2 _19770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13830_ _13677_/A _13828_/X _13830_/C VGND VGND VPWR VPWR _13830_/X sky130_fd_sc_hd__and3_4
XFILLER_63_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13761_ _13737_/A _13759_/X _13760_/X VGND VGND VPWR VPWR _13761_/X sky130_fd_sc_hd__and3_4
X_22959_ _22982_/A _22957_/Y _22958_/X VGND VGND VPWR VPWR _22959_/X sky130_fd_sc_hd__and3_4
XFILLER_95_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14657__A _11738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15500_ _12612_/A _15492_/X _15500_/C VGND VGND VPWR VPWR _15516_/B sky130_fd_sc_hd__and3_4
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18129__A _18129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12712_ _12198_/X _12710_/X _12711_/X VGND VGND VPWR VPWR _12712_/X sky130_fd_sc_hd__and3_4
X_16480_ _11770_/X _16480_/B _16479_/X VGND VGND VPWR VPWR _16481_/C sky130_fd_sc_hd__and3_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13692_ _14178_/A VGND VGND VPWR VPWR _14010_/A sky130_fd_sc_hd__buf_2
XFILLER_43_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15431_ _15431_/A _15429_/X _15431_/C VGND VGND VPWR VPWR _15435_/B sky130_fd_sc_hd__and3_4
X_12643_ _12643_/A _12643_/B VGND VGND VPWR VPWR _12644_/C sky130_fd_sc_hd__or2_4
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17968__A _18142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22099__A2 _22089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ _17447_/X _17455_/X _18217_/B VGND VGND VPWR VPWR _18151_/B sky130_fd_sc_hd__or3_4
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15362_ _14020_/A _15362_/B _15361_/X VGND VGND VPWR VPWR _15362_/X sky130_fd_sc_hd__and3_4
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12574_ _14009_/A VGND VGND VPWR VPWR _12575_/A sky130_fd_sc_hd__buf_2
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21846__A2 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20503__C1 _20502_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20394__A _21802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17101_ _17100_/X VGND VGND VPWR VPWR _17101_/X sky130_fd_sc_hd__buf_2
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ _11911_/A _14313_/B _14312_/X VGND VGND VPWR VPWR _14313_/X sky130_fd_sc_hd__and3_4
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ _24340_/Q _11524_/X VGND VGND VPWR VPWR _11525_/X sky130_fd_sc_hd__or2_4
X_18081_ _18081_/A _18081_/B VGND VGND VPWR VPWR _18081_/X sky130_fd_sc_hd__or2_4
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15293_ _14161_/A _15293_/B VGND VGND VPWR VPWR _15293_/X sky130_fd_sc_hd__or2_4
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14392__A _15592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12905__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17032_ _17105_/A _17032_/B VGND VGND VPWR VPWR _17032_/X sky130_fd_sc_hd__and2_4
X_14244_ _14204_/A _23081_/Q VGND VGND VPWR VPWR _14244_/X sky130_fd_sc_hd__or2_4
XFILLER_67_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14175_ _14175_/A VGND VGND VPWR VPWR _14202_/A sky130_fd_sc_hd__buf_2
XANTENNA__22271__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13126_ _13098_/A _23474_/Q VGND VGND VPWR VPWR _13126_/X sky130_fd_sc_hd__or2_4
XFILLER_113_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18983_ _11525_/X VGND VGND VPWR VPWR _18983_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13736__A _12652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13057_ _12892_/A _13034_/X _13041_/X _13048_/X _13056_/X VGND VGND VPWR VPWR _13057_/X
+ sky130_fd_sc_hd__a32o_4
X_17934_ _17801_/X _17246_/X _17807_/X _17847_/X VGND VGND VPWR VPWR _17934_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__12640__A _12640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12008_ _12008_/A _23486_/Q VGND VGND VPWR VPWR _12011_/B sky130_fd_sc_hd__or2_4
XFILLER_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17865_ _17244_/X _17226_/Y _17252_/X VGND VGND VPWR VPWR _17865_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21782__B2 _21737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19604_ _19826_/B VGND VGND VPWR VPWR _19822_/A sky130_fd_sc_hd__buf_2
X_16816_ _16743_/X _16814_/B _16815_/Y VGND VGND VPWR VPWR _16816_/X sky130_fd_sc_hd__a21o_4
X_17796_ _17962_/A VGND VGND VPWR VPWR _17796_/X sky130_fd_sc_hd__buf_2
XFILLER_94_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19535_ _19535_/A VGND VGND VPWR VPWR _19536_/B sky130_fd_sc_hd__inv_2
X_13959_ _13959_/A _23882_/Q VGND VGND VPWR VPWR _13959_/X sky130_fd_sc_hd__or2_4
X_16747_ _11729_/X VGND VGND VPWR VPWR _16747_/X sky130_fd_sc_hd__buf_2
XFILLER_46_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13471__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16678_ _16077_/A _16646_/X _16677_/X VGND VGND VPWR VPWR _16678_/X sky130_fd_sc_hd__and3_4
X_19466_ _19458_/X _19465_/X HRDATA[11] _19462_/X VGND VGND VPWR VPWR _19517_/A sky130_fd_sc_hd__o22a_4
XFILLER_35_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20742__C1 _20741_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22784__A _15120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18417_ _18416_/X VGND VGND VPWR VPWR _18417_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15629_ _15617_/A _15573_/B VGND VGND VPWR VPWR _15629_/X sky130_fd_sc_hd__or2_4
XFILLER_37_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17878__A _18390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19397_ _19396_/X _18463_/Y _19396_/X _24203_/Q VGND VGND VPWR VPWR _24203_/D sky130_fd_sc_hd__a2bb2o_4
X_18348_ _18348_/A _18348_/B VGND VGND VPWR VPWR _18349_/B sky130_fd_sc_hd__or2_4
XANTENNA__21837__A2 _21829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15398__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18279_ _18307_/A _18278_/X _17519_/Y VGND VGND VPWR VPWR _18279_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_11_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20310_ _20284_/X _20287_/X _20288_/X _20309_/Y VGND VGND VPWR VPWR _20310_/X sky130_fd_sc_hd__a211o_4
XFILLER_50_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21290_ _21289_/X _21283_/X _15146_/B _21230_/A VGND VGND VPWR VPWR _23905_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20241_ _20447_/A VGND VGND VPWR VPWR _20270_/A sky130_fd_sc_hd__inv_2
XFILLER_85_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18502__A _18443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24107__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20172_ _20074_/Y _20172_/B VGND VGND VPWR VPWR _20173_/B sky130_fd_sc_hd__or2_4
XFILLER_66_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15845__B _15845_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22024__A _22031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17763__D _17762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22014__A2 _22009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12550__A _13031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23931_ _23931_/CLK _21228_/X VGND VGND VPWR VPWR _23931_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24149__CLK _24223_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15861__A _13548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23862_ _23473_/CLK _21365_/X VGND VGND VPWR VPWR _12332_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15452__A1 _13594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22813_ _22862_/A VGND VGND VPWR VPWR _22813_/X sky130_fd_sc_hd__buf_2
XFILLER_72_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23793_ _23342_/CLK _23793_/D VGND VGND VPWR VPWR _13254_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_22_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14477__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21525__B2 _21515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22722__B1 _23064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24299__CLK _24299_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22744_ _24101_/Q VGND VGND VPWR VPWR _22744_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17788__A _18066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22675_ _21797_/A _22672_/X _23099_/Q _22669_/X VGND VGND VPWR VPWR _23099_/D sky130_fd_sc_hd__o22a_4
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24414_ _24435_/CLK _24414_/D HRESETn VGND VGND VPWR VPWR _24414_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21626_ _21590_/A VGND VGND VPWR VPWR _21626_/X sky130_fd_sc_hd__buf_2
XANTENNA__21103__A _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24345_ _24344_/CLK _24345_/D HRESETn VGND VGND VPWR VPWR _11530_/A sky130_fd_sc_hd__dfstp_4
X_21557_ _21555_/X _21556_/X _23753_/Q _21551_/X VGND VGND VPWR VPWR _21557_/X sky130_fd_sc_hd__o22a_4
XFILLER_21_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12725__A _12725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15101__A _14055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20508_ _22413_/A VGND VGND VPWR VPWR _20509_/A sky130_fd_sc_hd__buf_2
X_12290_ _12726_/A _24054_/Q VGND VGND VPWR VPWR _12290_/X sky130_fd_sc_hd__or2_4
X_24276_ _23326_/CLK _24276_/D HRESETn VGND VGND VPWR VPWR _19225_/A sky130_fd_sc_hd__dfrtp_4
X_21488_ _21467_/A VGND VGND VPWR VPWR _21488_/X sky130_fd_sc_hd__buf_2
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12444__B _12571_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23227_ _24059_/CLK _23227_/D VGND VGND VPWR VPWR _16806_/B sky130_fd_sc_hd__dfxtp_4
X_20439_ _20484_/A _20438_/X VGND VGND VPWR VPWR _20439_/X sky130_fd_sc_hd__or2_4
XANTENNA__14940__A _15072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23158_ _23313_/CLK _22582_/X VGND VGND VPWR VPWR _12274_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15755__B _15690_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22109_ _22107_/X _22101_/X _13312_/B _22108_/X VGND VGND VPWR VPWR _23440_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13556__A _13494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15980_ _15980_/A _15976_/X _15980_/C VGND VGND VPWR VPWR _15980_/X sky130_fd_sc_hd__or3_4
XANTENNA__22005__A2 _22002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23089_ _23564_/CLK _22689_/X VGND VGND VPWR VPWR _13193_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12460__A _12460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20016__A1 _19994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14931_ _14002_/A VGND VGND VPWR VPWR _14937_/A sky130_fd_sc_hd__buf_2
XFILLER_94_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21773__A _21752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13275__B _13274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21764__B2 _21759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15771__A _12765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14862_ _13986_/A _14858_/X _14861_/X VGND VGND VPWR VPWR _14862_/X sky130_fd_sc_hd__or3_4
X_17650_ _24135_/Q _17544_/X _17647_/X VGND VGND VPWR VPWR _17651_/B sky130_fd_sc_hd__o21ai_4
XFILLER_36_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13813_ _13813_/A _13809_/X _13813_/C VGND VGND VPWR VPWR _13813_/X sky130_fd_sc_hd__or3_4
X_16601_ _12152_/A VGND VGND VPWR VPWR _16799_/A sky130_fd_sc_hd__buf_2
X_17581_ _18066_/B _17565_/Y _17556_/X VGND VGND VPWR VPWR _17581_/Y sky130_fd_sc_hd__o21ai_4
X_14793_ _14816_/A _14789_/X _14793_/C VGND VGND VPWR VPWR _14793_/X sky130_fd_sc_hd__or3_4
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14387__A _15611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21516__B2 _21515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22713__B1 _23071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16532_ _12011_/A _16530_/X _16532_/C VGND VGND VPWR VPWR _16533_/C sky130_fd_sc_hd__and3_4
X_19320_ _19318_/X _18054_/X _19318_/X _24249_/Q VGND VGND VPWR VPWR _24249_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13291__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11804__A _11717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13744_ _15493_/A _23592_/Q VGND VGND VPWR VPWR _13746_/B sky130_fd_sc_hd__or2_4
XFILLER_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17196__A1 _15909_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23666__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16463_ _11673_/X _16454_/X _16462_/X VGND VGND VPWR VPWR _16463_/X sky130_fd_sc_hd__and3_4
X_19251_ _19251_/A VGND VGND VPWR VPWR _19251_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13675_ _12203_/A _13756_/B VGND VGND VPWR VPWR _13675_/X sky130_fd_sc_hd__or2_4
X_15414_ _13641_/A _15471_/B VGND VGND VPWR VPWR _15415_/C sky130_fd_sc_hd__or2_4
X_18202_ _18202_/A VGND VGND VPWR VPWR _18202_/X sky130_fd_sc_hd__buf_2
X_12626_ _12626_/A VGND VGND VPWR VPWR _12955_/A sky130_fd_sc_hd__buf_2
X_19182_ _24297_/Q _19118_/B _19181_/Y VGND VGND VPWR VPWR _19182_/X sky130_fd_sc_hd__o21a_4
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16394_ _12546_/A VGND VGND VPWR VPWR _16394_/X sky130_fd_sc_hd__buf_2
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18133_ _23016_/B _18132_/X _23016_/B _18132_/X VGND VGND VPWR VPWR _18133_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15345_ _13992_/A _15345_/B _15344_/X VGND VGND VPWR VPWR _15345_/X sky130_fd_sc_hd__or3_4
XFILLER_34_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21013__A _21012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12557_ _12922_/A _12556_/X VGND VGND VPWR VPWR _12557_/X sky130_fd_sc_hd__and2_4
XANTENNA__18696__A1 _18499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12635__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22492__A2 _22486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11508_ _24323_/Q _11508_/B VGND VGND VPWR VPWR _11508_/X sky130_fd_sc_hd__or2_4
X_18064_ _18205_/A _17572_/B VGND VGND VPWR VPWR _18064_/X sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_4_4_0_HCLK_A clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15276_ _14588_/X _15276_/B VGND VGND VPWR VPWR _15276_/X sky130_fd_sc_hd__or2_4
XFILLER_32_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12488_ _13031_/A VGND VGND VPWR VPWR _12872_/A sky130_fd_sc_hd__buf_2
XFILLER_32_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17015_ _17014_/X VGND VGND VPWR VPWR _17015_/X sky130_fd_sc_hd__buf_2
XANTENNA__24271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14227_ _14195_/A _14227_/B _14227_/C VGND VGND VPWR VPWR _14233_/B sky130_fd_sc_hd__and3_4
XANTENNA__22244__A2 _22243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14850__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24200__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14158_ _14158_/A _23209_/Q VGND VGND VPWR VPWR _14162_/B sky130_fd_sc_hd__or2_4
XFILLER_113_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13109_ _13109_/A _13109_/B _13109_/C VGND VGND VPWR VPWR _13110_/C sky130_fd_sc_hd__and3_4
XFILLER_98_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14089_ _14089_/A _23753_/Q VGND VGND VPWR VPWR _14090_/C sky130_fd_sc_hd__or2_4
X_18966_ _24344_/Q _11528_/X _18959_/Y VGND VGND VPWR VPWR _18966_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__20007__A1 _19994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17917_ _17910_/X _17913_/Y _17914_/X _17916_/Y VGND VGND VPWR VPWR _17917_/X sky130_fd_sc_hd__o22a_4
XFILLER_26_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18897_ _17194_/X _18891_/X _24368_/Q _18892_/X VGND VGND VPWR VPWR _24368_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16777__A _16747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17848_ _17802_/X _17232_/X _17804_/X _17228_/X VGND VGND VPWR VPWR _17848_/X sky130_fd_sc_hd__o22a_4
XFILLER_94_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17779_ _18063_/A VGND VGND VPWR VPWR _17779_/X sky130_fd_sc_hd__buf_2
XANTENNA__14297__A _14322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19518_ _24147_/Q _19459_/X HRDATA[21] _19460_/X VGND VGND VPWR VPWR _19518_/X sky130_fd_sc_hd__o22a_4
X_20790_ _20630_/A _20790_/B VGND VGND VPWR VPWR _20790_/Y sky130_fd_sc_hd__nor2_4
XFILLER_23_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17187__A1 _15782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22180__B2 _22176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19449_ _19449_/A VGND VGND VPWR VPWR _19449_/X sky130_fd_sc_hd__buf_2
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17401__A _22017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22460_ _22460_/A VGND VGND VPWR VPWR _22460_/X sky130_fd_sc_hd__buf_2
XANTENNA__22019__A _22052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21411_ _21232_/X _21405_/X _16280_/B _21409_/X VGND VGND VPWR VPWR _23833_/D sky130_fd_sc_hd__o22a_4
X_22391_ _22384_/X VGND VGND VPWR VPWR _22416_/A sky130_fd_sc_hd__buf_2
XANTENNA__12545__A _12553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24130_ _23522_/CLK _20008_/Y HRESETn VGND VGND VPWR VPWR _24130_/Q sky130_fd_sc_hd__dfrtp_4
X_21342_ _21285_/X _21340_/X _14819_/B _21337_/X VGND VGND VPWR VPWR _21342_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14173__A1 _12267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24061_ _23485_/CLK _24061_/D VGND VGND VPWR VPWR _24061_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15856__A _13548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19328__A _19328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21273_ _21843_/A VGND VGND VPWR VPWR _21273_/X sky130_fd_sc_hd__buf_2
XANTENNA__22235__A2 _22229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23012_ _22985_/X _16945_/Y _22997_/X _23011_/X VGND VGND VPWR VPWR _23013_/A sky130_fd_sc_hd__a211o_4
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20224_ _20644_/A _20224_/B VGND VGND VPWR VPWR _20224_/X sky130_fd_sc_hd__or2_4
XFILLER_85_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17111__B2 _17105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21994__A1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21994__B2 _21992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20155_ _20135_/Y _20136_/Y _11560_/X _20154_/X VGND VGND VPWR VPWR _20155_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15122__B1 _15120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23539__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13095__B _23986_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20086_ _20086_/A VGND VGND VPWR VPWR _20089_/A sky130_fd_sc_hd__inv_2
XFILLER_112_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21746__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23914_ _23692_/CLK _23914_/D VGND VGND VPWR VPWR _23914_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17414__A2 _17340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24369__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_HCLK_A clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23845_ _23845_/CLK _23845_/D VGND VGND VPWR VPWR _14487_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_25_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_50_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11790_ _11821_/A _11790_/B VGND VGND VPWR VPWR _11790_/X sky130_fd_sc_hd__or2_4
X_23776_ _23840_/CLK _23776_/D VGND VGND VPWR VPWR _23776_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14000__A _14000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20988_ _19769_/Y _20851_/X _19770_/X _20675_/X VGND VGND VPWR VPWR _20988_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22171__B2 _22169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22727_ _22727_/A VGND VGND VPWR VPWR _22750_/A sky130_fd_sc_hd__inv_2
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20182__B1 _19313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20721__A2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13460_ _11980_/A _13460_/B VGND VGND VPWR VPWR _13460_/X sky130_fd_sc_hd__and2_4
X_22658_ _22451_/X _22657_/X _14695_/B _22654_/X VGND VGND VPWR VPWR _23108_/D sky130_fd_sc_hd__o22a_4
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14654__B _14654_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12411_ _12398_/A _12409_/X _12411_/C VGND VGND VPWR VPWR _12411_/X sky130_fd_sc_hd__and3_4
X_21609_ _21602_/A VGND VGND VPWR VPWR _21609_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13391_ _11666_/X _13391_/B _13391_/C VGND VGND VPWR VPWR _13425_/B sky130_fd_sc_hd__or3_4
XANTENNA__22474__A2 _22472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22589_ _22420_/X _22586_/X _13165_/B _22583_/X VGND VGND VPWR VPWR _23153_/D sky130_fd_sc_hd__o22a_4
XFILLER_51_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12455__A _12852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15130_ _12252_/A _15128_/X _15129_/X VGND VGND VPWR VPWR _15130_/X sky130_fd_sc_hd__and3_4
XFILLER_16_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12342_ _13726_/A VGND VGND VPWR VPWR _12791_/A sky130_fd_sc_hd__buf_2
X_24328_ _24305_/CLK _19064_/X HRESETn VGND VGND VPWR VPWR _24328_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21682__B1 _23679_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15061_ _14068_/A _23743_/Q VGND VGND VPWR VPWR _15062_/C sky130_fd_sc_hd__or2_4
XANTENNA__15766__A _12795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12273_ _12233_/X VGND VGND VPWR VPWR _12710_/A sky130_fd_sc_hd__buf_2
X_24259_ _24321_/CLK _24259_/D HRESETn VGND VGND VPWR VPWR _24259_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18142__A _18142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14670__A _14071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14012_ _12568_/A _23754_/Q VGND VGND VPWR VPWR _14013_/C sky130_fd_sc_hd__or2_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18820_ _18842_/A VGND VGND VPWR VPWR _18835_/A sky130_fd_sc_hd__buf_2
XANTENNA__13286__A _15689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18850__A1 _17171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12190__A _13056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18751_ _18751_/A _18751_/B _18751_/C VGND VGND VPWR VPWR _18752_/A sky130_fd_sc_hd__and3_4
X_15963_ _16095_/A _15963_/B _15962_/X VGND VGND VPWR VPWR _15963_/X sky130_fd_sc_hd__or3_4
Xclkbuf_7_107_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR _23986_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16597__A _11675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17702_ _16973_/A VGND VGND VPWR VPWR _18459_/A sky130_fd_sc_hd__buf_2
X_14914_ _12250_/A _14914_/B _14914_/C VGND VGND VPWR VPWR _14914_/X sky130_fd_sc_hd__and3_4
XFILLER_49_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15894_ _13551_/X _15838_/B VGND VGND VPWR VPWR _15894_/X sky130_fd_sc_hd__or2_4
X_18682_ _24112_/Q _18681_/X _18610_/X VGND VGND VPWR VPWR _18682_/X sky130_fd_sc_hd__o21a_4
XFILLER_64_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17633_ _17077_/A _17633_/B VGND VGND VPWR VPWR _17633_/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13733__B _13630_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14845_ _14845_/A _14773_/B VGND VGND VPWR VPWR _14846_/C sky130_fd_sc_hd__or2_4
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15006__A _15006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14776_ _13959_/A _14776_/B VGND VGND VPWR VPWR _14778_/B sky130_fd_sc_hd__or2_4
X_17564_ _16235_/X _17564_/B VGND VGND VPWR VPWR _17564_/X sky130_fd_sc_hd__or2_4
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11988_ _16143_/A _11986_/X _11988_/C VGND VGND VPWR VPWR _11989_/C sky130_fd_sc_hd__and3_4
X_19303_ _19302_/X VGND VGND VPWR VPWR _19303_/X sky130_fd_sc_hd__buf_2
XFILLER_17_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13727_ _13735_/A _13727_/B VGND VGND VPWR VPWR _13730_/B sky130_fd_sc_hd__or2_4
X_16515_ _16444_/Y _16514_/X VGND VGND VPWR VPWR _16515_/X sky130_fd_sc_hd__and2_4
XFILLER_1_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17495_ _17495_/A VGND VGND VPWR VPWR _18332_/A sky130_fd_sc_hd__inv_2
XANTENNA__14845__A _14845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18317__A _18204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19234_ _24285_/Q _19234_/B VGND VGND VPWR VPWR _19236_/A sky130_fd_sc_hd__and2_4
X_13658_ _15442_/A _13658_/B _13658_/C VGND VGND VPWR VPWR _13658_/X sky130_fd_sc_hd__or3_4
X_16446_ _11715_/A _16381_/B VGND VGND VPWR VPWR _16447_/C sky130_fd_sc_hd__or2_4
XFILLER_13_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12609_ _12964_/A _12596_/X _12609_/C VGND VGND VPWR VPWR _12609_/X sky130_fd_sc_hd__or3_4
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16377_ _16302_/X _16377_/B VGND VGND VPWR VPWR _16377_/X sky130_fd_sc_hd__or2_4
X_19165_ _19165_/A VGND VGND VPWR VPWR _19165_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13589_ _13579_/X VGND VGND VPWR VPWR _13590_/B sky130_fd_sc_hd__inv_2
XANTENNA__12365__A _15484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20476__A1 _20468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15328_ _15333_/A _15263_/B VGND VGND VPWR VPWR _15329_/C sky130_fd_sc_hd__or2_4
X_18116_ _17910_/X _17982_/Y _17921_/X _17934_/Y VGND VGND VPWR VPWR _18116_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19096_ _19087_/X _19095_/X _19087_/X _19092_/A VGND VGND VPWR VPWR _19096_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15676__A _12742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15259_ _14315_/A _15259_/B VGND VGND VPWR VPWR _15259_/X sky130_fd_sc_hd__or2_4
X_18047_ _18047_/A _18046_/X VGND VGND VPWR VPWR _18047_/X sky130_fd_sc_hd__or2_4
XANTENNA__22217__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19618__B1 HRDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21425__B1 _23823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15395__B _15458_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13196__A _15706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21976__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19998_ _19994_/X _17661_/A _19976_/X _19997_/X VGND VGND VPWR VPWR _19999_/A sky130_fd_sc_hd__o22a_4
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18949_ _18923_/Y _18924_/Y _11532_/X VGND VGND VPWR VPWR _18949_/X sky130_fd_sc_hd__o21a_4
XFILLER_86_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21728__B2 _21723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21960_ _21852_/X _21959_/X _14683_/B _21956_/X VGND VGND VPWR VPWR _23524_/D sky130_fd_sc_hd__o22a_4
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16300__A _11851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20911_ _20616_/X _20899_/X _20757_/X _20910_/Y VGND VGND VPWR VPWR _20911_/X sky130_fd_sc_hd__a211o_4
XFILLER_94_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21891_ _21884_/A VGND VGND VPWR VPWR _21891_/X sky130_fd_sc_hd__buf_2
X_23630_ _23342_/CLK _23630_/D VGND VGND VPWR VPWR _15700_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20842_ _20223_/A VGND VGND VPWR VPWR _20842_/X sky130_fd_sc_hd__buf_2
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23561_ _23561_/CLK _23561_/D VGND VGND VPWR VPWR _23561_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20773_ _20773_/A VGND VGND VPWR VPWR _20773_/Y sky130_fd_sc_hd__inv_2
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14755__A _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21900__B2 _21898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22512_ _22460_/X _22507_/X _14905_/B _22476_/A VGND VGND VPWR VPWR _22512_/X sky130_fd_sc_hd__o22a_4
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23492_ _23433_/CLK _23492_/D VGND VGND VPWR VPWR _14646_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22443_ _22442_/X _22440_/X _13696_/B _22435_/X VGND VGND VPWR VPWR _22443_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12275__A _12238_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24122__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18124__A3 _18120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21588__A _21595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21664__B1 _15838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22374_ _22134_/X _22368_/X _14511_/B _22372_/X VGND VGND VPWR VPWR _22374_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17332__A1 _14988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24113_ _24199_/CLK _24113_/D HRESETn VGND VGND VPWR VPWR _16964_/A sky130_fd_sc_hd__dfrtp_4
X_21325_ _21256_/X _21319_/X _23887_/Q _21323_/X VGND VGND VPWR VPWR _21325_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14490__A _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23361__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24044_ _24044_/CLK _21040_/X VGND VGND VPWR VPWR _15490_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19085__A1 _18965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21256_ _21256_/A VGND VGND VPWR VPWR _21256_/X sky130_fd_sc_hd__buf_2
XFILLER_89_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20207_ _20206_/X VGND VGND VPWR VPWR _20421_/A sky130_fd_sc_hd__buf_2
XFILLER_89_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11619__A _11618_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18832__A1 _12430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21187_ _21180_/A VGND VGND VPWR VPWR _21187_/X sky130_fd_sc_hd__buf_2
X_20138_ IRQ[15] VGND VGND VPWR VPWR _20138_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22212__A _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13834__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12960_ _12596_/A _12958_/X _12960_/C VGND VGND VPWR VPWR _12964_/B sky130_fd_sc_hd__and3_4
X_20069_ _20069_/A VGND VGND VPWR VPWR _20069_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16210__A _16194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21195__A2 _21190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11911_ _11911_/A VGND VGND VPWR VPWR _11912_/A sky130_fd_sc_hd__buf_2
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12891_ _12891_/A _12887_/X _12890_/X VGND VGND VPWR VPWR _12892_/B sky130_fd_sc_hd__or3_4
XFILLER_98_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14630_ _11929_/A _14626_/X _14630_/C VGND VGND VPWR VPWR _14630_/X sky130_fd_sc_hd__or3_4
X_11842_ _11842_/A VGND VGND VPWR VPWR _11842_/X sky130_fd_sc_hd__buf_2
X_23828_ _23315_/CLK _23828_/D VGND VGND VPWR VPWR _23828_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19371__A2_N _17953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22144__B2 _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14561_ _13770_/A _14553_/X _14561_/C VGND VGND VPWR VPWR _14561_/X sky130_fd_sc_hd__and3_4
X_11773_ _11729_/X VGND VGND VPWR VPWR _11773_/X sky130_fd_sc_hd__buf_2
X_23759_ _24047_/CLK _23759_/D VGND VGND VPWR VPWR _13435_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14665__A _14679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22695__A2 _22693_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18137__A _18137_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13512_ _12591_/X VGND VGND VPWR VPWR _13558_/A sky130_fd_sc_hd__buf_2
X_16300_ _11851_/X _16299_/X VGND VGND VPWR VPWR _16300_/X sky130_fd_sc_hd__and2_4
X_17280_ _17902_/B VGND VGND VPWR VPWR _17280_/Y sky130_fd_sc_hd__inv_2
X_14492_ _11842_/A _11618_/A _14461_/X _11596_/A _14491_/X VGND VGND VPWR VPWR _14492_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22882__A _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16231_ _16231_/A _16231_/B _16231_/C VGND VGND VPWR VPWR _16232_/C sky130_fd_sc_hd__or3_4
X_13443_ _13437_/X _13530_/B VGND VGND VPWR VPWR _13443_/X sky130_fd_sc_hd__or2_4
XFILLER_55_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15582__B1 _11596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19848__B1 _19592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12185__A _12184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16162_ _13388_/A VGND VGND VPWR VPWR _16162_/X sky130_fd_sc_hd__buf_2
XFILLER_70_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13374_ _13357_/X _13372_/X _13374_/C VGND VGND VPWR VPWR _13381_/B sky130_fd_sc_hd__and3_4
XANTENNA__17695__B _17375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15113_ _11710_/A _23615_/Q VGND VGND VPWR VPWR _15113_/X sky130_fd_sc_hd__or2_4
X_12325_ _12740_/A _12323_/X _12325_/C VGND VGND VPWR VPWR _12325_/X sky130_fd_sc_hd__and3_4
XANTENNA__15496__A _13735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16093_ _16097_/A _23735_/Q VGND VGND VPWR VPWR _16094_/C sky130_fd_sc_hd__or2_4
XANTENNA__12913__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15044_ _13951_/A _23839_/Q VGND VGND VPWR VPWR _15045_/C sky130_fd_sc_hd__or2_4
X_19921_ _19916_/X _24144_/Q _19917_/X _20939_/B VGND VGND VPWR VPWR _24144_/D sky130_fd_sc_hd__o22a_4
X_12256_ _13678_/A VGND VGND VPWR VPWR _12257_/A sky130_fd_sc_hd__buf_2
XFILLER_68_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21958__B2 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19852_ _19730_/A _19846_/B _19621_/A _19846_/B VGND VGND VPWR VPWR _19852_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18823__A1 _12184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12187_ _12186_/X VGND VGND VPWR VPWR _12187_/X sky130_fd_sc_hd__buf_2
XFILLER_110_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18803_ _18789_/A VGND VGND VPWR VPWR _18803_/X sky130_fd_sc_hd__buf_2
X_19783_ _19419_/X _19782_/X _16652_/A _19678_/X VGND VGND VPWR VPWR _19783_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19324__A2_N _18168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16995_ _16969_/A VGND VGND VPWR VPWR _16998_/A sky130_fd_sc_hd__buf_2
XFILLER_84_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22122__A _20747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18734_ _18713_/A _18733_/X VGND VGND VPWR VPWR _18734_/Y sky130_fd_sc_hd__nor2_4
XFILLER_95_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15946_ _15976_/A _15944_/X _15946_/C VGND VGND VPWR VPWR _15946_/X sky130_fd_sc_hd__and3_4
XFILLER_7_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16120__A _16147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21186__A2 _21183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24352__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18665_ _18607_/X _18610_/X _18607_/X _18610_/X VGND VGND VPWR VPWR _18665_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18051__A2 _18020_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15877_ _15884_/A _15815_/B VGND VGND VPWR VPWR _15877_/X sky130_fd_sc_hd__or2_4
XFILLER_64_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20933__A2 _20924_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22776__B _17032_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17616_ _17609_/Y _17615_/X _17323_/X VGND VGND VPWR VPWR _17616_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19339__A2_N _18455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19431__A _19433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14828_ _13690_/A _14826_/X _14828_/C VGND VGND VPWR VPWR _14828_/X sky130_fd_sc_hd__and3_4
X_18596_ _18557_/A VGND VGND VPWR VPWR _22913_/B sky130_fd_sc_hd__inv_2
XFILLER_91_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22135__B2 _22132_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23234__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17547_ _16376_/X _17549_/B VGND VGND VPWR VPWR _17547_/X sky130_fd_sc_hd__or2_4
X_14759_ _12883_/A _14759_/B VGND VGND VPWR VPWR _14760_/C sky130_fd_sc_hd__or2_4
XANTENNA__14575__A _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17478_ _16640_/X _17364_/X _17365_/X VGND VGND VPWR VPWR _17479_/B sky130_fd_sc_hd__o21a_4
X_19217_ _19217_/A _19217_/B VGND VGND VPWR VPWR _19218_/B sky130_fd_sc_hd__and2_4
X_16429_ _16087_/X _16427_/X _16428_/X VGND VGND VPWR VPWR _16433_/B sky130_fd_sc_hd__and3_4
XANTENNA__12095__A _12068_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22438__A2 _22428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16790__A _11782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19148_ _24314_/Q _19134_/X _19147_/Y VGND VGND VPWR VPWR _19148_/X sky130_fd_sc_hd__o21a_4
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21201__A _21180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13919__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19079_ _19079_/A VGND VGND VPWR VPWR _19079_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21110_ _21110_/A VGND VGND VPWR VPWR _21110_/Y sky130_fd_sc_hd__inv_2
X_22090_ _22088_/X _22089_/X _15969_/B _22084_/X VGND VGND VPWR VPWR _22090_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16014__B _23352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21041_ _21027_/A VGND VGND VPWR VPWR _21041_/X sky130_fd_sc_hd__buf_2
XFILLER_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22610__A2 _22607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15853__B _15792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14300__A1 _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13654__A _13654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22992_ _22998_/A _22992_/B VGND VGND VPWR VPWR _22994_/B sky130_fd_sc_hd__or2_4
XANTENNA__22967__A _22967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22374__B2 _22372_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21943_ _21823_/X _21938_/X _23536_/Q _21942_/X VGND VGND VPWR VPWR _23536_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_7_0_HCLK_A clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21874_ _21791_/X _21873_/X _23581_/Q _21870_/X VGND VGND VPWR VPWR _23581_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22126__B2 _22120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23485_/CLK _23613_/D VGND VGND VPWR VPWR _23613_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _20578_/A VGND VGND VPWR VPWR _20825_/X sky130_fd_sc_hd__buf_2
XFILLER_93_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22677__A2 _22672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14485__A _15404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19542__A2 _19877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23544_ _23539_/CLK _21932_/X VGND VGND VPWR VPWR _23544_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20756_ _20802_/A _20755_/X VGND VGND VPWR VPWR _20756_/X sky130_fd_sc_hd__or2_4
XFILLER_93_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11621__B _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23475_ _23699_/CLK _22039_/X VGND VGND VPWR VPWR _12980_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22429__A2 _22428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20687_ _20494_/X _20685_/X _24332_/Q _20686_/X VGND VGND VPWR VPWR _20687_/X sky130_fd_sc_hd__o22a_4
XFILLER_7_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22426_ _22425_/X _22416_/X _13427_/B _22423_/X VGND VGND VPWR VPWR _23247_/D sky130_fd_sc_hd__o22a_4
XFILLER_6_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21101__A2 _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22207__A _22207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14932__B _14868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13829__A _13645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21111__A _21583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22357_ _22105_/X _22354_/X _13149_/B _22351_/X VGND VGND VPWR VPWR _23281_/D sky130_fd_sc_hd__o22a_4
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12733__A _12713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12110_ _11971_/A _23869_/Q VGND VGND VPWR VPWR _12110_/X sky130_fd_sc_hd__or2_4
X_21308_ _21227_/X _21305_/X _23899_/Q _21302_/X VGND VGND VPWR VPWR _23899_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13090_ _13065_/A VGND VGND VPWR VPWR _13115_/A sky130_fd_sc_hd__buf_2
X_22288_ _22127_/X _22286_/X _13702_/B _22283_/X VGND VGND VPWR VPWR _22288_/X sky130_fd_sc_hd__o22a_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12041_ _11903_/A VGND VGND VPWR VPWR _16714_/A sky130_fd_sc_hd__buf_2
X_24027_ _23515_/CLK _24027_/D VGND VGND VPWR VPWR _24027_/Q sky130_fd_sc_hd__dfxtp_4
X_21239_ _20464_/A VGND VGND VPWR VPWR _21239_/X sky130_fd_sc_hd__buf_2
XANTENNA__23107__CLK _23107_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18805__A1 _17297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22601__A2 _22600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20612__A1 _20511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23038__A _18000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20612__B2 _20592_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15800_ _15823_/A _15798_/X _15799_/X VGND VGND VPWR VPWR _15800_/X sky130_fd_sc_hd__and3_4
XFILLER_24_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13564__A _12753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13992_ _13992_/A VGND VGND VPWR VPWR _14037_/A sky130_fd_sc_hd__buf_2
X_16780_ _16045_/A _16762_/X _16780_/C VGND VGND VPWR VPWR _16780_/X sky130_fd_sc_hd__or3_4
XANTENNA__14379__B _14379_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12943_ _12974_/A _12943_/B VGND VGND VPWR VPWR _12943_/X sky130_fd_sc_hd__or2_4
X_15731_ _12765_/X _15729_/X _15730_/X VGND VGND VPWR VPWR _15735_/B sky130_fd_sc_hd__and3_4
XFILLER_59_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18450_ _18216_/X _17349_/A _18448_/X _18398_/X _18449_/Y VGND VGND VPWR VPWR _18450_/X
+ sky130_fd_sc_hd__a32o_4
X_12874_ _12874_/A _12953_/B VGND VGND VPWR VPWR _12875_/C sky130_fd_sc_hd__or2_4
X_15662_ _12725_/A _15724_/B VGND VGND VPWR VPWR _15662_/X sky130_fd_sc_hd__or2_4
XANTENNA__16595__A2 _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17401_ _22017_/B VGND VGND VPWR VPWR _20197_/B sky130_fd_sc_hd__inv_2
XFILLER_27_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11825_ _11746_/X VGND VGND VPWR VPWR _11834_/A sky130_fd_sc_hd__buf_2
X_14613_ _14146_/X _14613_/B _14612_/X VGND VGND VPWR VPWR _14613_/X sky130_fd_sc_hd__or3_4
XFILLER_2_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15593_ _15617_/A _24011_/Q VGND VGND VPWR VPWR _15595_/B sky130_fd_sc_hd__or2_4
X_18381_ _18381_/A VGND VGND VPWR VPWR _18381_/X sky130_fd_sc_hd__buf_2
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12908__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11812__A _11692_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _13711_/X _14544_/B _14543_/X VGND VGND VPWR VPWR _14544_/X sky130_fd_sc_hd__and3_4
X_17332_ _14988_/X _17220_/A _17330_/X _17331_/X VGND VGND VPWR VPWR _17332_/X sky130_fd_sc_hd__o22a_4
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11818_/A _24030_/Q VGND VGND VPWR VPWR _11761_/B sky130_fd_sc_hd__or2_4
XFILLER_72_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18741__B1 _18864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _12533_/A _14471_/X _14475_/C VGND VGND VPWR VPWR _14475_/X sky130_fd_sc_hd__or3_4
X_17263_ _17039_/X _17262_/X _17043_/X VGND VGND VPWR VPWR _17263_/Y sky130_fd_sc_hd__o21ai_4
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _13231_/A VGND VGND VPWR VPWR _15774_/A sky130_fd_sc_hd__buf_2
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19002_ _19002_/A VGND VGND VPWR VPWR _19002_/X sky130_fd_sc_hd__buf_2
XANTENNA__20844__B _20844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13426_ _13350_/Y _13425_/X VGND VGND VPWR VPWR _13426_/X sky130_fd_sc_hd__and2_4
X_16214_ _16198_/A _16210_/X _16213_/X VGND VGND VPWR VPWR _16215_/C sky130_fd_sc_hd__or3_4
X_17194_ _13425_/X VGND VGND VPWR VPWR _17194_/X sky130_fd_sc_hd__buf_2
XANTENNA__22117__A _20696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16145_ _16145_/A _23095_/Q VGND VGND VPWR VPWR _16147_/B sky130_fd_sc_hd__or2_4
X_13357_ _12769_/A VGND VGND VPWR VPWR _13357_/X sky130_fd_sc_hd__buf_2
XANTENNA__13739__A _12612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12308_ _12747_/A VGND VGND VPWR VPWR _12705_/A sky130_fd_sc_hd__buf_2
X_16076_ _16231_/A _16076_/B _16075_/X VGND VGND VPWR VPWR _16077_/C sky130_fd_sc_hd__or3_4
XFILLER_115_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21956__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13288_ _13283_/X _23728_/Q VGND VGND VPWR VPWR _13289_/C sky130_fd_sc_hd__or2_4
XFILLER_29_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15027_ _14151_/A _23807_/Q VGND VGND VPWR VPWR _15028_/C sky130_fd_sc_hd__or2_4
X_19904_ _24157_/Q _19899_/X _20224_/B _19903_/X VGND VGND VPWR VPWR _24157_/D sky130_fd_sc_hd__o22a_4
X_12239_ _12238_/X VGND VGND VPWR VPWR _12240_/A sky130_fd_sc_hd__buf_2
XANTENNA__15954__A _15980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24032__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16769__B _16708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19835_ _19877_/A _19867_/B VGND VGND VPWR VPWR _19835_/X sky130_fd_sc_hd__or2_4
XFILLER_25_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13474__A _11913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19766_ _19766_/A _19766_/B VGND VGND VPWR VPWR _19766_/X sky130_fd_sc_hd__and2_4
X_16978_ _17681_/A _16978_/B VGND VGND VPWR VPWR _16979_/B sky130_fd_sc_hd__or2_4
XFILLER_96_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22787__A _14786_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22356__A1 _22103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21159__A2 _21154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22356__B2 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18717_ _17101_/X _17258_/Y _18249_/A _18716_/X VGND VGND VPWR VPWR _18718_/A sky130_fd_sc_hd__a211o_4
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21691__A _21705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15929_ _12503_/A VGND VGND VPWR VPWR _15929_/X sky130_fd_sc_hd__buf_2
X_19697_ _19419_/A VGND VGND VPWR VPWR _19697_/X sky130_fd_sc_hd__buf_2
XFILLER_80_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17232__B1 _14723_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19772__A2 _19592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18648_ _17743_/A _18647_/X _17743_/A _18647_/X VGND VGND VPWR VPWR _18648_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18579_ _18621_/B _18578_/X VGND VGND VPWR VPWR _18579_/X sky130_fd_sc_hd__or2_4
XANTENNA__22659__A2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12818__A _12802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20610_ _20610_/A VGND VGND VPWR VPWR _21256_/A sky130_fd_sc_hd__buf_2
XFILLER_33_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11722__A _13998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21590_ _21590_/A VGND VGND VPWR VPWR _21605_/A sky130_fd_sc_hd__buf_2
XANTENNA__21331__A2 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16009__B _23256_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20541_ _24402_/Q _20405_/X _24434_/Q _20449_/X VGND VGND VPWR VPWR _20541_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23260_ _23260_/CLK _22395_/X VGND VGND VPWR VPWR _16602_/B sky130_fd_sc_hd__dfxtp_4
X_20472_ _20470_/Y _20521_/B VGND VGND VPWR VPWR _20472_/X sky130_fd_sc_hd__or2_4
XFILLER_105_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22211_ _22081_/X _22208_/X _16791_/B _22205_/X VGND VGND VPWR VPWR _23387_/D sky130_fd_sc_hd__o22a_4
XFILLER_69_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_15_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR _23433_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21095__B2 _21093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23191_ _23313_/CLK _22531_/X VGND VGND VPWR VPWR _16096_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12553__A _12553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_78_0_HCLK clkbuf_7_78_0_HCLK/A VGND VGND VPWR VPWR _23931_/CLK sky130_fd_sc_hd__clkbuf_1
X_22142_ _22141_/X _22137_/X _15277_/B _22132_/X VGND VGND VPWR VPWR _23426_/D sky130_fd_sc_hd__o22a_4
XFILLER_69_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15864__A _13554_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22073_ _20276_/A VGND VGND VPWR VPWR _22073_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19336__A _19336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21024_ _20419_/X _21023_/X _24056_/Q _21020_/X VGND VGND VPWR VPWR _21024_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22595__B2 _22590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15583__B _15522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22697__A _22683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22975_ _22982_/A _22975_/B _22974_/X VGND VGND VPWR VPWR _22975_/X sky130_fd_sc_hd__and3_4
XFILLER_112_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21926_ _21795_/X _21924_/X _23548_/Q _21921_/X VGND VGND VPWR VPWR _21926_/X sky130_fd_sc_hd__o22a_4
XFILLER_76_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21857_ _21287_/A VGND VGND VPWR VPWR _21857_/X sky130_fd_sc_hd__buf_2
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__A _12728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11610_/A VGND VGND VPWR VPWR _11611_/A sky130_fd_sc_hd__buf_2
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _20704_/X _20807_/Y _19212_/A _20325_/X VGND VGND VPWR VPWR _20808_/X sky130_fd_sc_hd__o22a_4
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12590_ _13731_/A VGND VGND VPWR VPWR _12964_/A sky130_fd_sc_hd__buf_2
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21788_ _21787_/X VGND VGND VPWR VPWR _21788_/X sky130_fd_sc_hd__buf_2
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21322__A2 _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _11541_/A IRQ[2] VGND VGND VPWR VPWR _11541_/Y sky130_fd_sc_hd__nand2_4
X_23527_ _23591_/CLK _21955_/X VGND VGND VPWR VPWR _23527_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20739_ _20305_/X VGND VGND VPWR VPWR _20739_/X sky130_fd_sc_hd__buf_2
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _11798_/A _14243_/X _14260_/C VGND VGND VPWR VPWR _14260_/X sky130_fd_sc_hd__or3_4
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23458_ _23907_/CLK _23458_/D VGND VGND VPWR VPWR _15296_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14662__B _14662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13211_ _13211_/A _13211_/B _13210_/X VGND VGND VPWR VPWR _13219_/B sky130_fd_sc_hd__or3_4
X_22409_ _22408_/X _22404_/X _12206_/B _22399_/X VGND VGND VPWR VPWR _23254_/D sky130_fd_sc_hd__o22a_4
X_14191_ _11738_/A VGND VGND VPWR VPWR _14201_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17829__A2 _17827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23389_ _23100_/CLK _22209_/X VGND VGND VPWR VPWR _12162_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12463__A _12865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13142_ _12720_/A _13140_/X _13141_/X VGND VGND VPWR VPWR _13142_/X sky130_fd_sc_hd__and3_4
XFILLER_100_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21776__A _21740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20680__A _20447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15774__A _15774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13073_ _12613_/A VGND VGND VPWR VPWR _13082_/A sky130_fd_sc_hd__buf_2
X_17950_ _18171_/A VGND VGND VPWR VPWR _17950_/X sky130_fd_sc_hd__buf_2
XFILLER_65_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21389__A2 _21383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12024_ _12024_/A _23870_/Q VGND VGND VPWR VPWR _12025_/C sky130_fd_sc_hd__or2_4
X_16901_ _16524_/Y _16900_/X _16817_/X _16897_/X VGND VGND VPWR VPWR _16902_/A sky130_fd_sc_hd__a211o_4
X_17881_ _16935_/X _17775_/X _17006_/X _17880_/X VGND VGND VPWR VPWR _17881_/X sky130_fd_sc_hd__o22a_4
XFILLER_61_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19620_ _19645_/A VGND VGND VPWR VPWR _19808_/A sky130_fd_sc_hd__inv_2
X_16832_ _16824_/D _13593_/X _13580_/Y VGND VGND VPWR VPWR _16832_/X sky130_fd_sc_hd__o21a_4
XFILLER_117_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22338__B2 _22337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19551_ _19551_/A VGND VGND VPWR VPWR _19551_/X sky130_fd_sc_hd__buf_2
XANTENNA__19203__A1 _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16763_ _16772_/A _23931_/Q VGND VGND VPWR VPWR _16763_/X sky130_fd_sc_hd__or2_4
X_13975_ _12217_/A _13975_/B _13974_/X VGND VGND VPWR VPWR _13979_/B sky130_fd_sc_hd__and3_4
XFILLER_81_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18502_ _18443_/A VGND VGND VPWR VPWR _18697_/A sky130_fd_sc_hd__buf_2
XFILLER_111_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15714_ _13129_/A _15652_/B VGND VGND VPWR VPWR _15714_/X sky130_fd_sc_hd__or2_4
X_12926_ _12926_/A _23507_/Q VGND VGND VPWR VPWR _12926_/X sky130_fd_sc_hd__or2_4
X_19482_ _19598_/A _19561_/A VGND VGND VPWR VPWR _19538_/A sky130_fd_sc_hd__or2_4
X_16694_ _16714_/A _16759_/B VGND VGND VPWR VPWR _16695_/C sky130_fd_sc_hd__or2_4
XFILLER_59_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21561__A2 _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14837__B _14779_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18433_ _18340_/X _18431_/X _18377_/X _18432_/X VGND VGND VPWR VPWR _18433_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21016__A _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15645_ _13918_/A _15645_/B _15645_/C VGND VGND VPWR VPWR _15645_/X sky130_fd_sc_hd__and3_4
X_12857_ _12851_/A _12857_/B VGND VGND VPWR VPWR _12857_/X sky130_fd_sc_hd__or2_4
XFILLER_76_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12638__A _12638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18309__A3 _18305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21849__B1 _14304_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11808_ _11820_/A _11808_/B _11808_/C VGND VGND VPWR VPWR _11809_/C sky130_fd_sc_hd__and3_4
X_18364_ _17837_/X _18109_/X _17846_/X _18112_/X VGND VGND VPWR VPWR _18364_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12788_ _12799_/A _23924_/Q VGND VGND VPWR VPWR _12788_/X sky130_fd_sc_hd__or2_4
X_15576_ _15576_/A _23691_/Q VGND VGND VPWR VPWR _15576_/X sky130_fd_sc_hd__or2_4
XANTENNA__21313__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22510__B2 _22504_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17315_/A VGND VGND VPWR VPWR _17618_/C sky130_fd_sc_hd__buf_2
X_11739_ _13706_/A VGND VGND VPWR VPWR _11740_/A sky130_fd_sc_hd__buf_2
X_14527_ _14519_/X _14450_/B VGND VGND VPWR VPWR _14527_/X sky130_fd_sc_hd__or2_4
XANTENNA__15949__A _13437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18295_ _18295_/A _17510_/B VGND VGND VPWR VPWR _18298_/B sky130_fd_sc_hd__nor2_4
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17246_ _17222_/X _17815_/A _17826_/A _17218_/X VGND VGND VPWR VPWR _17246_/X sky130_fd_sc_hd__o22a_4
X_14458_ _15404_/A _14458_/B _14458_/C VGND VGND VPWR VPWR _14459_/C sky130_fd_sc_hd__and3_4
X_13409_ _13358_/X _13340_/B VGND VGND VPWR VPWR _13411_/B sky130_fd_sc_hd__or2_4
XANTENNA__13469__A _13437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21077__B2 _21072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14389_ _13886_/A _14365_/X _14389_/C VGND VGND VPWR VPWR _14423_/B sky130_fd_sc_hd__or3_4
X_17177_ _17141_/X _17174_/X _17163_/A _17176_/X VGND VGND VPWR VPWR _17177_/X sky130_fd_sc_hd__o22a_4
X_16128_ _16108_/A _24055_/Q VGND VGND VPWR VPWR _16129_/C sky130_fd_sc_hd__or2_4
XANTENNA__21686__A _21690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20590__A _20590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22026__B1 _23484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15684__A _12720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16059_ _11684_/X _16055_/X _16058_/X VGND VGND VPWR VPWR _16060_/C sky130_fd_sc_hd__or3_4
XFILLER_88_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19818_ _19818_/A VGND VGND VPWR VPWR _19846_/B sky130_fd_sc_hd__buf_2
XANTENNA__11717__A _16072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23572__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19749_ _19554_/X _19740_/X _19746_/Y _19581_/X _19748_/Y VGND VGND VPWR VPWR _19749_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_84_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17205__B1 _15909_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13932__A _13611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22760_ _22730_/Y _22758_/B VGND VGND VPWR VPWR _22763_/B sky130_fd_sc_hd__or2_4
XFILLER_25_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21552__A2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21711_ _21541_/X _21705_/X _13530_/B _21709_/X VGND VGND VPWR VPWR _23663_/D sky130_fd_sc_hd__o22a_4
X_22691_ _20591_/A _22686_/X _13340_/B _22690_/X VGND VGND VPWR VPWR _23088_/D sky130_fd_sc_hd__o22a_4
XFILLER_94_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12548__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24430_ _24334_/CLK _18791_/X HRESETn VGND VGND VPWR VPWR _24430_/Q sky130_fd_sc_hd__dfrtp_4
X_21642_ _21506_/X _21641_/X _23709_/Q _21638_/X VGND VGND VPWR VPWR _23709_/D sky130_fd_sc_hd__o22a_4
XFILLER_40_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22501__B2 _22497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24361_ _24330_/CLK _18908_/X HRESETn VGND VGND VPWR VPWR _24361_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__15859__A _13572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21573_ _21572_/X _21568_/X _15260_/B _21563_/X VGND VGND VPWR VPWR _23746_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23312_ _23699_/CLK _22314_/X VGND VGND VPWR VPWR _13304_/B sky130_fd_sc_hd__dfxtp_4
X_20524_ _20468_/X _20523_/Y _24275_/Q _20301_/X VGND VGND VPWR VPWR _20524_/X sky130_fd_sc_hd__o22a_4
X_24292_ _24293_/CLK _24292_/D HRESETn VGND VGND VPWR VPWR _19113_/A sky130_fd_sc_hd__dfrtp_4
X_23243_ _24011_/CLK _23243_/D VGND VGND VPWR VPWR _15522_/B sky130_fd_sc_hd__dfxtp_4
X_20455_ _20321_/X _20454_/X _24310_/Q _20330_/X VGND VGND VPWR VPWR _20455_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12283__A _13025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20815__A1 _24231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23174_ _23494_/CLK _22555_/X VGND VGND VPWR VPWR _14275_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20386_ _20291_/X _20386_/B VGND VGND VPWR VPWR _20386_/Y sky130_fd_sc_hd__nor2_4
XFILLER_88_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22125_ _22125_/A VGND VGND VPWR VPWR _22125_/X sky130_fd_sc_hd__buf_2
XFILLER_106_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22056_ _22035_/A VGND VGND VPWR VPWR _22056_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_8_0_HCLK clkbuf_6_4_0_HCLK/X VGND VGND VPWR VPWR _24066_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_88_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20579__B1 _24432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21007_ _21007_/A _20197_/B _21212_/B VGND VGND VPWR VPWR _21008_/A sky130_fd_sc_hd__or3_4
XFILLER_88_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21240__B2 _21230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17995__A1 _17989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14938__A _13998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13760_ _12652_/A _13760_/B VGND VGND VPWR VPWR _13760_/X sky130_fd_sc_hd__or2_4
X_22958_ _18453_/X _22950_/X VGND VGND VPWR VPWR _22958_/X sky130_fd_sc_hd__or2_4
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12711_ _12711_/A _12711_/B VGND VGND VPWR VPWR _12711_/X sky130_fd_sc_hd__or2_4
X_21909_ _21852_/X _21908_/X _23556_/Q _21905_/X VGND VGND VPWR VPWR _23556_/D sky130_fd_sc_hd__o22a_4
X_13691_ _13880_/A VGND VGND VPWR VPWR _13699_/A sky130_fd_sc_hd__buf_2
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22889_ _22980_/A VGND VGND VPWR VPWR _22889_/X sky130_fd_sc_hd__buf_2
XANTENNA__12458__A _12458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12642_ _12604_/A _12525_/B VGND VGND VPWR VPWR _12642_/X sky130_fd_sc_hd__or2_4
X_15430_ _15430_/A _23820_/Q VGND VGND VPWR VPWR _15431_/C sky130_fd_sc_hd__or2_4
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15361_ _11638_/A _15361_/B _15360_/X VGND VGND VPWR VPWR _15361_/X sky130_fd_sc_hd__or3_4
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23051__A _23051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12573_ _13708_/A VGND VGND VPWR VPWR _14009_/A sky130_fd_sc_hd__buf_2
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14673__A _14673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18172__A1 _16945_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17100_ _17161_/A VGND VGND VPWR VPWR _17100_/X sky130_fd_sc_hd__buf_2
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11524_ _11524_/A _18996_/A VGND VGND VPWR VPWR _11524_/X sky130_fd_sc_hd__or2_4
X_14312_ _15556_/A _23398_/Q VGND VGND VPWR VPWR _14312_/X sky130_fd_sc_hd__or2_4
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15292_ _14158_/A _15292_/B VGND VGND VPWR VPWR _15292_/X sky130_fd_sc_hd__or2_4
X_18080_ _17794_/X _18075_/Y _18076_/X _18079_/X VGND VGND VPWR VPWR _18080_/X sky130_fd_sc_hd__a211o_4
XFILLER_12_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23445__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22890__A _20196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _14243_/A _14243_/B _14242_/X VGND VGND VPWR VPWR _14243_/X sky130_fd_sc_hd__and3_4
X_17031_ _17033_/A VGND VGND VPWR VPWR _17032_/B sky130_fd_sc_hd__buf_2
XANTENNA__13289__A _12540_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12193__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14174_ _11839_/X _11615_/X _14129_/X _11594_/A _14173_/X VGND VGND VPWR VPWR _14174_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_119_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_61_0_HCLK clkbuf_6_30_0_HCLK/X VGND VGND VPWR VPWR _23889_/CLK sky130_fd_sc_hd__clkbuf_1
X_13125_ _13101_/A _13121_/X _13124_/X VGND VGND VPWR VPWR _13133_/B sky130_fd_sc_hd__or3_4
X_18982_ _18982_/A VGND VGND VPWR VPWR _18982_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12921__A _13041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22559__B2 _22554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13056_ _13056_/A _13055_/X VGND VGND VPWR VPWR _13056_/X sky130_fd_sc_hd__and2_4
X_17933_ _17933_/A VGND VGND VPWR VPWR _17933_/X sky130_fd_sc_hd__buf_2
XFILLER_26_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16238__A1 _16155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12640__B _12640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12007_ _11916_/X VGND VGND VPWR VPWR _12011_/A sky130_fd_sc_hd__buf_2
XFILLER_94_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15009__A _15032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21231__B2 _21230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17864_ _17864_/A VGND VGND VPWR VPWR _17864_/X sky130_fd_sc_hd__buf_2
XFILLER_94_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19603_ _19603_/A _19638_/A VGND VGND VPWR VPWR _19826_/B sky130_fd_sc_hd__or2_4
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21782__A2 _21755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16815_ _16815_/A VGND VGND VPWR VPWR _16815_/Y sky130_fd_sc_hd__inv_2
X_17795_ _17860_/A VGND VGND VPWR VPWR _17962_/A sky130_fd_sc_hd__buf_2
XANTENNA__14848__A _11669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19534_ _19793_/A VGND VGND VPWR VPWR _19534_/X sky130_fd_sc_hd__buf_2
XFILLER_47_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17224__A _17224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13752__A _12937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16746_ _11782_/A _16744_/X _16746_/C VGND VGND VPWR VPWR _16746_/X sky130_fd_sc_hd__and3_4
X_13958_ _14172_/A _13933_/X _13941_/X _13948_/X _13957_/X VGND VGND VPWR VPWR _13958_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_34_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12909_ _12874_/A _12909_/B VGND VGND VPWR VPWR _12910_/C sky130_fd_sc_hd__or2_4
X_19465_ _24153_/Q _19459_/X HRDATA[27] _19460_/X VGND VGND VPWR VPWR _19465_/X sky130_fd_sc_hd__o22a_4
X_16677_ _16677_/A _16661_/X _16676_/X VGND VGND VPWR VPWR _16677_/X sky130_fd_sc_hd__or3_4
XFILLER_62_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13889_ _13911_/A _13887_/X _13888_/X VGND VGND VPWR VPWR _13889_/X sky130_fd_sc_hd__and3_4
XFILLER_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18416_ _18011_/X _18383_/B _18413_/Y _18016_/X _22962_/B VGND VGND VPWR VPWR _18416_/X
+ sky130_fd_sc_hd__a32o_4
X_15628_ _15628_/A _15620_/X _15627_/X VGND VGND VPWR VPWR _15644_/B sky130_fd_sc_hd__and3_4
XFILLER_59_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24220__CLK _24187_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19396_ _19385_/A VGND VGND VPWR VPWR _19396_/X sky130_fd_sc_hd__buf_2
X_18347_ _18533_/A _16999_/C VGND VGND VPWR VPWR _18348_/B sky130_fd_sc_hd__or2_4
XANTENNA__15679__A _12713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22495__B1 _15831_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15559_ _14283_/A _23115_/Q VGND VGND VPWR VPWR _15559_/X sky130_fd_sc_hd__or2_4
XFILLER_33_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14583__A _15028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18163__B2 _18162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18278_ _18332_/A _18330_/A _17517_/X VGND VGND VPWR VPWR _18278_/X sky130_fd_sc_hd__o21a_4
X_17229_ _16814_/B _17137_/X _15381_/X _17138_/X VGND VGND VPWR VPWR _17229_/X sky130_fd_sc_hd__o22a_4
XFILLER_11_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17894__A _17893_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13199__A _13004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20240_ _20492_/A VGND VGND VPWR VPWR _20240_/X sky130_fd_sc_hd__buf_2
XFILLER_102_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13927__A _13927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20171_ _20105_/A _20171_/B VGND VGND VPWR VPWR _20172_/B sky130_fd_sc_hd__and2_4
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12750__A3 _12732_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12831__A _12753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16303__A _12837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19816__A1_N _19531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23930_ _23706_/CLK _21231_/X VGND VGND VPWR VPWR _16404_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19614__A HRDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23861_ _24021_/CLK _21367_/X VGND VGND VPWR VPWR _12661_/B sky130_fd_sc_hd__dfxtp_4
X_22812_ _22792_/X _22812_/B VGND VGND VPWR VPWR HWDATA[12] sky130_fd_sc_hd__nor2_4
XANTENNA__23318__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13662__A _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23792_ _24047_/CLK _21475_/X VGND VGND VPWR VPWR _13341_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21525__A2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22743_ SYSTICKCLKDIV[5] VGND VGND VPWR VPWR _22743_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12278__A _13025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22674_ _21795_/A _22672_/X _23100_/Q _22669_/X VGND VGND VPWR VPWR _23100_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23468__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24413_ _24435_/CLK _24413_/D HRESETn VGND VGND VPWR VPWR _20296_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21625_ _21565_/X _21619_/X _14502_/B _21623_/X VGND VGND VPWR VPWR _21625_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14493__A _14492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24344_ _24344_/CLK _18970_/X HRESETn VGND VGND VPWR VPWR _24344_/Q sky130_fd_sc_hd__dfstp_4
X_21556_ _21556_/A VGND VGND VPWR VPWR _21556_/X sky130_fd_sc_hd__buf_2
XANTENNA__24329__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20507_ _24212_/Q _20398_/X _20506_/Y VGND VGND VPWR VPWR _22413_/A sky130_fd_sc_hd__o21a_4
X_24275_ _23326_/CLK _19258_/X HRESETn VGND VGND VPWR VPWR _24275_/Q sky130_fd_sc_hd__dfrtp_4
X_21487_ _21275_/X _21484_/X _13829_/B _21481_/X VGND VGND VPWR VPWR _21487_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23226_ _23313_/CLK _22477_/X VGND VGND VPWR VPWR _16430_/B sky130_fd_sc_hd__dfxtp_4
X_20438_ _24247_/Q _20421_/X _20437_/X VGND VGND VPWR VPWR _20438_/X sky130_fd_sc_hd__o21a_4
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22215__A _22222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14940__B _14882_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_48_0_HCLK clkbuf_6_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_48_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23157_ _23157_/CLK _22584_/X VGND VGND VPWR VPWR _12620_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17309__A _14723_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21461__B2 _21460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20369_ _20209_/X _20359_/Y _20367_/X _20368_/Y _20233_/X VGND VGND VPWR VPWR _20369_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12741__A _15820_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22108_ _22108_/A VGND VGND VPWR VPWR _22108_/X sky130_fd_sc_hd__buf_2
X_23088_ _23920_/CLK _23088_/D VGND VGND VPWR VPWR _13340_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_62_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20016__A2 _17672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14930_ _12340_/A _14866_/B VGND VGND VPWR VPWR _14930_/X sky130_fd_sc_hd__or2_4
X_22039_ _21816_/X _22038_/X _12980_/B _22035_/X VGND VGND VPWR VPWR _22039_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19524__A _19481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21764__A2 _21762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23046__A _23051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14861_ _12216_/A _14859_/X _14861_/C VGND VGND VPWR VPWR _14861_/X sky130_fd_sc_hd__and3_4
XFILLER_48_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16600_ _11692_/X VGND VGND VPWR VPWR _16621_/A sky130_fd_sc_hd__buf_2
XANTENNA__13572__A _13572_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13812_ _13624_/A _13812_/B _13812_/C VGND VGND VPWR VPWR _13813_/C sky130_fd_sc_hd__and3_4
Xclkbuf_4_3_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17580_ _17101_/X VGND VGND VPWR VPWR _18107_/A sky130_fd_sc_hd__buf_2
XFILLER_21_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14792_ _12575_/A _14790_/X _14791_/X VGND VGND VPWR VPWR _14793_/C sky130_fd_sc_hd__and3_4
XANTENNA__21516__A2 _21508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22713__B2 _22668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16531_ _16536_/A _23740_/Q VGND VGND VPWR VPWR _16532_/C sky130_fd_sc_hd__or2_4
XANTENNA__13291__B _13291_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13743_ _13711_/X _13741_/X _13742_/X VGND VGND VPWR VPWR _13743_/X sky130_fd_sc_hd__and3_4
XFILLER_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19250_ _24279_/Q _19251_/A _19249_/Y VGND VGND VPWR VPWR _19250_/X sky130_fd_sc_hd__o21a_4
X_16462_ _16363_/X _16457_/X _16462_/C VGND VGND VPWR VPWR _16462_/X sky130_fd_sc_hd__or3_4
XFILLER_31_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13674_ _15442_/A _13674_/B _13673_/X VGND VGND VPWR VPWR _13674_/X sky130_fd_sc_hd__or3_4
XFILLER_32_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18201_ _18199_/X _18200_/X _18199_/X _18200_/X VGND VGND VPWR VPWR _19382_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15413_ _15413_/A _23916_/Q VGND VGND VPWR VPWR _15415_/B sky130_fd_sc_hd__or2_4
X_12625_ _12948_/A _12625_/B _12624_/X VGND VGND VPWR VPWR _12625_/X sky130_fd_sc_hd__or3_4
X_19181_ _19181_/A VGND VGND VPWR VPWR _19181_/Y sky130_fd_sc_hd__inv_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22477__B1 _16430_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16393_ _16121_/A _16389_/X _16393_/C VGND VGND VPWR VPWR _16393_/X sky130_fd_sc_hd__or3_4
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12916__A _13009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18132_ _18174_/C _18174_/D _18132_/C VGND VGND VPWR VPWR _18132_/X sky130_fd_sc_hd__and3_4
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12556_ _12556_/A _12556_/B _12555_/X VGND VGND VPWR VPWR _12556_/X sky130_fd_sc_hd__or3_4
X_15344_ _14009_/A _15342_/X _15344_/C VGND VGND VPWR VPWR _15344_/X sky130_fd_sc_hd__and3_4
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11507_ _19092_/A _11506_/Y VGND VGND VPWR VPWR _11508_/B sky130_fd_sc_hd__or2_4
XFILLER_32_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18063_ _18063_/A VGND VGND VPWR VPWR _18267_/A sky130_fd_sc_hd__buf_2
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15011__B _23551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12487_ _13022_/A VGND VGND VPWR VPWR _13031_/A sky130_fd_sc_hd__buf_2
X_15275_ _14994_/A _15273_/X _15274_/X VGND VGND VPWR VPWR _15279_/B sky130_fd_sc_hd__and3_4
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17014_ _17014_/A VGND VGND VPWR VPWR _17014_/X sky130_fd_sc_hd__buf_2
X_14226_ _14182_/A _23945_/Q VGND VGND VPWR VPWR _14227_/C sky130_fd_sc_hd__or2_4
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22125__A _22125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14157_ _15006_/A VGND VGND VPWR VPWR _14158_/A sky130_fd_sc_hd__buf_2
XFILLER_119_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13747__A _13747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13108_ _13080_/A _24050_/Q VGND VGND VPWR VPWR _13109_/C sky130_fd_sc_hd__or2_4
XFILLER_119_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14088_ _14083_/A _23177_/Q VGND VGND VPWR VPWR _14088_/X sky130_fd_sc_hd__or2_4
X_18965_ _18965_/A VGND VGND VPWR VPWR _18965_/X sky130_fd_sc_hd__buf_2
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13039_ _13016_/A _13039_/B VGND VGND VPWR VPWR _13040_/C sky130_fd_sc_hd__or2_4
X_17916_ _17916_/A VGND VGND VPWR VPWR _17916_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18896_ _13270_/X _18891_/X _19010_/A _18892_/X VGND VGND VPWR VPWR _24369_/D sky130_fd_sc_hd__o22a_4
XFILLER_117_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17847_ _17814_/X _17229_/X _17815_/X _17217_/X VGND VGND VPWR VPWR _17847_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14578__A _14145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20963__B1 _20576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13482__A _13442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17778_ _18240_/A VGND VGND VPWR VPWR _18063_/A sky130_fd_sc_hd__buf_2
XFILLER_19_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22795__A _18720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19517_ _19517_/A VGND VGND VPWR VPWR _19672_/D sky130_fd_sc_hd__buf_2
X_16729_ _12068_/X _16729_/B _16729_/C VGND VGND VPWR VPWR _16729_/X sky130_fd_sc_hd__and3_4
XFILLER_81_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23610__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12098__A _12098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16793__A _16747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22180__A2 _22179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19448_ _19419_/X _19445_/X _18016_/X _19447_/X VGND VGND VPWR VPWR _24190_/D sky130_fd_sc_hd__o22a_4
XFILLER_91_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21204__A _21168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19379_ _18652_/A VGND VGND VPWR VPWR _19379_/X sky130_fd_sc_hd__buf_2
XANTENNA__12826__A _12826_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21410_ _21229_/X _21405_/X _16421_/B _21409_/X VGND VGND VPWR VPWR _23834_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15202__A _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22390_ _20314_/A VGND VGND VPWR VPWR _22390_/X sky130_fd_sc_hd__buf_2
X_21341_ _21282_/X _21340_/X _14688_/B _21337_/X VGND VGND VPWR VPWR _23876_/D sky130_fd_sc_hd__o22a_4
XFILLER_11_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24060_ _24092_/CLK _24060_/D VGND VGND VPWR VPWR _24060_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24399__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21272_ _21270_/X _21271_/X _23913_/Q _21266_/X VGND VGND VPWR VPWR _21272_/X sky130_fd_sc_hd__o22a_4
XFILLER_2_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24116__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22035__A _22035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23011_ _22989_/A _23008_/Y _23011_/C VGND VGND VPWR VPWR _23011_/X sky130_fd_sc_hd__and3_4
XANTENNA__18232__B _16999_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20223_ _20223_/A HRDATA[15] VGND VGND VPWR VPWR _20223_/X sky130_fd_sc_hd__or2_4
XANTENNA__13657__A _15431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21443__B2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12561__A _13770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17111__A2 _17032_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21994__A2 _21988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15122__A1 _14918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20154_ _20137_/Y _20138_/Y _11551_/X _20153_/X VGND VGND VPWR VPWR _20154_/X sky130_fd_sc_hd__o22a_4
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15122__B2 _15121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15872__A _13500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23140__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20085_ _19884_/X _20084_/X _19303_/X _17724_/X VGND VGND VPWR VPWR _24115_/D sky130_fd_sc_hd__a22oi_4
XANTENNA__13684__A1 _13594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21746__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23913_ _23561_/CLK _21272_/X VGND VGND VPWR VPWR _23913_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15591__B _15530_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23844_ _23907_/CLK _23844_/D VGND VGND VPWR VPWR _14635_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23775_ _23217_/CLK _23775_/D VGND VGND VPWR VPWR _23775_/Q sky130_fd_sc_hd__dfxtp_4
X_20987_ _20841_/X _20986_/X VGND VGND VPWR VPWR _20987_/X sky130_fd_sc_hd__and2_4
XFILLER_26_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22171__A2 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22726_ _19909_/A _22714_/X _23064_/B _22721_/Y VGND VGND VPWR VPWR _24104_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20182__A1 _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21114__A _21118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22657_ _22621_/A VGND VGND VPWR VPWR _22657_/X sky130_fd_sc_hd__buf_2
XANTENNA__12736__A _15693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12410_ _12419_/A _12329_/B VGND VGND VPWR VPWR _12411_/C sky130_fd_sc_hd__or2_4
XFILLER_40_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21608_ _21536_/X _21605_/X _13141_/B _21602_/X VGND VGND VPWR VPWR _23729_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15112__A _15105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13390_ _12822_/A _13381_/X _13389_/X VGND VGND VPWR VPWR _13391_/C sky130_fd_sc_hd__and3_4
Xclkbuf_4_11_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22588_ _22418_/X _22586_/X _13089_/B _22583_/X VGND VGND VPWR VPWR _23154_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12341_ _12341_/A VGND VGND VPWR VPWR _13726_/A sky130_fd_sc_hd__buf_2
X_21539_ _21527_/A VGND VGND VPWR VPWR _21539_/X sky130_fd_sc_hd__buf_2
X_24327_ _24305_/CLK _24327_/D HRESETn VGND VGND VPWR VPWR _19065_/A sky130_fd_sc_hd__dfstp_4
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21682__B2 _21637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15060_ _12341_/A _23167_/Q VGND VGND VPWR VPWR _15062_/B sky130_fd_sc_hd__or2_4
X_12272_ _13054_/A _12270_/X _12271_/X VGND VGND VPWR VPWR _12278_/B sky130_fd_sc_hd__and3_4
X_24258_ _24321_/CLK _19292_/X HRESETn VGND VGND VPWR VPWR _24258_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14011_ _14813_/A _14011_/B VGND VGND VPWR VPWR _14011_/X sky130_fd_sc_hd__or2_4
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23209_ _23433_/CLK _22501_/X VGND VGND VPWR VPWR _23209_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13567__A _13500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21434__B2 _21430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22631__B1 _16131_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24189_ _24165_/CLK _19492_/Y HRESETn VGND VGND VPWR VPWR _17343_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18750_ _18750_/A _18750_/B _18327_/A _18750_/D VGND VGND VPWR VPWR _18751_/C sky130_fd_sc_hd__or4_4
XANTENNA__15782__A _15712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15962_ _15986_/A _15960_/X _15961_/X VGND VGND VPWR VPWR _15962_/X sky130_fd_sc_hd__and3_4
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21198__B1 _23945_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17701_ _16974_/A _17354_/X _16974_/A _17354_/X VGND VGND VPWR VPWR _17701_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14913_ _15011_/A _23840_/Q VGND VGND VPWR VPWR _14914_/C sky130_fd_sc_hd__or2_4
X_18681_ _18681_/A _18556_/X VGND VGND VPWR VPWR _18681_/X sky130_fd_sc_hd__and2_4
X_15893_ _13529_/X _15893_/B _15892_/X VGND VGND VPWR VPWR _15893_/X sky130_fd_sc_hd__and3_4
XANTENNA__23633__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17632_ _17261_/X _18746_/A _18107_/A _17631_/X VGND VGND VPWR VPWR _17633_/B sky130_fd_sc_hd__o22a_4
XFILLER_97_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14844_ _14021_/A _14772_/B VGND VGND VPWR VPWR _14846_/B sky130_fd_sc_hd__or2_4
XFILLER_17_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17563_ _17560_/Y _17015_/X _17022_/X _17653_/B VGND VGND VPWR VPWR _17564_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22698__B1 _15573_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11534__B IRQ[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14775_ _13647_/A _14771_/X _14774_/X VGND VGND VPWR VPWR _14775_/X sky130_fd_sc_hd__or3_4
XFILLER_63_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11987_ _11962_/X _11781_/B VGND VGND VPWR VPWR _11988_/C sky130_fd_sc_hd__or2_4
XFILLER_95_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19302_ _19317_/A VGND VGND VPWR VPWR _19302_/X sky130_fd_sc_hd__buf_2
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19563__B1 HRDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16514_ _16513_/X VGND VGND VPWR VPWR _16514_/X sky130_fd_sc_hd__buf_2
XFILLER_72_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13726_ _13726_/A VGND VGND VPWR VPWR _13735_/A sky130_fd_sc_hd__buf_2
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23783__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17494_ _17490_/Y _17493_/Y VGND VGND VPWR VPWR _17495_/A sky130_fd_sc_hd__or2_4
XANTENNA__21370__B1 _23859_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14845__B _14773_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19233_ _24284_/Q _19233_/B VGND VGND VPWR VPWR _19234_/B sky130_fd_sc_hd__and2_4
X_16445_ _11702_/A _16380_/B VGND VGND VPWR VPWR _16445_/X sky130_fd_sc_hd__or2_4
X_13657_ _15431_/A _13655_/X _13656_/X VGND VGND VPWR VPWR _13658_/C sky130_fd_sc_hd__and3_4
XANTENNA__16118__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12646__A _12646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15022__A _14588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12608_ _12963_/A _12604_/X _12607_/X VGND VGND VPWR VPWR _12609_/C sky130_fd_sc_hd__and3_4
X_19164_ _24306_/Q _19165_/A _19163_/Y VGND VGND VPWR VPWR _24306_/D sky130_fd_sc_hd__o21a_4
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21959__A _21919_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16376_ _16377_/B VGND VGND VPWR VPWR _16376_/X sky130_fd_sc_hd__buf_2
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13588_ _13588_/A VGND VGND VPWR VPWR _15927_/B sky130_fd_sc_hd__inv_2
XFILLER_9_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18115_ _18114_/X VGND VGND VPWR VPWR _18115_/Y sky130_fd_sc_hd__inv_2
X_15327_ _15332_/A _15262_/B VGND VGND VPWR VPWR _15329_/B sky130_fd_sc_hd__or2_4
X_12539_ _12500_/X _12653_/B VGND VGND VPWR VPWR _12540_/C sky130_fd_sc_hd__or2_4
X_19095_ _18965_/A _19093_/X _19094_/Y _19084_/X VGND VGND VPWR VPWR _19095_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22870__B1 _17339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19429__A _19429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18046_ _18425_/A _17993_/X _18425_/A _17990_/X VGND VGND VPWR VPWR _18046_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15258_ _14145_/A _15254_/X _15257_/X VGND VGND VPWR VPWR _15258_/X sky130_fd_sc_hd__or3_4
XFILLER_12_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24375__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14580__B _14662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14209_ _14218_/A VGND VGND VPWR VPWR _14210_/A sky130_fd_sc_hd__buf_2
XANTENNA__21425__B2 _21423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15189_ _15201_/A _15128_/B VGND VGND VPWR VPWR _15189_/X sky130_fd_sc_hd__or2_4
XANTENNA__21976__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_31_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19997_ _18169_/X _19985_/X _19995_/Y _19996_/X VGND VGND VPWR VPWR _19997_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15692__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18948_ _18937_/X _18947_/X _18937_/X _24348_/Q VGND VGND VPWR VPWR _18948_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21728__A2 _21726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18879_ _11837_/X _18875_/X _24382_/Q _18878_/X VGND VGND VPWR VPWR _24382_/D sky130_fd_sc_hd__o22a_4
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20910_ _20910_/A VGND VGND VPWR VPWR _20910_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21890_ _21821_/X _21887_/X _23569_/Q _21884_/X VGND VGND VPWR VPWR _21890_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20841_ _20214_/Y VGND VGND VPWR VPWR _20841_/X sky130_fd_sc_hd__buf_2
XFILLER_39_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18508__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23560_ _23304_/CLK _21903_/X VGND VGND VPWR VPWR _23560_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20772_ _18528_/X _20653_/X _20758_/X _20771_/Y VGND VGND VPWR VPWR _20773_/A sky130_fd_sc_hd__a211o_4
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22511_ _22458_/X _22507_/X _15243_/B _22476_/A VGND VGND VPWR VPWR _23201_/D sky130_fd_sc_hd__o22a_4
XFILLER_39_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21900__A2 _21894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23491_ _23907_/CLK _23491_/D VGND VGND VPWR VPWR _14788_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12556__A _12556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22442_ _22127_/A VGND VGND VPWR VPWR _22442_/X sky130_fd_sc_hd__buf_2
XANTENNA__21869__A _21884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22373_ _22131_/X _22368_/X _14279_/B _22372_/X VGND VGND VPWR VPWR _23270_/D sky130_fd_sc_hd__o22a_4
XFILLER_30_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15867__A _13546_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21664__B2 _21659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14771__A _13800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18243__A _18297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_113_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR _24088_/CLK sky130_fd_sc_hd__clkbuf_1
X_24112_ _24199_/CLK _20131_/Y HRESETn VGND VGND VPWR VPWR _24112_/Q sky130_fd_sc_hd__dfrtp_4
X_21324_ _21253_/X _21319_/X _13318_/B _21323_/X VGND VGND VPWR VPWR _21324_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15586__B _23339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24043_ _23688_/CLK _21042_/X VGND VGND VPWR VPWR _15556_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21255_ _21253_/X _21247_/X _13308_/B _21254_/X VGND VGND VPWR VPWR _23920_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12291__A _12695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20206_ _20206_/A _17025_/A VGND VGND VPWR VPWR _20206_/X sky130_fd_sc_hd__or2_4
XFILLER_89_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21186_ _20574_/X _21183_/X _23953_/Q _21180_/X VGND VGND VPWR VPWR _23953_/D sky130_fd_sc_hd__o22a_4
XFILLER_46_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23656__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20137_ _24430_/Q VGND VGND VPWR VPWR _20137_/Y sky130_fd_sc_hd__inv_2
X_20068_ _19379_/X _16998_/A _20048_/X _20067_/X VGND VGND VPWR VPWR _20069_/A sky130_fd_sc_hd__o22a_4
X_11910_ _15578_/A VGND VGND VPWR VPWR _11911_/A sky130_fd_sc_hd__buf_2
XFILLER_98_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15107__A _15107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12890_ _12890_/A _12888_/X _12890_/C VGND VGND VPWR VPWR _12890_/X sky130_fd_sc_hd__and3_4
XANTENNA__14011__A _14813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11841_ _11841_/A VGND VGND VPWR VPWR _11842_/A sky130_fd_sc_hd__buf_2
X_23827_ _23827_/CLK _23827_/D VGND VGND VPWR VPWR _23827_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18418__A _18418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22144__A2 _22137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17322__A _15381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11772_ _16215_/A VGND VGND VPWR VPWR _11772_/X sky130_fd_sc_hd__buf_2
X_14560_ _13747_/A _14556_/X _14560_/C VGND VGND VPWR VPWR _14561_/C sky130_fd_sc_hd__or3_4
XFILLER_57_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23758_ _23922_/CLK _23758_/D VGND VGND VPWR VPWR _15722_/B sky130_fd_sc_hd__dfxtp_4
X_13511_ _12951_/A VGND VGND VPWR VPWR _13511_/X sky130_fd_sc_hd__buf_2
X_22709_ _21855_/A _22707_/X _14776_/B _22704_/X VGND VGND VPWR VPWR _23075_/D sky130_fd_sc_hd__o22a_4
X_14491_ _13026_/A _14468_/X _14475_/X _14482_/X _14490_/X VGND VGND VPWR VPWR _14491_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12466__A _12917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23689_ _23847_/CLK _23689_/D VGND VGND VPWR VPWR _23689_/Q sky130_fd_sc_hd__dfxtp_4
X_16230_ _16180_/A _16230_/B _16230_/C VGND VGND VPWR VPWR _16231_/C sky130_fd_sc_hd__and3_4
XFILLER_70_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13442_ _12466_/X VGND VGND VPWR VPWR _13442_/X sky130_fd_sc_hd__buf_2
XFILLER_70_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15582__A1 _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13373_ _13383_/A _23568_/Q VGND VGND VPWR VPWR _13374_/C sky130_fd_sc_hd__or2_4
X_16161_ _16194_/A _16158_/X _16161_/C VGND VGND VPWR VPWR _16161_/X sky130_fd_sc_hd__and3_4
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15777__A _12672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23186__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_24_0_HCLK_A clkbuf_5_24_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18153__A _18153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15112_ _15105_/A _23199_/Q VGND VGND VPWR VPWR _15112_/X sky130_fd_sc_hd__or2_4
X_12324_ _12739_/A _12424_/B VGND VGND VPWR VPWR _12325_/C sky130_fd_sc_hd__or2_4
X_16092_ _16127_/A _16092_/B VGND VGND VPWR VPWR _16094_/B sky130_fd_sc_hd__or2_4
XFILLER_114_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12255_ _12709_/A VGND VGND VPWR VPWR _12255_/X sky130_fd_sc_hd__buf_2
X_15043_ _11611_/A _23679_/Q VGND VGND VPWR VPWR _15045_/B sky130_fd_sc_hd__or2_4
X_19920_ _19916_/X _24145_/Q _19917_/X _20539_/B VGND VGND VPWR VPWR _19920_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21407__B2 _21402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21958__A2 _21952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19851_ _19818_/A _19730_/D VGND VGND VPWR VPWR _19851_/X sky130_fd_sc_hd__or2_4
XFILLER_9_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12186_ _12115_/X _12186_/B VGND VGND VPWR VPWR _12186_/X sky130_fd_sc_hd__or2_4
XANTENNA__22080__B2 _22072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_18_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22403__A _20418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18802_ _18788_/A VGND VGND VPWR VPWR _18802_/X sky130_fd_sc_hd__buf_2
X_19782_ _19494_/X _19771_/X _19781_/X VGND VGND VPWR VPWR _19782_/X sky130_fd_sc_hd__o21a_4
XFILLER_95_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16994_ _24190_/Q VGND VGND VPWR VPWR _17889_/A sky130_fd_sc_hd__inv_2
XFILLER_7_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18733_ _17862_/A _18732_/X _18183_/X _18368_/X VGND VGND VPWR VPWR _18733_/X sky130_fd_sc_hd__o22a_4
XFILLER_114_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15945_ _15952_/A _23768_/Q VGND VGND VPWR VPWR _15946_/C sky130_fd_sc_hd__or2_4
XFILLER_23_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18664_ _18160_/A _18658_/X _18660_/X _18662_/Y _18663_/X VGND VGND VPWR VPWR _18664_/X
+ sky130_fd_sc_hd__a32o_4
X_15876_ _15876_/A _23885_/Q VGND VGND VPWR VPWR _15876_/X sky130_fd_sc_hd__or2_4
X_17615_ _17610_/Y _17614_/X _17326_/X VGND VGND VPWR VPWR _17615_/X sky130_fd_sc_hd__o21a_4
X_14827_ _13851_/A _23811_/Q VGND VGND VPWR VPWR _14828_/C sky130_fd_sc_hd__or2_4
XANTENNA__22776__C _20196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18595_ _18557_/X VGND VGND VPWR VPWR _18595_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22135__A2 _22125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13760__A _12652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17546_ _17542_/Y _17015_/X _17022_/X _17646_/B VGND VGND VPWR VPWR _17549_/B sky130_fd_sc_hd__o22a_4
X_14758_ _14758_/A _14758_/B VGND VGND VPWR VPWR _14758_/X sky130_fd_sc_hd__or2_4
XFILLER_17_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13709_ _13709_/A VGND VGND VPWR VPWR _13710_/A sky130_fd_sc_hd__buf_2
XFILLER_36_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17477_ _13493_/X VGND VGND VPWR VPWR _17477_/Y sky130_fd_sc_hd__inv_2
X_14689_ _14672_/A _14689_/B VGND VGND VPWR VPWR _14689_/X sky130_fd_sc_hd__or2_4
XFILLER_60_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19216_ _19216_/A _19216_/B VGND VGND VPWR VPWR _19217_/B sky130_fd_sc_hd__and2_4
X_16428_ _16397_/X _24090_/Q VGND VGND VPWR VPWR _16428_/X sky130_fd_sc_hd__or2_4
X_19147_ _19135_/X VGND VGND VPWR VPWR _19147_/Y sky130_fd_sc_hd__inv_2
X_16359_ _11702_/A _16296_/B VGND VGND VPWR VPWR _16361_/B sky130_fd_sc_hd__or2_4
XANTENNA__21646__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18063__A _18063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14591__A _14161_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19078_ _19076_/Y _19077_/Y _11511_/B VGND VGND VPWR VPWR _19078_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12823__B _12823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18029_ _18421_/A VGND VGND VPWR VPWR _18137_/A sky130_fd_sc_hd__buf_2
XANTENNA__13000__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21040_ _20697_/X _21037_/X _15490_/B _21034_/X VGND VGND VPWR VPWR _21040_/X sky130_fd_sc_hd__o22a_4
XFILLER_47_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17407__A _14073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22991_ _22990_/X VGND VGND VPWR VPWR HADDR[18] sky130_fd_sc_hd__inv_2
XFILLER_80_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22374__A2 _22368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21942_ _21935_/A VGND VGND VPWR VPWR _21942_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_38_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR _23365_/CLK sky130_fd_sc_hd__clkbuf_1
X_21873_ _21887_/A VGND VGND VPWR VPWR _21873_/X sky130_fd_sc_hd__buf_2
XFILLER_110_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14766__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22126__A2 _22125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13670__A _13670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _20226_/A _20823_/X _20617_/X VGND VGND VPWR VPWR _20824_/Y sky130_fd_sc_hd__o21ai_4
X_23612_ _23515_/CLK _23612_/D VGND VGND VPWR VPWR _23612_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20755_ _20641_/X _20753_/X _20755_/C VGND VGND VPWR VPWR _20755_/X sky130_fd_sc_hd__and3_4
X_23543_ _23539_/CLK _23543_/D VGND VGND VPWR VPWR _23543_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12286__A _12211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21885__B2 _21884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24454__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23474_ _23986_/CLK _22040_/X VGND VGND VPWR VPWR _23474_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20686_ _20303_/X VGND VGND VPWR VPWR _20686_/X sky130_fd_sc_hd__buf_2
XFILLER_50_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22425_ _20610_/A VGND VGND VPWR VPWR _22425_/X sky130_fd_sc_hd__buf_2
XANTENNA__15597__A _15643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22356_ _22103_/X _22354_/X _23282_/Q _22351_/X VGND VGND VPWR VPWR _22356_/X sky130_fd_sc_hd__o22a_4
X_21307_ _21225_/X _21305_/X _23900_/Q _21302_/X VGND VGND VPWR VPWR _21307_/X sky130_fd_sc_hd__o22a_4
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22287_ _22124_/X _22286_/X _23337_/Q _22283_/X VGND VGND VPWR VPWR _23337_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12040_ _16713_/A _12118_/B VGND VGND VPWR VPWR _12040_/X sky130_fd_sc_hd__or2_4
X_24026_ _24026_/CLK _24026_/D VGND VGND VPWR VPWR _16390_/B sky130_fd_sc_hd__dfxtp_4
X_21238_ _21237_/X _21235_/X _16181_/B _21230_/X VGND VGND VPWR VPWR _21238_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22062__B2 _22056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17317__A _17143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21169_ _21183_/A VGND VGND VPWR VPWR _21169_/X sky130_fd_sc_hd__buf_2
XFILLER_104_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23038__B _23038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13991_ _13991_/A VGND VGND VPWR VPWR _14071_/A sky130_fd_sc_hd__buf_2
XFILLER_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15730_ _15725_/A _15674_/B VGND VGND VPWR VPWR _15730_/X sky130_fd_sc_hd__or2_4
X_12942_ _12949_/A _23923_/Q VGND VGND VPWR VPWR _12942_/X sky130_fd_sc_hd__or2_4
XFILLER_46_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21573__B1 _15260_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15661_ _12688_/A _15661_/B _15661_/C VGND VGND VPWR VPWR _15665_/B sky130_fd_sc_hd__and3_4
X_12873_ _13032_/A VGND VGND VPWR VPWR _12874_/A sky130_fd_sc_hd__buf_2
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17400_ _24165_/Q VGND VGND VPWR VPWR _22017_/B sky130_fd_sc_hd__buf_2
XFILLER_2_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19518__B1 HRDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14612_ _14727_/A _14610_/X _14612_/C VGND VGND VPWR VPWR _14612_/X sky130_fd_sc_hd__and3_4
X_11824_ _11824_/A _11820_/X _11823_/X VGND VGND VPWR VPWR _11835_/B sky130_fd_sc_hd__or3_4
X_18380_ _11628_/X VGND VGND VPWR VPWR _18381_/A sky130_fd_sc_hd__buf_2
X_15592_ _15592_/A _15590_/X _15591_/X VGND VGND VPWR VPWR _15592_/X sky130_fd_sc_hd__and3_4
XFILLER_37_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14395__B _14305_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17221_/Y _17130_/A VGND VGND VPWR VPWR _17331_/X sky130_fd_sc_hd__and2_4
X_14543_ _14519_/X _14473_/B VGND VGND VPWR VPWR _14543_/X sky130_fd_sc_hd__or2_4
XFILLER_18_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11754_/X VGND VGND VPWR VPWR _11818_/A sky130_fd_sc_hd__buf_2
XANTENNA__12196__A _12196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18741__A1 _12031_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _17262_/A _17561_/B VGND VGND VPWR VPWR _17262_/X sky130_fd_sc_hd__and2_4
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14474_ _12494_/A _14474_/B _14473_/X VGND VGND VPWR VPWR _14475_/C sky130_fd_sc_hd__and3_4
XFILLER_70_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11686_ _12421_/A VGND VGND VPWR VPWR _13231_/A sky130_fd_sc_hd__buf_2
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19001_ _18988_/X _19000_/X _18988_/X _11524_/A VGND VGND VPWR VPWR _19001_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16213_ _16162_/X _16211_/X _16212_/X VGND VGND VPWR VPWR _16213_/X sky130_fd_sc_hd__and3_4
XFILLER_35_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13425_ _11658_/X _13425_/B _13424_/X VGND VGND VPWR VPWR _13425_/X sky130_fd_sc_hd__and3_4
XANTENNA__23821__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21302__A _21301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17193_ _17192_/Y _17161_/X _13278_/X _17138_/X VGND VGND VPWR VPWR _17193_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21628__B2 _21623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16144_ _16130_/A _16144_/B _16143_/X VGND VGND VPWR VPWR _16144_/X sky130_fd_sc_hd__or3_4
X_13356_ _13351_/X _13353_/X _13356_/C VGND VGND VPWR VPWR _13356_/X sky130_fd_sc_hd__and3_4
XFILLER_115_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12307_ _12307_/A VGND VGND VPWR VPWR _12747_/A sky130_fd_sc_hd__buf_2
XFILLER_114_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16075_ _16180_/A _16075_/B _16074_/X VGND VGND VPWR VPWR _16075_/X sky130_fd_sc_hd__and3_4
X_13287_ _13286_/X _13287_/B VGND VGND VPWR VPWR _13287_/X sky130_fd_sc_hd__or2_4
X_15026_ _15026_/A _23103_/Q VGND VGND VPWR VPWR _15028_/B sky130_fd_sc_hd__or2_4
X_19903_ _22723_/A VGND VGND VPWR VPWR _19903_/X sky130_fd_sc_hd__buf_2
X_12238_ _15447_/A VGND VGND VPWR VPWR _12238_/X sky130_fd_sc_hd__buf_2
XANTENNA__22053__B2 _22049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13755__A _12612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12169_ _12169_/A _12169_/B _12168_/X VGND VGND VPWR VPWR _12169_/X sky130_fd_sc_hd__and3_4
X_19834_ _19775_/Y _19826_/B _19817_/C _19703_/A VGND VGND VPWR VPWR _19834_/X sky130_fd_sc_hd__o22a_4
XFILLER_96_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17480__A1 _17477_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17480__B2 _17479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16977_ _17680_/A _16977_/B VGND VGND VPWR VPWR _16978_/B sky130_fd_sc_hd__or2_4
X_19765_ _19759_/B _19765_/B VGND VGND VPWR VPWR _19766_/B sky130_fd_sc_hd__or2_4
XANTENNA__22356__A2 _22354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15970__A _15948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15928_ _15928_/A VGND VGND VPWR VPWR _15928_/X sky130_fd_sc_hd__buf_2
X_18716_ _18728_/B _18716_/B VGND VGND VPWR VPWR _18716_/X sky130_fd_sc_hd__and2_4
XFILLER_77_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19696_ _19683_/X _19759_/B _19581_/X _19695_/Y VGND VGND VPWR VPWR _19696_/X sky130_fd_sc_hd__a211o_4
XANTENNA__20367__A1 _18000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21564__B1 _14276_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17232__A1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18647_ _17742_/X _17743_/B _17729_/X VGND VGND VPWR VPWR _18647_/X sky130_fd_sc_hd__o21a_4
X_15859_ _13572_/A _15851_/X _15858_/X VGND VGND VPWR VPWR _15859_/X sky130_fd_sc_hd__and3_4
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19509__B1 HRDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13490__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18578_ _18578_/A _17606_/X VGND VGND VPWR VPWR _18578_/X sky130_fd_sc_hd__or2_4
X_17529_ _17156_/Y _17523_/Y _17476_/C _17528_/X VGND VGND VPWR VPWR _17530_/A sky130_fd_sc_hd__o22a_4
XFILLER_75_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20540_ _20229_/A _20539_/X _20284_/X VGND VGND VPWR VPWR _20540_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_32_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16743__B1 _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20471_ _20471_/A VGND VGND VPWR VPWR _20521_/B sky130_fd_sc_hd__buf_2
XANTENNA__12834__A _12769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22210_ _22079_/X _22208_/X _16657_/B _22205_/X VGND VGND VPWR VPWR _23388_/D sky130_fd_sc_hd__o22a_4
XFILLER_101_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23190_ _23313_/CLK _23190_/D VGND VGND VPWR VPWR _12228_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21095__A2 _21089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22292__B2 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12553__B _12660_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22141_ _22456_/A VGND VGND VPWR VPWR _22141_/X sky130_fd_sc_hd__buf_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22044__A1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22072_ _22071_/X VGND VGND VPWR VPWR _22072_/X sky130_fd_sc_hd__buf_2
XFILLER_82_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22044__B2 _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18748__A1_N _17057_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18799__A1 _17178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21023_ _21030_/A VGND VGND VPWR VPWR _21023_/X sky130_fd_sc_hd__buf_2
XANTENNA__13665__A _12211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22595__A2 _22593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22978__A _22978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15880__A _15892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19748__B1 _20539_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22974_ _18375_/X _22950_/X VGND VGND VPWR VPWR _22974_/X sky130_fd_sc_hd__or2_4
XFILLER_83_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21925_ _21791_/X _21924_/X _23549_/Q _21921_/X VGND VGND VPWR VPWR _21925_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11913__A _12464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21856_ _21855_/X _21853_/X _14758_/B _21848_/X VGND VGND VPWR VPWR _23587_/D sky130_fd_sc_hd__o22a_4
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _20807_/A VGND VGND VPWR VPWR _20807_/Y sky130_fd_sc_hd__inv_2
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21787_ _21812_/A VGND VGND VPWR VPWR _21787_/X sky130_fd_sc_hd__buf_2
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21858__B2 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _11540_/A IRQ[0] VGND VGND VPWR VPWR _11540_/X sky130_fd_sc_hd__and2_4
X_23526_ _23781_/CLK _23526_/D VGND VGND VPWR VPWR _14289_/B sky130_fd_sc_hd__dfxtp_4
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20738_ _20733_/X _20737_/X _24330_/Q _20686_/X VGND VGND VPWR VPWR _20738_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20530__A1 _18256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20669_ _24205_/Q _20614_/X _20668_/X VGND VGND VPWR VPWR _20670_/A sky130_fd_sc_hd__o21a_4
X_23457_ _23391_/CLK _22063_/X VGND VGND VPWR VPWR _15240_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12744__A _12744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ _13214_/A _13210_/B _13210_/C VGND VGND VPWR VPWR _13210_/X sky130_fd_sc_hd__and3_4
XANTENNA__23994__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15120__A _14918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22408_ _20463_/A VGND VGND VPWR VPWR _22408_/X sky130_fd_sc_hd__buf_2
XFILLER_32_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14190_ _14190_/A _14190_/B _14190_/C VGND VGND VPWR VPWR _14190_/X sky130_fd_sc_hd__or3_4
X_23388_ _23100_/CLK _23388_/D VGND VGND VPWR VPWR _16657_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12463__B _12463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13141_ _12240_/X _13141_/B VGND VGND VPWR VPWR _13141_/X sky130_fd_sc_hd__or2_4
XFILLER_30_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22339_ _22368_/A VGND VGND VPWR VPWR _22354_/A sky130_fd_sc_hd__buf_2
XANTENNA__19338__A2_N _18432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13072_ _13101_/A _13072_/B _13071_/X VGND VGND VPWR VPWR _13072_/X sky130_fd_sc_hd__or3_4
XFILLER_69_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12023_ _11901_/X VGND VGND VPWR VPWR _12024_/A sky130_fd_sc_hd__buf_2
X_16900_ _15927_/B _16899_/X _16520_/X VGND VGND VPWR VPWR _16900_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24009_ _23494_/CLK _21097_/X VGND VGND VPWR VPWR _24009_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13575__A _13574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17880_ _17777_/X _17790_/Y _17872_/X _17876_/Y _17879_/X VGND VGND VPWR VPWR _17880_/X
+ sky130_fd_sc_hd__a32o_4
X_16831_ _16518_/X _16830_/X _16518_/X _16830_/X VGND VGND VPWR VPWR _16831_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13294__B _24016_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19550_ HRDATA[28] VGND VGND VPWR VPWR _20342_/B sky130_fd_sc_hd__buf_2
XANTENNA__15790__A _12458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16762_ _16597_/X _16753_/X _16761_/X VGND VGND VPWR VPWR _16762_/X sky130_fd_sc_hd__and3_4
X_13974_ _12209_/A _24074_/Q VGND VGND VPWR VPWR _13974_/X sky130_fd_sc_hd__or2_4
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18501_ _18499_/X _17601_/A _18500_/X VGND VGND VPWR VPWR _18501_/X sky130_fd_sc_hd__a21o_4
X_15713_ _15712_/X VGND VGND VPWR VPWR _15713_/Y sky130_fd_sc_hd__inv_2
X_12925_ _12958_/A _12925_/B VGND VGND VPWR VPWR _12925_/X sky130_fd_sc_hd__or2_4
X_19481_ _19481_/A _19481_/B VGND VGND VPWR VPWR _19481_/X sky130_fd_sc_hd__and2_4
X_16693_ _16713_/A _24027_/Q VGND VGND VPWR VPWR _16695_/B sky130_fd_sc_hd__or2_4
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12919__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20201__A _20279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18432_ _17753_/C _17753_/B _17753_/C _17753_/B VGND VGND VPWR VPWR _18432_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11823__A _11823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15644_ _11799_/A _15644_/B _15644_/C VGND VGND VPWR VPWR _15645_/C sky130_fd_sc_hd__or3_4
XFILLER_73_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_21_0_HCLK clkbuf_6_10_0_HCLK/X VGND VGND VPWR VPWR _24162_/CLK sky130_fd_sc_hd__clkbuf_1
X_12856_ _11912_/A VGND VGND VPWR VPWR _12859_/A sky130_fd_sc_hd__buf_2
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_84_0_HCLK clkbuf_6_42_0_HCLK/X VGND VGND VPWR VPWR _24435_/CLK sky130_fd_sc_hd__clkbuf_1
X_11807_ _11819_/A _24062_/Q VGND VGND VPWR VPWR _11808_/C sky130_fd_sc_hd__or2_4
X_18363_ _18362_/X VGND VGND VPWR VPWR _18363_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15575_ _12861_/A _15573_/X _15574_/X VGND VGND VPWR VPWR _15575_/X sky130_fd_sc_hd__and3_4
XANTENNA__21849__B2 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15014__B _23423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12787_ _12787_/A _12787_/B _12787_/C VGND VGND VPWR VPWR _12807_/B sky130_fd_sc_hd__and3_4
XFILLER_109_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _18587_/B _17608_/A VGND VGND VPWR VPWR _17315_/A sky130_fd_sc_hd__and2_4
XANTENNA__22510__A2 _22507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14526_ _13695_/X _22325_/A VGND VGND VPWR VPWR _14528_/B sky130_fd_sc_hd__or2_4
XANTENNA__17510__A _13278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _11738_/A VGND VGND VPWR VPWR _13706_/A sky130_fd_sc_hd__buf_2
X_18294_ _18239_/A _17512_/A VGND VGND VPWR VPWR _18294_/X sky130_fd_sc_hd__or2_4
XFILLER_109_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ _17825_/A VGND VGND VPWR VPWR _17911_/A sky130_fd_sc_hd__buf_2
X_14457_ _13608_/A _14520_/B VGND VGND VPWR VPWR _14458_/C sky130_fd_sc_hd__or2_4
X_11669_ _11669_/A VGND VGND VPWR VPWR _11670_/A sky130_fd_sc_hd__buf_2
XANTENNA__12654__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15030__A _15030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _12822_/A _13408_/B _13408_/C VGND VGND VPWR VPWR _13424_/B sky130_fd_sc_hd__and3_4
XANTENNA__22274__A1 _22103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17176_ _15648_/X _17131_/X _17175_/Y _17133_/X VGND VGND VPWR VPWR _17176_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22274__B2 _22269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14388_ _15628_/A _14388_/B _14387_/X VGND VGND VPWR VPWR _14389_/C sky130_fd_sc_hd__and3_4
XANTENNA__11565__A2 IRQ[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16127_ _16127_/A _23607_/Q VGND VGND VPWR VPWR _16129_/B sky130_fd_sc_hd__or2_4
XANTENNA__15965__A _15956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13339_ _13483_/A _13334_/X _13338_/X VGND VGND VPWR VPWR _13339_/X sky130_fd_sc_hd__or3_4
XANTENNA__19437__A HRDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18341__A _16977_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16058_ _16058_/A _16058_/B _16058_/C VGND VGND VPWR VPWR _16058_/X sky130_fd_sc_hd__and3_4
XFILLER_83_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15009_ _15032_/A _15009_/B _15009_/C VGND VGND VPWR VPWR _15009_/X sky130_fd_sc_hd__or3_4
XANTENNA__13485__A _12905_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22577__A2 _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19817_ _19442_/B _19793_/B _19817_/C VGND VGND VPWR VPWR _19817_/X sky130_fd_sc_hd__and3_4
XFILLER_110_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19748_ _19497_/X HRDATA[3] _20539_/B _19496_/X VGND VGND VPWR VPWR _19748_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_38_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19679_ _19419_/X _19677_/X _11599_/X _19678_/X VGND VGND VPWR VPWR _19679_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11733__A _16072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21710_ _21538_/X _21705_/X _23664_/Q _21709_/X VGND VGND VPWR VPWR _23664_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15205__A _14252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19900__A _22978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22690_ _22683_/A VGND VGND VPWR VPWR _22690_/X sky130_fd_sc_hd__buf_2
XFILLER_53_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21641_ _21662_/A VGND VGND VPWR VPWR _21641_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22501__A2 _22500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21572_ _21287_/A VGND VGND VPWR VPWR _21572_/X sky130_fd_sc_hd__buf_2
X_24360_ _24330_/CLK _24360_/D HRESETn VGND VGND VPWR VPWR _19062_/A sky130_fd_sc_hd__dfstp_4
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22038__A _22031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20523_ _20522_/X VGND VGND VPWR VPWR _20523_/Y sky130_fd_sc_hd__inv_2
X_23311_ _23311_/CLK _22315_/X VGND VGND VPWR VPWR _23311_/Q sky130_fd_sc_hd__dfxtp_4
X_24291_ _24290_/CLK _19194_/X HRESETn VGND VGND VPWR VPWR _19112_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_53_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12564__A _12965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20454_ _20322_/X _20452_/X _11527_/A _20453_/X VGND VGND VPWR VPWR _20454_/X sky130_fd_sc_hd__o22a_4
X_23242_ _24011_/CLK _23242_/D VGND VGND VPWR VPWR _13995_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21877__A _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20781__A HRDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23173_ _23557_/CLK _22556_/X VGND VGND VPWR VPWR _14505_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15875__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19347__A _19336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20385_ _20292_/X _20384_/X _19134_/A _20305_/X VGND VGND VPWR VPWR _20386_/B sky130_fd_sc_hd__o22a_4
XANTENNA__18251__A _17874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22124_ _20778_/A VGND VGND VPWR VPWR _22124_/X sky130_fd_sc_hd__buf_2
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22055_ _21845_/X _22052_/X _23463_/Q _22049_/X VGND VGND VPWR VPWR _23463_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11908__A _14998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20579__B2 _20449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21006_ _21296_/A VGND VGND VPWR VPWR _21112_/B sky130_fd_sc_hd__buf_2
XFILLER_43_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21240__A2 _21235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21528__B1 _12463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22957_ _22962_/A _18437_/Y VGND VGND VPWR VPWR _22957_/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12739__A _12739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12710_ _12710_/A _23156_/Q VGND VGND VPWR VPWR _12710_/X sky130_fd_sc_hd__or2_4
XANTENNA__15115__A _15115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11643__A _15114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21908_ _21901_/A VGND VGND VPWR VPWR _21908_/X sky130_fd_sc_hd__buf_2
X_13690_ _13690_/A VGND VGND VPWR VPWR _13880_/A sky130_fd_sc_hd__buf_2
X_22888_ _22888_/A _19414_/A VGND VGND VPWR VPWR _22980_/A sky130_fd_sc_hd__or2_4
XANTENNA__12458__B _12445_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12641_ _12982_/A _12639_/X _12641_/C VGND VGND VPWR VPWR _12641_/X sky130_fd_sc_hd__and3_4
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21839_ _21838_/X _21829_/X _23594_/Q _21836_/X VGND VGND VPWR VPWR _23594_/D sky130_fd_sc_hd__o22a_4
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14954__A _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15360_ _14009_/A _15360_/B _15359_/X VGND VGND VPWR VPWR _15360_/X sky130_fd_sc_hd__and3_4
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _12967_/A _12564_/X _12571_/X VGND VGND VPWR VPWR _12572_/X sky130_fd_sc_hd__and3_4
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20503__A1 _18222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15769__B _15769_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ _15536_/A _14311_/B VGND VGND VPWR VPWR _14313_/B sky130_fd_sc_hd__or2_4
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _24338_/Q _11522_/X VGND VGND VPWR VPWR _18996_/A sky130_fd_sc_hd__or2_4
X_23509_ _23315_/CLK _21986_/X VGND VGND VPWR VPWR _12571_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15291_ _12860_/A _15289_/X _15291_/C VGND VGND VPWR VPWR _15291_/X sky130_fd_sc_hd__and3_4
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17030_ _17024_/C _17030_/B _17009_/A _17285_/A VGND VGND VPWR VPWR _17033_/A sky130_fd_sc_hd__or4_4
X_14242_ _14190_/A _14237_/X _14242_/C VGND VGND VPWR VPWR _14242_/X sky130_fd_sc_hd__or3_4
XANTENNA__21787__A _21812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22256__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20691__A _24236_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24172__CLK _24299_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15785__A _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14173_ _12267_/X _14136_/X _14145_/X _14163_/X _14172_/X VGND VGND VPWR VPWR _14173_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18475__A3 _18471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13124_ _13100_/A _13124_/B _13123_/X VGND VGND VPWR VPWR _13124_/X sky130_fd_sc_hd__and3_4
XANTENNA__22008__B2 _22006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18981_ _18971_/X _18980_/X _18971_/X _11527_/A VGND VGND VPWR VPWR _24342_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22559__A2 _22557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13055_ _13055_/A _13051_/X _13055_/C VGND VGND VPWR VPWR _13055_/X sky130_fd_sc_hd__or3_4
X_17932_ _17932_/A VGND VGND VPWR VPWR _17932_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21767__B1 _15570_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12006_ _12112_/A _12006_/B _12005_/X VGND VGND VPWR VPWR _12006_/X sky130_fd_sc_hd__or3_4
XFILLER_79_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16238__A2 _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17863_ _17863_/A VGND VGND VPWR VPWR _17864_/A sky130_fd_sc_hd__buf_2
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22411__A _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19602_ _19598_/A _19599_/B VGND VGND VPWR VPWR _19638_/A sky130_fd_sc_hd__or2_4
X_16814_ _16743_/X _16814_/B VGND VGND VPWR VPWR _16815_/A sky130_fd_sc_hd__or2_4
X_17794_ _17794_/A VGND VGND VPWR VPWR _17794_/X sky130_fd_sc_hd__buf_2
XANTENNA__20990__B2 _20449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16745_ _16618_/X _23515_/Q VGND VGND VPWR VPWR _16746_/C sky130_fd_sc_hd__or2_4
X_19533_ _19450_/A VGND VGND VPWR VPWR _19793_/A sky130_fd_sc_hd__buf_2
XANTENNA__21027__A _21027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13957_ _13957_/A _13957_/B VGND VGND VPWR VPWR _13957_/X sky130_fd_sc_hd__and2_4
XANTENNA__12649__A _12951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12908_ _12872_/A _12980_/B VGND VGND VPWR VPWR _12910_/B sky130_fd_sc_hd__or2_4
X_19464_ _19742_/A VGND VGND VPWR VPWR _19464_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15025__A _14119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19720__A _19873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16676_ _16597_/X _16668_/X _16675_/X VGND VGND VPWR VPWR _16676_/X sky130_fd_sc_hd__and3_4
X_13888_ _13895_/A _23943_/Q VGND VGND VPWR VPWR _13888_/X sky130_fd_sc_hd__or2_4
XANTENNA__20742__A1 _18506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15627_ _15611_/A _15623_/X _15627_/C VGND VGND VPWR VPWR _15627_/X sky130_fd_sc_hd__or3_4
X_18415_ _24123_/Q _18414_/Y _16976_/B VGND VGND VPWR VPWR _22962_/B sky130_fd_sc_hd__o21a_4
X_12839_ _12787_/A _12831_/X _12839_/C VGND VGND VPWR VPWR _12839_/X sky130_fd_sc_hd__and3_4
X_19395_ _19392_/X _18439_/Y _19392_/X _24204_/Q VGND VGND VPWR VPWR _19395_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18346_ _16970_/A VGND VGND VPWR VPWR _18533_/A sky130_fd_sc_hd__buf_2
XANTENNA__17240__A _18249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15558_ _15558_/A _15554_/X _15557_/X VGND VGND VPWR VPWR _15558_/X sky130_fd_sc_hd__or3_4
XANTENNA__22495__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14509_ _14554_/A _14442_/B VGND VGND VPWR VPWR _14509_/X sky130_fd_sc_hd__or2_4
X_18277_ _18153_/Y _17513_/A _17516_/Y VGND VGND VPWR VPWR _18330_/A sky130_fd_sc_hd__o21a_4
X_15489_ _13735_/A _23596_/Q VGND VGND VPWR VPWR _15491_/B sky130_fd_sc_hd__or2_4
XANTENNA__12384__A _12958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17228_ _17144_/Y _17155_/X _17143_/X _17186_/X VGND VGND VPWR VPWR _17228_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22247__B2 _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17894__B _16977_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15695__A _15695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17159_ _17152_/X _17153_/X _17154_/X _17158_/X VGND VGND VPWR VPWR _17159_/X sky130_fd_sc_hd__o22a_4
X_20170_ _18940_/A _20169_/X VGND VGND VPWR VPWR _20171_/B sky130_fd_sc_hd__or2_4
XFILLER_115_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11728__A _11727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14104__A _14315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17415__A _14263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23860_ _24084_/CLK _21368_/X VGND VGND VPWR VPWR _23860_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22811_ _17339_/Y _22794_/X _22796_/X _22810_/X VGND VGND VPWR VPWR _22812_/B sky130_fd_sc_hd__o22a_4
XFILLER_38_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23791_ _23859_/CLK _21476_/X VGND VGND VPWR VPWR _13485_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24045__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22742_ SYSTICKCLKDIV[6] _22741_/A _22740_/Y _22741_/Y VGND VGND VPWR VPWR _22746_/C
+ sky130_fd_sc_hd__o22a_4
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22673_ _21791_/A _22672_/X _23101_/Q _22669_/X VGND VGND VPWR VPWR _23101_/D sky130_fd_sc_hd__o22a_4
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14774__A _13654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24412_ _24277_/CLK _24412_/D HRESETn VGND VGND VPWR VPWR _24412_/Q sky130_fd_sc_hd__dfrtp_4
X_21624_ _21562_/X _21619_/X _14272_/B _21623_/X VGND VGND VPWR VPWR _21624_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22991__A _22990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19351__B2 _20888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24343_ _24334_/CLK _18977_/X HRESETn VGND VGND VPWR VPWR _11528_/A sky130_fd_sc_hd__dfstp_4
X_21555_ _21555_/A VGND VGND VPWR VPWR _21555_/X sky130_fd_sc_hd__buf_2
XANTENNA__12294__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20506_ _20588_/A _20505_/X VGND VGND VPWR VPWR _20506_/Y sky130_fd_sc_hd__nand2_4
X_21486_ _21273_/X _21484_/X _13757_/B _21481_/X VGND VGND VPWR VPWR _21486_/X sky130_fd_sc_hd__o22a_4
X_24274_ _23326_/CLK _24274_/D HRESETn VGND VGND VPWR VPWR _19223_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22238__B2 _22233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20437_ _20376_/X _20423_/X _20288_/X _20436_/Y VGND VGND VPWR VPWR _20437_/X sky130_fd_sc_hd__a211o_4
X_23225_ _23130_/CLK _23225_/D VGND VGND VPWR VPWR _16289_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21997__B1 _23501_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20368_ _24250_/Q VGND VGND VPWR VPWR _20368_/Y sky130_fd_sc_hd__inv_2
X_23156_ _23157_/CLK _22585_/X VGND VGND VPWR VPWR _23156_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12741__B _12737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22107_ _20590_/A VGND VGND VPWR VPWR _22107_/X sky130_fd_sc_hd__buf_2
XANTENNA__11638__A _11638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23087_ _23859_/CLK _22692_/X VGND VGND VPWR VPWR _13484_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__19805__A _19877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20299_ _20407_/A _20296_/Y _20298_/X _18931_/A _20253_/X VGND VGND VPWR VPWR _20300_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14014__A _14021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22038_ _22031_/A VGND VGND VPWR VPWR _22038_/X sky130_fd_sc_hd__buf_2
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14949__A _15072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14860_ _13984_/A _14860_/B VGND VGND VPWR VPWR _14861_/C sky130_fd_sc_hd__or2_4
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17325__A _15251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13811_ _15430_/A _24039_/Q VGND VGND VPWR VPWR _13812_/C sky130_fd_sc_hd__or2_4
X_14791_ _13862_/A _14791_/B VGND VGND VPWR VPWR _14791_/X sky130_fd_sc_hd__or2_4
X_23989_ _24021_/CLK _21131_/X VGND VGND VPWR VPWR _12628_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_112_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12469__A _12518_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18917__A1 _15379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16530_ _16538_/A _16608_/B VGND VGND VPWR VPWR _16530_/X sky130_fd_sc_hd__or2_4
XANTENNA__22713__A2 _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13742_ _13697_/X _13652_/B VGND VGND VPWR VPWR _13742_/X sky130_fd_sc_hd__or2_4
XFILLER_16_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16461_ _16499_/A _16459_/X _16460_/X VGND VGND VPWR VPWR _16462_/C sky130_fd_sc_hd__and3_4
X_13673_ _13631_/A _13671_/X _13673_/C VGND VGND VPWR VPWR _13673_/X sky130_fd_sc_hd__and3_4
XFILLER_71_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14684__A _15592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18200_ _18174_/C _18174_/D _18174_/B VGND VGND VPWR VPWR _18200_/X sky130_fd_sc_hd__and3_4
X_15412_ _15412_/A _15408_/X _15412_/C VGND VGND VPWR VPWR _15412_/X sky130_fd_sc_hd__or3_4
X_12624_ _12947_/A _12620_/X _12623_/X VGND VGND VPWR VPWR _12624_/X sky130_fd_sc_hd__and3_4
X_19180_ _24298_/Q _19181_/A _19179_/Y VGND VGND VPWR VPWR _24298_/D sky130_fd_sc_hd__o21a_4
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16392_ _15948_/A _16390_/X _16391_/X VGND VGND VPWR VPWR _16393_/C sky130_fd_sc_hd__and3_4
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18131_ _24132_/Q _18132_/C _16984_/X VGND VGND VPWR VPWR _23016_/B sky130_fd_sc_hd__o21a_4
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19342__B2 _20743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15343_ _12567_/A _15343_/B VGND VGND VPWR VPWR _15344_/C sky130_fd_sc_hd__or2_4
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12555_ _13017_/A _12555_/B _12554_/X VGND VGND VPWR VPWR _12555_/X sky130_fd_sc_hd__and3_4
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23562__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11506_ _11506_/A VGND VGND VPWR VPWR _11506_/Y sky130_fd_sc_hd__inv_2
X_18062_ _18062_/A _17559_/A VGND VGND VPWR VPWR _18062_/X sky130_fd_sc_hd__or2_4
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15274_ _14165_/A _15274_/B VGND VGND VPWR VPWR _15274_/X sky130_fd_sc_hd__or2_4
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ _13622_/A VGND VGND VPWR VPWR _13022_/A sky130_fd_sc_hd__buf_2
XFILLER_89_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22406__A _20441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17013_ _17013_/A VGND VGND VPWR VPWR _17014_/A sky130_fd_sc_hd__buf_2
X_14225_ _14225_/A _23881_/Q VGND VGND VPWR VPWR _14227_/B sky130_fd_sc_hd__or2_4
XFILLER_32_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12932__A _12958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14156_ _15013_/A VGND VGND VPWR VPWR _15006_/A sky130_fd_sc_hd__buf_2
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13107_ _13119_/A _23602_/Q VGND VGND VPWR VPWR _13109_/B sky130_fd_sc_hd__or2_4
XFILLER_84_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14087_ _13956_/A VGND VGND VPWR VPWR _14136_/A sky130_fd_sc_hd__buf_2
X_18964_ _18994_/A VGND VGND VPWR VPWR _18965_/A sky130_fd_sc_hd__buf_2
XFILLER_80_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13038_ _13015_/A _23378_/Q VGND VGND VPWR VPWR _13040_/B sky130_fd_sc_hd__or2_4
X_17915_ _17817_/X _17207_/X _17825_/X _17189_/X VGND VGND VPWR VPWR _17916_/A sky130_fd_sc_hd__o22a_4
XFILLER_26_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17773__A1_N _11629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18895_ _13274_/X _18891_/X _24370_/Q _18892_/X VGND VGND VPWR VPWR _18895_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22141__A _22456_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13763__A _12935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17846_ _17845_/X VGND VGND VPWR VPWR _17846_/X sky130_fd_sc_hd__buf_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14989_ _14121_/A _15052_/B VGND VGND VPWR VPWR _14991_/B sky130_fd_sc_hd__or2_4
X_17777_ _18062_/A _17270_/X VGND VGND VPWR VPWR _17777_/X sky130_fd_sc_hd__or2_4
XANTENNA__12379__A _13211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18908__A1 _14261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24335__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22795__B _18752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19516_ _19516_/A VGND VGND VPWR VPWR _19861_/A sky130_fd_sc_hd__buf_2
XFILLER_93_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16728_ _12065_/X _24091_/Q VGND VGND VPWR VPWR _16729_/C sky130_fd_sc_hd__or2_4
XANTENNA__21912__B1 _23553_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16659_ _16640_/X _16657_/X _16659_/C VGND VGND VPWR VPWR _16659_/X sky130_fd_sc_hd__and3_4
X_19447_ _19678_/A VGND VGND VPWR VPWR _19447_/X sky130_fd_sc_hd__buf_2
XFILLER_62_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14594__A _15037_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18066__A _18066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_54_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19378_ _19378_/A VGND VGND VPWR VPWR _19378_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18329_ _17483_/X _18274_/C VGND VGND VPWR VPWR _18329_/X sky130_fd_sc_hd__or2_4
XANTENNA__15202__B _23553_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21340_ _21300_/A VGND VGND VPWR VPWR _21340_/X sky130_fd_sc_hd__buf_2
X_21271_ _21271_/A VGND VGND VPWR VPWR _21271_/X sky130_fd_sc_hd__buf_2
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13938__A _13959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16314__A _16185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12842__A _12752_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20222_ _20214_/Y _20618_/B VGND VGND VPWR VPWR _20226_/A sky130_fd_sc_hd__and2_4
X_23010_ _18193_/X _23017_/B VGND VGND VPWR VPWR _23011_/C sky130_fd_sc_hd__or2_4
XANTENNA__21443__A2 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16033__B _15967_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20153_ _20139_/Y _20140_/Y _11549_/X _20152_/X VGND VGND VPWR VPWR _20153_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19625__A _19866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20084_ _19957_/X _20082_/X _20083_/X _18602_/Y _19931_/B VGND VGND VPWR VPWR _20084_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_58_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14769__A _15413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23912_ _23079_/CLK _21274_/X VGND VGND VPWR VPWR _13723_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13673__A _13631_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22986__A _23015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23843_ _23270_/CLK _23843_/D VGND VGND VPWR VPWR _14780_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12289__A _12725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23774_ _23774_/CLK _23774_/D VGND VGND VPWR VPWR _21498_/A sky130_fd_sc_hd__dfxtp_4
X_20986_ _20842_/X _20984_/X _20985_/X HRDATA[8] _20847_/X VGND VGND VPWR VPWR _20986_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22725_ _22898_/A _22724_/X _19201_/X _19380_/X VGND VGND VPWR VPWR _22725_/X sky130_fd_sc_hd__o22a_4
XFILLER_26_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20182__A2 _16997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22656_ _22449_/X _22650_/X _14539_/B _22654_/X VGND VGND VPWR VPWR _22656_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22459__B2 _22386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16208__B _16131_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21607_ _21534_/X _21605_/X _23730_/Q _21602_/X VGND VGND VPWR VPWR _21607_/X sky130_fd_sc_hd__o22a_4
XFILLER_16_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15112__B _23199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22587_ _22415_/X _22586_/X _12945_/B _22583_/X VGND VGND VPWR VPWR _22587_/X sky130_fd_sc_hd__o22a_4
XFILLER_90_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14009__A _14009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21131__B2 _21130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12340_ _12340_/A VGND VGND VPWR VPWR _12341_/A sky130_fd_sc_hd__buf_2
X_24326_ _24305_/CLK _24326_/D HRESETn VGND VGND VPWR VPWR _11511_/A sky130_fd_sc_hd__dfstp_4
X_21538_ _20591_/A VGND VGND VPWR VPWR _21538_/X sky130_fd_sc_hd__buf_2
XANTENNA__17886__B2 _11629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21682__A2 _21662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22226__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21130__A _21130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12271_ _12240_/A _12271_/B VGND VGND VPWR VPWR _12271_/X sky130_fd_sc_hd__or2_4
X_24257_ _24321_/CLK _19294_/X HRESETn VGND VGND VPWR VPWR _24257_/Q sky130_fd_sc_hd__dfrtp_4
X_21469_ _21244_/X _21463_/X _23796_/Q _21467_/X VGND VGND VPWR VPWR _21469_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12752__A _12751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14010_ _14010_/A VGND VGND VPWR VPWR _14813_/A sky130_fd_sc_hd__buf_2
X_23208_ _23304_/CLK _23208_/D VGND VGND VPWR VPWR _13766_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21434__A2 _21433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24188_ _24165_/CLK _24188_/D HRESETn VGND VGND VPWR VPWR _17412_/A sky130_fd_sc_hd__dfrtp_4
X_23139_ _23433_/CLK _23139_/D VGND VGND VPWR VPWR _23139_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24210__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15961_ _15957_/A _23544_/Q VGND VGND VPWR VPWR _15961_/X sky130_fd_sc_hd__or2_4
XFILLER_1_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15782__B _15782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23057__A _19953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14679__A _14679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21198__B2 _21194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14912_ _14912_/A _14912_/B VGND VGND VPWR VPWR _14914_/B sky130_fd_sc_hd__or2_4
X_17700_ _17699_/X _17375_/X _17696_/B VGND VGND VPWR VPWR _17753_/B sky130_fd_sc_hd__a21bo_4
XFILLER_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15892_ _15892_/A _15836_/B VGND VGND VPWR VPWR _15892_/X sky130_fd_sc_hd__or2_4
X_18680_ _18679_/X VGND VGND VPWR VPWR _18680_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14398__B _14308_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14843_ _12575_/A _14841_/X _14842_/X VGND VGND VPWR VPWR _14843_/X sky130_fd_sc_hd__and3_4
X_17631_ _17267_/X _17630_/X _17785_/B VGND VGND VPWR VPWR _17631_/X sky130_fd_sc_hd__o21a_4
XFILLER_5_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12199__A _12198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17562_ _17039_/X _17561_/X _17043_/X VGND VGND VPWR VPWR _17653_/B sky130_fd_sc_hd__o21ai_4
XFILLER_1_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14774_ _13654_/A _14774_/B _14774_/C VGND VGND VPWR VPWR _14774_/X sky130_fd_sc_hd__and3_4
XFILLER_40_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11986_ _11983_/A _11779_/B VGND VGND VPWR VPWR _11986_/X sky130_fd_sc_hd__or2_4
XFILLER_16_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22698__B2 _22697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16513_ _11658_/X _16513_/B _16513_/C VGND VGND VPWR VPWR _16513_/X sky130_fd_sc_hd__and3_4
X_19301_ _22888_/A VGND VGND VPWR VPWR _19317_/A sky130_fd_sc_hd__buf_2
X_13725_ _13765_/A _13723_/X _13725_/C VGND VGND VPWR VPWR _13725_/X sky130_fd_sc_hd__and3_4
XFILLER_75_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21305__A _21319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17493_ _17492_/X VGND VGND VPWR VPWR _17493_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12927__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21370__B2 _21366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11831__A _11821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16444_ _16443_/X VGND VGND VPWR VPWR _16444_/Y sky130_fd_sc_hd__inv_2
X_19232_ _19232_/A _19231_/X VGND VGND VPWR VPWR _19233_/B sky130_fd_sc_hd__and2_4
XANTENNA__15303__A _14588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13656_ _13630_/A _13745_/B VGND VGND VPWR VPWR _13656_/X sky130_fd_sc_hd__or2_4
XANTENNA__16118__B _16186_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12607_ _12643_/A _12607_/B VGND VGND VPWR VPWR _12607_/X sky130_fd_sc_hd__or2_4
X_19163_ _19163_/A VGND VGND VPWR VPWR _19163_/Y sky130_fd_sc_hd__inv_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16375_ _16374_/X VGND VGND VPWR VPWR _16377_/B sky130_fd_sc_hd__inv_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ _12432_/X _12678_/Y _12434_/A _13586_/Y VGND VGND VPWR VPWR _13588_/A sky130_fd_sc_hd__a211o_4
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21122__B2 _21116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18114_ _17962_/A _18110_/X _17836_/A _18113_/X VGND VGND VPWR VPWR _18114_/X sky130_fd_sc_hd__o22a_4
X_15326_ _14178_/A VGND VGND VPWR VPWR _15332_/A sky130_fd_sc_hd__buf_2
X_12538_ _12497_/X _12651_/B VGND VGND VPWR VPWR _12540_/B sky130_fd_sc_hd__or2_4
X_19094_ _19094_/A VGND VGND VPWR VPWR _19094_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22136__A _20892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18045_ _17242_/A VGND VGND VPWR VPWR _18425_/A sky130_fd_sc_hd__buf_2
X_15257_ _11909_/A _15255_/X _15256_/X VGND VGND VPWR VPWR _15257_/X sky130_fd_sc_hd__and3_4
XANTENNA__13758__A _15495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12469_ _12518_/A VGND VGND VPWR VPWR _12868_/A sky130_fd_sc_hd__buf_2
XANTENNA__23308__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12662__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14208_ _14247_/A _23145_/Q VGND VGND VPWR VPWR _14208_/X sky130_fd_sc_hd__or2_4
XANTENNA__21425__A2 _21419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15188_ _14183_/A _15186_/X _15188_/C VGND VGND VPWR VPWR _15188_/X sky130_fd_sc_hd__and3_4
XFILLER_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12381__B _12248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20633__B1 _20632_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14139_ _14138_/X _23113_/Q VGND VGND VPWR VPWR _14141_/B sky130_fd_sc_hd__or2_4
XFILLER_10_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19445__A _19445_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16301__A1 _11982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19996_ _19996_/A VGND VGND VPWR VPWR _19996_/X sky130_fd_sc_hd__buf_2
XFILLER_113_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18947_ _18941_/X _18943_/X _18944_/Y _18946_/X VGND VGND VPWR VPWR _18947_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14589__A _14588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21189__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18878_ _18892_/A VGND VGND VPWR VPWR _18878_/X sky130_fd_sc_hd__buf_2
XFILLER_67_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17829_ _17825_/X _17827_/X _17806_/X _17828_/X VGND VGND VPWR VPWR _17829_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20840_ _20750_/X _20838_/X _14320_/B _20839_/X VGND VGND VPWR VPWR _20840_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22689__A1 _20574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22689__B2 _22683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20771_ _20715_/A _20771_/B VGND VGND VPWR VPWR _20771_/Y sky130_fd_sc_hd__nor2_4
XFILLER_39_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12837__A _12837_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21361__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22510_ _22456_/X _22507_/X _15299_/B _22504_/X VGND VGND VPWR VPWR _23202_/D sky130_fd_sc_hd__o22a_4
XFILLER_50_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15213__A _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11741__A _12613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23490_ _23907_/CLK _23490_/D VGND VGND VPWR VPWR _15253_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18109__A2 _17919_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22441_ _22439_/X _22440_/X _14078_/B _22435_/X VGND VGND VPWR VPWR _23241_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22372_ _22351_/A VGND VGND VPWR VPWR _22372_/X sky130_fd_sc_hd__buf_2
XANTENNA__21664__A2 _21662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24111_ _24199_/CLK _20179_/Y HRESETn VGND VGND VPWR VPWR _18681_/A sky130_fd_sc_hd__dfrtp_4
X_21323_ _21316_/A VGND VGND VPWR VPWR _21323_/X sky130_fd_sc_hd__buf_2
XANTENNA__13668__A _15436_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12572__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16044__A _16215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24233__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21254_ _21242_/A VGND VGND VPWR VPWR _21254_/X sky130_fd_sc_hd__buf_2
X_24042_ _23915_/CLK _24042_/D VGND VGND VPWR VPWR _24042_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22613__B2 _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20205_ _20399_/A VGND VGND VPWR VPWR _20370_/A sky130_fd_sc_hd__buf_2
XANTENNA__15883__A _15876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21185_ _20553_/X _21183_/X _23954_/Q _21180_/X VGND VGND VPWR VPWR _23954_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19355__A _19370_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20136_ IRQ[17] VGND VGND VPWR VPWR _20136_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14854__A1 _14786_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24131__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20067_ _18573_/X _20057_/X _20066_/Y _19929_/X VGND VGND VPWR VPWR _20067_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20927__A1 _20403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14606__A1 _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11840_ _11839_/X VGND VGND VPWR VPWR _11841_/A sky130_fd_sc_hd__buf_2
X_23826_ _23826_/CLK _23826_/D VGND VGND VPWR VPWR _13112_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11771_ _11770_/X VGND VGND VPWR VPWR _16215_/A sky130_fd_sc_hd__buf_2
X_23757_ _23922_/CLK _23757_/D VGND VGND VPWR VPWR _15792_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20969_ _20425_/A _20965_/X _20967_/X _20968_/Y _20473_/A VGND VGND VPWR VPWR _20970_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12747__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24381__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16219__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13510_ _12413_/X _13508_/X _13510_/C VGND VGND VPWR VPWR _13510_/X sky130_fd_sc_hd__and3_4
X_22708_ _21282_/A _22707_/X _14703_/B _22704_/X VGND VGND VPWR VPWR _22708_/X sky130_fd_sc_hd__o22a_4
X_14490_ _13597_/X _14490_/B VGND VGND VPWR VPWR _14490_/X sky130_fd_sc_hd__and2_4
X_23688_ _23688_/CLK _23688_/D VGND VGND VPWR VPWR _13759_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13441_ _13483_/A _13436_/X _13441_/C VGND VGND VPWR VPWR _13441_/X sky130_fd_sc_hd__or3_4
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22882__C _22932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22639_ _22420_/X _22636_/X _13178_/B _22633_/X VGND VGND VPWR VPWR _23121_/D sky130_fd_sc_hd__o22a_4
XFILLER_107_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21104__B2 _21100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16160_ _16159_/X _23511_/Q VGND VGND VPWR VPWR _16161_/C sky130_fd_sc_hd__or2_4
XFILLER_31_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13372_ _13358_/X _13308_/B VGND VGND VPWR VPWR _13372_/X sky130_fd_sc_hd__or2_4
X_15111_ _15107_/A _15109_/X _15110_/X VGND VGND VPWR VPWR _15115_/B sky130_fd_sc_hd__and3_4
X_12323_ _12738_/A _12323_/B VGND VGND VPWR VPWR _12323_/X sky130_fd_sc_hd__or2_4
X_24309_ _24301_/CLK _19158_/X HRESETn VGND VGND VPWR VPWR _24309_/Q sky130_fd_sc_hd__dfrtp_4
X_16091_ _16091_/A VGND VGND VPWR VPWR _16127_/A sky130_fd_sc_hd__buf_2
XFILLER_86_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15042_ _13955_/A _15040_/X _15042_/C VGND VGND VPWR VPWR _15042_/X sky130_fd_sc_hd__and3_4
XANTENNA__21795__A _21795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12254_ _13670_/A VGND VGND VPWR VPWR _12709_/A sky130_fd_sc_hd__buf_2
XANTENNA__16889__A _16822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15793__A _12859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19850_ _19849_/X VGND VGND VPWR VPWR _19850_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12185_ _12184_/X VGND VGND VPWR VPWR _12186_/B sky130_fd_sc_hd__inv_2
XANTENNA__18284__B2 _18283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18801_ _14425_/A _18795_/X _24422_/Q _18796_/X VGND VGND VPWR VPWR _24422_/D sky130_fd_sc_hd__o22a_4
X_19781_ _19580_/X _19772_/X _19774_/X _19780_/X VGND VGND VPWR VPWR _19781_/X sky130_fd_sc_hd__or4_4
X_16993_ _16937_/X _16991_/B _16992_/Y VGND VGND VPWR VPWR _16993_/X sky130_fd_sc_hd__a21o_4
XANTENNA__20204__A _16929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11826__A _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18732_ _17969_/X _18731_/X _17975_/X _18143_/X VGND VGND VPWR VPWR _18732_/X sky130_fd_sc_hd__o22a_4
X_15944_ _15939_/A _16019_/B VGND VGND VPWR VPWR _15944_/X sky130_fd_sc_hd__or2_4
XFILLER_42_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11545__B IRQ[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15875_ _11665_/X _15859_/X _15875_/C VGND VGND VPWR VPWR _15907_/B sky130_fd_sc_hd__or3_4
X_18663_ _18662_/A _18662_/B _17634_/X VGND VGND VPWR VPWR _18663_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19712__B HRDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14826_ _13872_/A _14762_/B VGND VGND VPWR VPWR _14826_/X sky130_fd_sc_hd__or2_4
X_17614_ _17611_/Y _17613_/Y _17329_/X VGND VGND VPWR VPWR _17614_/X sky130_fd_sc_hd__o21a_4
XFILLER_40_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18594_ _18593_/X VGND VGND VPWR VPWR _18594_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14757_ _12449_/A _14757_/B _14756_/X VGND VGND VPWR VPWR _14757_/X sky130_fd_sc_hd__and3_4
X_17545_ _17544_/X VGND VGND VPWR VPWR _17646_/B sky130_fd_sc_hd__inv_2
X_11969_ _12008_/A _11790_/B VGND VGND VPWR VPWR _11969_/X sky130_fd_sc_hd__or2_4
XFILLER_45_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16129__A _16109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21343__B2 _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13708_ _13708_/A VGND VGND VPWR VPWR _13709_/A sky130_fd_sc_hd__buf_2
XANTENNA__15033__A _13925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17476_ _18254_/A _17456_/Y _17476_/C _18191_/A VGND VGND VPWR VPWR _17476_/X sky130_fd_sc_hd__or4_4
X_14688_ _15105_/A _14688_/B VGND VGND VPWR VPWR _14690_/B sky130_fd_sc_hd__or2_4
XFILLER_32_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19215_ _19215_/A _19215_/B VGND VGND VPWR VPWR _19216_/B sky130_fd_sc_hd__and2_4
X_13639_ _12302_/A VGND VGND VPWR VPWR _13647_/A sky130_fd_sc_hd__buf_2
X_16427_ _16091_/A _16427_/B VGND VGND VPWR VPWR _16427_/X sky130_fd_sc_hd__or2_4
XFILLER_38_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15968__A _13477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16358_ _16303_/X _16356_/X _16358_/C VGND VGND VPWR VPWR _16358_/X sky130_fd_sc_hd__and3_4
X_19146_ _24315_/Q _19135_/X _19145_/Y VGND VGND VPWR VPWR _24315_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21646__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15309_ _14782_/A _15305_/X _15308_/X VGND VGND VPWR VPWR _15309_/X sky130_fd_sc_hd__or3_4
XFILLER_69_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16289_ _15939_/A _16289_/B VGND VGND VPWR VPWR _16291_/B sky130_fd_sc_hd__or2_4
X_19077_ _11510_/B VGND VGND VPWR VPWR _19077_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12392__A _12392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18028_ _17090_/X _17550_/B VGND VGND VPWR VPWR _18031_/C sky130_fd_sc_hd__nor2_4
XFILLER_114_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23280__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19979_ _19970_/X _17951_/A _19976_/X _19978_/X VGND VGND VPWR VPWR _19979_/X sky130_fd_sc_hd__o22a_4
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15208__A _15201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11736__A _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19903__A _22723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22990_ _22985_/X _17674_/A _22967_/X _22989_/X VGND VGND VPWR VPWR _22990_/X sky130_fd_sc_hd__a211o_4
XFILLER_68_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14112__A _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20909__A1 _18664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21941_ _21821_/X _21938_/X _23537_/Q _21935_/X VGND VGND VPWR VPWR _23537_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20385__A2 _20384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21872_ _21901_/A VGND VGND VPWR VPWR _21887_/A sky130_fd_sc_hd__buf_2
XFILLER_58_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _23515_/CLK _23611_/D VGND VGND VPWR VPWR _23611_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _20642_/X _20823_/B _20823_/C VGND VGND VPWR VPWR _20823_/X sky130_fd_sc_hd__and3_4
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12567__A _12567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21334__B2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22531__B1 _16096_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23542_ _23539_/CLK _21934_/X VGND VGND VPWR VPWR _12263_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20754_ _20754_/A _20754_/B VGND VGND VPWR VPWR _20755_/C sky130_fd_sc_hd__or2_4
XFILLER_23_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15878__A _12413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23473_ _23473_/CLK _22041_/X VGND VGND VPWR VPWR _23473_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20685_ _20622_/X _20684_/X _19217_/A _20497_/X VGND VGND VPWR VPWR _20685_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14782__A _14782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_24_0_HCLK clkbuf_5_24_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21098__B1 _24008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22424_ _22422_/X _22416_/X _13282_/B _22423_/X VGND VGND VPWR VPWR _22424_/X sky130_fd_sc_hd__o22a_4
X_22355_ _22100_/X _22354_/X _23283_/Q _22351_/X VGND VGND VPWR VPWR _22355_/X sky130_fd_sc_hd__o22a_4
X_21306_ _21221_/X _21305_/X _23901_/Q _21302_/X VGND VGND VPWR VPWR _21306_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24383__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22286_ _22286_/A VGND VGND VPWR VPWR _22286_/X sky130_fd_sc_hd__buf_2
XFILLER_105_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22504__A _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22598__B1 _23147_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24025_ _23514_/CLK _21074_/X VGND VGND VPWR VPWR _24025_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21237_ _20442_/A VGND VGND VPWR VPWR _21237_/X sky130_fd_sc_hd__buf_2
XANTENNA__22062__A2 _22059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19463__B1 HRDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16502__A _16203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16816__A2 _16814_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21168_ _21168_/A VGND VGND VPWR VPWR _21183_/A sky130_fd_sc_hd__buf_2
XANTENNA__20024__A _20000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20119_ _11547_/B _20117_/X _20118_/Y VGND VGND VPWR VPWR _20119_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15118__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13990_ _13989_/X VGND VGND VPWR VPWR _14074_/A sky130_fd_sc_hd__inv_2
X_21099_ _20819_/X _21096_/X _13859_/B _21093_/X VGND VGND VPWR VPWR _24007_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12941_ _13083_/A _12931_/X _12941_/C VGND VGND VPWR VPWR _12957_/B sky130_fd_sc_hd__and3_4
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14957__A _13998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21573__B2 _21563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13861__A _14810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15660_ _12286_/X _15722_/B VGND VGND VPWR VPWR _15661_/C sky130_fd_sc_hd__or2_4
X_12872_ _12872_/A _22311_/A VGND VGND VPWR VPWR _12875_/B sky130_fd_sc_hd__or2_4
XFILLER_73_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14611_ _11894_/A _14692_/B VGND VGND VPWR VPWR _14612_/C sky130_fd_sc_hd__or2_4
X_11823_ _11823_/A _11821_/X _11822_/X VGND VGND VPWR VPWR _11823_/X sky130_fd_sc_hd__and3_4
X_23809_ _23487_/CLK _23809_/D VGND VGND VPWR VPWR _23809_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15591_ _15584_/A _15530_/B VGND VGND VPWR VPWR _15591_/X sky130_fd_sc_hd__or2_4
XFILLER_2_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12477__A _13029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21325__B2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17330_ _17330_/A _17329_/X VGND VGND VPWR VPWR _17330_/X sky130_fd_sc_hd__and2_4
XFILLER_14_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _13695_/X _14472_/B VGND VGND VPWR VPWR _14544_/B sky130_fd_sc_hd__or2_4
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _16064_/A VGND VGND VPWR VPWR _11754_/X sky130_fd_sc_hd__buf_2
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17242_/A VGND VGND VPWR VPWR _17261_/X sky130_fd_sc_hd__buf_2
XANTENNA__15788__A _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _13020_/A _14473_/B VGND VGND VPWR VPWR _14473_/X sky130_fd_sc_hd__or2_4
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11684_/X VGND VGND VPWR VPWR _11685_/X sky130_fd_sc_hd__buf_2
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16212_ _16227_/A _16135_/B VGND VGND VPWR VPWR _16212_/X sky130_fd_sc_hd__or2_4
X_19000_ _18994_/X _18997_/X _18998_/Y _18999_/X VGND VGND VPWR VPWR _19000_/X sky130_fd_sc_hd__o22a_4
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ _11800_/X _13424_/B _13423_/X VGND VGND VPWR VPWR _13424_/X sky130_fd_sc_hd__or3_4
X_17192_ _17191_/X VGND VGND VPWR VPWR _17192_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21628__A2 _21626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16143_ _16143_/A _16143_/B _16143_/C VGND VGND VPWR VPWR _16143_/X sky130_fd_sc_hd__and3_4
XFILLER_10_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20836__B1 _20835_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13355_ _13354_/X _23504_/Q VGND VGND VPWR VPWR _13356_/C sky130_fd_sc_hd__or2_4
X_12306_ _15448_/A VGND VGND VPWR VPWR _12307_/A sky130_fd_sc_hd__buf_2
X_16074_ _11745_/X _16070_/X _16073_/X VGND VGND VPWR VPWR _16074_/X sky130_fd_sc_hd__or3_4
X_13286_ _15689_/A VGND VGND VPWR VPWR _13286_/X sky130_fd_sc_hd__buf_2
XFILLER_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15025_ _14119_/X _15021_/X _15024_/X VGND VGND VPWR VPWR _15025_/X sky130_fd_sc_hd__or3_4
X_19902_ _19901_/X VGND VGND VPWR VPWR _22723_/A sky130_fd_sc_hd__buf_2
X_12237_ _12209_/A VGND VGND VPWR VPWR _15447_/A sky130_fd_sc_hd__buf_2
XANTENNA__17508__A _13278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18257__B2 _18256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22053__A2 _22052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_44_0_HCLK clkbuf_6_22_0_HCLK/X VGND VGND VPWR VPWR _23910_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12940__A _12964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19833_ _19832_/X VGND VGND VPWR VPWR _19833_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12168_ _12168_/A _23805_/Q VGND VGND VPWR VPWR _12168_/X sky130_fd_sc_hd__or2_4
XFILLER_81_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16131__B _16131_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15028__A _15028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19764_ _19766_/A _19789_/B _19721_/Y VGND VGND VPWR VPWR _19764_/X sky130_fd_sc_hd__a21o_4
X_12099_ _12068_/X _12099_/B _12099_/C VGND VGND VPWR VPWR _12105_/B sky130_fd_sc_hd__and3_4
X_16976_ _17694_/A _16976_/B VGND VGND VPWR VPWR _16977_/B sky130_fd_sc_hd__or2_4
XFILLER_110_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20869__A _22134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18715_ _17782_/Y _18714_/X _17329_/X VGND VGND VPWR VPWR _18715_/X sky130_fd_sc_hd__o21a_4
XFILLER_7_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15927_ _15927_/A _15927_/B _15926_/X VGND VGND VPWR VPWR _15928_/A sky130_fd_sc_hd__and3_4
X_19695_ _19694_/X VGND VGND VPWR VPWR _19695_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21564__B2 _21563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13771__A _11799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18646_ _17006_/A _18641_/Y _16935_/A _18645_/X VGND VGND VPWR VPWR _18646_/X sky130_fd_sc_hd__o22a_4
XFILLER_65_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15858_ _15882_/A _15854_/X _15858_/C VGND VGND VPWR VPWR _15858_/X sky130_fd_sc_hd__or3_4
X_14809_ _13694_/A _14739_/B VGND VGND VPWR VPWR _14809_/X sky130_fd_sc_hd__or2_4
X_18577_ _16929_/X VGND VGND VPWR VPWR _18577_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12387__A _12386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15789_ _12859_/A _15787_/X _15789_/C VGND VGND VPWR VPWR _15790_/C sky130_fd_sc_hd__and3_4
XANTENNA__22513__B1 _23199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17528_ _18191_/A _17526_/X _17527_/Y VGND VGND VPWR VPWR _17528_/X sky130_fd_sc_hd__o21a_4
XFILLER_75_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15698__A _12737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17459_ _17688_/B VGND VGND VPWR VPWR _17459_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16743__A1 _11844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22816__A1 _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20470_ _20470_/A VGND VGND VPWR VPWR _20470_/Y sky130_fd_sc_hd__inv_2
X_19129_ _19129_/A _19129_/B VGND VGND VPWR VPWR _19129_/X sky130_fd_sc_hd__and2_4
XANTENNA__22292__A2 _22286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14107__A _14318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13011__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22140_ _22139_/X _22137_/X _14806_/B _22132_/X VGND VGND VPWR VPWR _22140_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13946__A _12509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22071_ _22108_/A VGND VGND VPWR VPWR _22071_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17418__A _14261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22044__A2 _22038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12850__A _12850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21022_ _20394_/X _21016_/X _24057_/Q _21020_/X VGND VGND VPWR VPWR _24057_/D sky130_fd_sc_hd__o22a_4
XFILLER_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_1_0_HCLK clkbuf_6_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19748__A1 _19497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15880__B _15818_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22973_ _17893_/X _16977_/B _22998_/A _18231_/Y VGND VGND VPWR VPWR _22975_/B sky130_fd_sc_hd__a211o_4
XFILLER_110_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14777__A _13960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13493__B1 _11596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23176__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18249__A _18249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13681__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21924_ _21938_/A VGND VGND VPWR VPWR _21924_/X sky130_fd_sc_hd__buf_2
XFILLER_112_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21855_ _21855_/A VGND VGND VPWR VPWR _21855_/X sky130_fd_sc_hd__buf_2
XFILLER_71_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12297__A _15685_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21307__B2 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _20654_/X _20803_/Y _20805_/X _19068_/Y _20709_/X VGND VGND VPWR VPWR _20807_/A
+ sky130_fd_sc_hd__a32o_4
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21858__A2 _21853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21786_ _21792_/A VGND VGND VPWR VPWR _21812_/A sky130_fd_sc_hd__inv_2
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23525_ _24008_/CLK _21958_/X VGND VGND VPWR VPWR _14450_/B sky130_fd_sc_hd__dfxtp_4
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19920__B2 _20539_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20737_ _20622_/X _20735_/X _19215_/A _20736_/X VGND VGND VPWR VPWR _20737_/X sky130_fd_sc_hd__o22a_4
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15401__A _12450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23456_ _23840_/CLK _23456_/D VGND VGND VPWR VPWR _23456_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20668_ _20534_/A _20667_/X VGND VGND VPWR VPWR _20668_/X sky130_fd_sc_hd__or2_4
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22407_ _22406_/X _22404_/X _16158_/B _22399_/X VGND VGND VPWR VPWR _22407_/X sky130_fd_sc_hd__o22a_4
XFILLER_32_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23387_ _23100_/CLK _23387_/D VGND VGND VPWR VPWR _16791_/B sky130_fd_sc_hd__dfxtp_4
X_20599_ _20598_/X VGND VGND VPWR VPWR _20599_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14017__A _12599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20961__B _20400_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13140_ _12693_/A _13140_/B VGND VGND VPWR VPWR _13140_/X sky130_fd_sc_hd__or2_4
X_22338_ _22332_/Y _22337_/X _22073_/X _22337_/X VGND VGND VPWR VPWR _23294_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13071_ _13128_/A _13071_/B _13070_/X VGND VGND VPWR VPWR _13071_/X sky130_fd_sc_hd__and3_4
XANTENNA__17328__A _14988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19436__B1 HRDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22269_ _22269_/A VGND VGND VPWR VPWR _22269_/X sky130_fd_sc_hd__buf_2
XFILLER_2_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16232__A _11658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12022_ _12022_/A _23710_/Q VGND VGND VPWR VPWR _12025_/B sky130_fd_sc_hd__or2_4
X_24008_ _24008_/CLK _21098_/X VGND VGND VPWR VPWR _24008_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21794__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16830_ _16519_/A _16829_/X _16377_/X VGND VGND VPWR VPWR _16830_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19543__A _19829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13973_ _13643_/A _23466_/Q VGND VGND VPWR VPWR _13975_/B sky130_fd_sc_hd__or2_4
X_16761_ _11834_/A _16756_/X _16761_/C VGND VGND VPWR VPWR _16761_/X sky130_fd_sc_hd__or3_4
XFILLER_20_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14687__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18500_ _18442_/A VGND VGND VPWR VPWR _18500_/X sky130_fd_sc_hd__buf_2
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12924_ _11842_/X _12681_/X _12893_/X _11596_/X _12923_/X VGND VGND VPWR VPWR _12924_/X
+ sky130_fd_sc_hd__a32o_4
X_15712_ _12189_/X _12681_/X _15681_/X _12281_/X _15711_/X VGND VGND VPWR VPWR _15712_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_47_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16692_ _16715_/A _16692_/B _16692_/C VGND VGND VPWR VPWR _16696_/B sky130_fd_sc_hd__and3_4
X_19480_ _19742_/A VGND VGND VPWR VPWR _19481_/A sky130_fd_sc_hd__buf_2
XFILLER_46_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18411__B2 _18410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12919__B _23859_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18431_ _18314_/X _18417_/Y _18357_/X _18430_/X VGND VGND VPWR VPWR _18431_/X sky130_fd_sc_hd__o22a_4
X_12855_ _12458_/A _12849_/X _12855_/C VGND VGND VPWR VPWR _12855_/X sky130_fd_sc_hd__or3_4
X_15643_ _15643_/A _15643_/B _15643_/C VGND VGND VPWR VPWR _15644_/C sky130_fd_sc_hd__and3_4
XFILLER_62_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11806_ _11818_/A _23614_/Q VGND VGND VPWR VPWR _11808_/B sky130_fd_sc_hd__or2_4
X_15574_ _15574_/A _23787_/Q VGND VGND VPWR VPWR _15574_/X sky130_fd_sc_hd__or2_4
X_18362_ _18244_/A _18362_/B _18360_/Y _18361_/X VGND VGND VPWR VPWR _18362_/X sky130_fd_sc_hd__or4_4
XANTENNA__21849__A2 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12786_ _12771_/X _12775_/X _12785_/X VGND VGND VPWR VPWR _12787_/C sky130_fd_sc_hd__or3_4
XANTENNA__12000__A _11943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14494_/X _14523_/X _14524_/X VGND VGND VPWR VPWR _14525_/X sky130_fd_sc_hd__and3_4
X_17313_ _14429_/B _17313_/B VGND VGND VPWR VPWR _17608_/A sky130_fd_sc_hd__nand2_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11737_/A VGND VGND VPWR VPWR _11738_/A sky130_fd_sc_hd__inv_2
XANTENNA__19911__B2 _20754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _18234_/B _22987_/B _18236_/B VGND VGND VPWR VPWR _18293_/X sky130_fd_sc_hd__o21a_4
XFILLER_30_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12935__A _12935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _15399_/A _14518_/B VGND VGND VPWR VPWR _14458_/B sky130_fd_sc_hd__or2_4
X_17244_ _17824_/A VGND VGND VPWR VPWR _17244_/X sky130_fd_sc_hd__buf_2
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _13991_/A VGND VGND VPWR VPWR _11669_/A sky130_fd_sc_hd__buf_2
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _11681_/X _13403_/X _13407_/C VGND VGND VPWR VPWR _13408_/C sky130_fd_sc_hd__or3_4
XFILLER_11_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17175_ _13274_/X VGND VGND VPWR VPWR _17175_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14387_ _15611_/A _14380_/X _14387_/C VGND VGND VPWR VPWR _14387_/X sky130_fd_sc_hd__or3_4
XANTENNA__22274__A2 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11599_ _11598_/X VGND VGND VPWR VPWR _11599_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16126_ _16140_/A _16126_/B _16126_/C VGND VGND VPWR VPWR _16130_/B sky130_fd_sc_hd__and3_4
XFILLER_115_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13338_ _13467_/A _13336_/X _13338_/C VGND VGND VPWR VPWR _13338_/X sky130_fd_sc_hd__and3_4
XANTENNA__21482__B1 _23787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16057_ _16050_/A _23416_/Q VGND VGND VPWR VPWR _16058_/C sky130_fd_sc_hd__or2_4
XANTENNA__13766__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13269_ _11656_/A _13237_/X _13268_/X VGND VGND VPWR VPWR _13270_/A sky130_fd_sc_hd__and3_4
XANTENNA__12670__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16142__A _16139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15008_ _14748_/A _15006_/X _15008_/C VGND VGND VPWR VPWR _15009_/C sky130_fd_sc_hd__and3_4
XFILLER_44_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22798__B _15051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19816_ _19531_/X _19815_/X _16913_/X _19531_/X VGND VGND VPWR VPWR _19816_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19747_ HRDATA[19] VGND VGND VPWR VPWR _20539_/B sky130_fd_sc_hd__buf_2
X_16959_ _24117_/Q VGND VGND VPWR VPWR _16969_/A sky130_fd_sc_hd__inv_2
XANTENNA__21537__A1 _21536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14597__A _13600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21537__B2 _21527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22734__B1 SYSTICKCLKDIV[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19678_ _19678_/A VGND VGND VPWR VPWR _19678_/X sky130_fd_sc_hd__buf_2
XFILLER_53_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12829__B _23860_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18629_ _17321_/Y _17616_/X VGND VGND VPWR VPWR _18629_/Y sky130_fd_sc_hd__nand2_4
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13006__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21640_ _21636_/A VGND VGND VPWR VPWR _21662_/A sky130_fd_sc_hd__buf_2
XANTENNA__21223__A _21247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21571_ _21570_/X _21568_/X _14733_/B _21563_/X VGND VGND VPWR VPWR _23747_/D sky130_fd_sc_hd__o22a_4
XFILLER_60_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23310_ _23692_/CLK _23310_/D VGND VGND VPWR VPWR _15669_/B sky130_fd_sc_hd__dfxtp_4
X_20522_ _20425_/X _20519_/Y _20521_/X _18998_/Y _20473_/X VGND VGND VPWR VPWR _20522_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_20_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24290_ _24290_/CLK _19196_/X HRESETn VGND VGND VPWR VPWR _19111_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_53_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23241_ _23978_/CLK _23241_/D VGND VGND VPWR VPWR _14078_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_20_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20453_ _20453_/A VGND VGND VPWR VPWR _20453_/X sky130_fd_sc_hd__buf_2
XFILLER_119_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23172_ _23107_/CLK _23172_/D VGND VGND VPWR VPWR _14661_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20384_ _20293_/X _20383_/X _11530_/A _20303_/X VGND VGND VPWR VPWR _20384_/X sky130_fd_sc_hd__o22a_4
XFILLER_106_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22123_ _22122_/X _22113_/X _14027_/B _22120_/X VGND VGND VPWR VPWR _23434_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12580__A _12980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22054_ _21843_/X _22052_/X _23464_/Q _22049_/X VGND VGND VPWR VPWR _23464_/D sky130_fd_sc_hd__o22a_4
XFILLER_62_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20579__A2 _20405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21005_ _21005_/A VGND VGND VPWR VPWR _21348_/A sky130_fd_sc_hd__buf_2
XFILLER_82_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_90_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR _23515_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_75_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23811__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21528__B2 _21527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22725__B1 _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11924__A _11924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22956_ _23015_/A VGND VGND VPWR VPWR _22982_/A sky130_fd_sc_hd__buf_2
XFILLER_60_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12739__B _12836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21907_ _21850_/X _21901_/X _14516_/B _21905_/X VGND VGND VPWR VPWR _23557_/D sky130_fd_sc_hd__o22a_4
XFILLER_71_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22887_ _22719_/X VGND VGND VPWR VPWR _22887_/X sky130_fd_sc_hd__buf_2
X_12640_ _12640_/A _12640_/B VGND VGND VPWR VPWR _12641_/C sky130_fd_sc_hd__or2_4
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21838_ _20748_/A VGND VGND VPWR VPWR _21838_/X sky130_fd_sc_hd__buf_2
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22229__A _22222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21133__A _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12571_ _12959_/A _12571_/B VGND VGND VPWR VPWR _12571_/X sky130_fd_sc_hd__or2_4
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21769_ _21740_/A VGND VGND VPWR VPWR _21769_/X sky130_fd_sc_hd__buf_2
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12755__A _13726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16227__A _16227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14310_ _15534_/A _14308_/X _14309_/X VGND VGND VPWR VPWR _14310_/X sky130_fd_sc_hd__and3_4
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21700__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11522_ _24337_/Q _19008_/A VGND VGND VPWR VPWR _11522_/X sky130_fd_sc_hd__or2_4
X_23508_ _23315_/CLK _21987_/X VGND VGND VPWR VPWR _23508_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15290_ _14152_/A _15290_/B VGND VGND VPWR VPWR _15291_/C sky130_fd_sc_hd__or2_4
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14241_ _14206_/A _14239_/X _14241_/C VGND VGND VPWR VPWR _14242_/C sky130_fd_sc_hd__and3_4
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23439_ _23859_/CLK _22111_/X VGND VGND VPWR VPWR _13457_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19657__B1 _19722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14172_ _14172_/A _14171_/X VGND VGND VPWR VPWR _14172_/X sky130_fd_sc_hd__and2_4
XANTENNA__15785__B _23501_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13123_ _13115_/A _13123_/B VGND VGND VPWR VPWR _13123_/X sky130_fd_sc_hd__or2_4
XANTENNA__22008__A2 _22002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19409__B1 _19380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18980_ _18965_/X _18978_/Y _18979_/Y _18968_/X VGND VGND VPWR VPWR _18980_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12490__A _13020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18880__A1 _12184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23341__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22899__A _23015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13054_ _13054_/A _13054_/B _13054_/C VGND VGND VPWR VPWR _13055_/C sky130_fd_sc_hd__and3_4
X_17931_ _17862_/X _17918_/X _17836_/X _17930_/X VGND VGND VPWR VPWR _17932_/A sky130_fd_sc_hd__o22a_4
XFILLER_79_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16897__A _16897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12005_ _11966_/X _12005_/B _12005_/C VGND VGND VPWR VPWR _12005_/X sky130_fd_sc_hd__and3_4
XFILLER_117_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21767__B2 _21766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17862_ _17862_/A VGND VGND VPWR VPWR _17862_/X sky130_fd_sc_hd__buf_2
XFILLER_117_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19601_ _19630_/A VGND VGND VPWR VPWR _19603_/A sky130_fd_sc_hd__buf_2
X_16813_ _16812_/X VGND VGND VPWR VPWR _16814_/B sky130_fd_sc_hd__inv_2
XFILLER_93_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17793_ _18082_/A VGND VGND VPWR VPWR _17794_/A sky130_fd_sc_hd__buf_2
X_19532_ _19493_/X _19529_/X _17028_/A _19531_/X VGND VGND VPWR VPWR _24188_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15306__A _13925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11834__A _11834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16744_ _16629_/X _16744_/B VGND VGND VPWR VPWR _16744_/X sky130_fd_sc_hd__or2_4
X_13956_ _13956_/A _13956_/B _13956_/C VGND VGND VPWR VPWR _13957_/B sky130_fd_sc_hd__or3_4
XFILLER_59_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14210__A _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22192__B2 _22190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12907_ _12876_/A _12903_/X _12907_/C VGND VGND VPWR VPWR _12907_/X sky130_fd_sc_hd__or3_4
X_19463_ _19458_/X _19461_/X HRDATA[12] _19462_/X VGND VGND VPWR VPWR _19742_/A sky130_fd_sc_hd__o22a_4
X_13887_ _13887_/A _13807_/B VGND VGND VPWR VPWR _13887_/X sky130_fd_sc_hd__or2_4
X_16675_ _16622_/A _16675_/B _16674_/X VGND VGND VPWR VPWR _16675_/X sky130_fd_sc_hd__or3_4
X_18414_ _16975_/B VGND VGND VPWR VPWR _18414_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12838_ _12771_/X _12838_/B _12837_/X VGND VGND VPWR VPWR _12839_/C sky130_fd_sc_hd__or3_4
X_15626_ _15626_/A _15624_/X _15625_/X VGND VGND VPWR VPWR _15627_/C sky130_fd_sc_hd__and3_4
X_19394_ _19392_/X _18417_/Y _19392_/X _24205_/Q VGND VGND VPWR VPWR _19394_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22139__A _20915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18747__A1_N _17007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18345_ _16972_/A VGND VGND VPWR VPWR _18349_/A sky130_fd_sc_hd__buf_2
XFILLER_37_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ _12769_/A _12769_/B _12769_/C VGND VGND VPWR VPWR _12769_/X sky130_fd_sc_hd__and3_4
X_15557_ _15571_/A _15555_/X _15557_/C VGND VGND VPWR VPWR _15557_/X sky130_fd_sc_hd__and3_4
XANTENNA__22495__A2 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16137__A _16113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508_ _13890_/A VGND VGND VPWR VPWR _14554_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_2_1_0_HCLK_A clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21978__A _21970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15488_ _13765_/A _15486_/X _15487_/X VGND VGND VPWR VPWR _15488_/X sky130_fd_sc_hd__and3_4
X_18276_ _17512_/A _18275_/X VGND VGND VPWR VPWR _18276_/X sky130_fd_sc_hd__or2_4
XFILLER_15_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17227_ _17227_/A VGND VGND VPWR VPWR _17824_/A sky130_fd_sc_hd__buf_2
X_14439_ _12441_/A _14505_/B VGND VGND VPWR VPWR _14441_/B sky130_fd_sc_hd__or2_4
XANTENNA__22247__A2 _22243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17894__C _16999_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17158_ _13920_/X _17155_/X _17156_/Y _17157_/X VGND VGND VPWR VPWR _17158_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17123__A1 _15120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17123__B2 _17122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24358__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16109_ _16109_/A _16109_/B _16108_/X VGND VGND VPWR VPWR _16113_/B sky130_fd_sc_hd__and3_4
XANTENNA__13496__A _15876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17089_ _17088_/X VGND VGND VPWR VPWR _18101_/A sky130_fd_sc_hd__buf_2
XANTENNA__21758__A1 _21536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_14_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21758__B2 _21752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16600__A _11692_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21218__A _21230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22810_ _22807_/A _14786_/Y VGND VGND VPWR VPWR _22810_/X sky130_fd_sc_hd__or2_4
XFILLER_61_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11744__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15216__A _14243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23790_ _23342_/CLK _23790_/D VGND VGND VPWR VPWR _15763_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22741_ _22741_/A VGND VGND VPWR VPWR _22741_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_1_HCLK clkbuf_1_0_1_HCLK/A VGND VGND VPWR VPWR clkbuf_2_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21930__B2 _21928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19337__A2_N _18410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17431__A _15646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22672_ _22686_/A VGND VGND VPWR VPWR _22672_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22049__A _22035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24411_ _24277_/CLK _18825_/X HRESETn VGND VGND VPWR VPWR _24411_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23214__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21623_ _21602_/A VGND VGND VPWR VPWR _21623_/X sky130_fd_sc_hd__buf_2
XANTENNA__24156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12575__A _12575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24342_ _24334_/CLK _24342_/D HRESETn VGND VGND VPWR VPWR _11527_/A sky130_fd_sc_hd__dfstp_4
X_21554_ _21553_/X _21544_/X _23754_/Q _21551_/X VGND VGND VPWR VPWR _21554_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20792__A _20792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20505_ _20444_/X _20491_/Y _20503_/X _20504_/Y _20459_/X VGND VGND VPWR VPWR _20505_/X
+ sky130_fd_sc_hd__a32o_4
X_24273_ _23326_/CLK _24273_/D HRESETn VGND VGND VPWR VPWR _24273_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22238__A2 _22236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21485_ _21270_/X _21484_/X _23785_/Q _21481_/X VGND VGND VPWR VPWR _21485_/X sky130_fd_sc_hd__o22a_4
X_23224_ _23313_/CLK _22480_/X VGND VGND VPWR VPWR _15992_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13923__A1 _13837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21446__B1 _23807_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20436_ _20436_/A VGND VGND VPWR VPWR _20436_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21997__B2 _21992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23155_ _23155_/CLK _22587_/X VGND VGND VPWR VPWR _12945_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18862__A1 _15121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20367_ _18000_/X _20238_/X _20319_/X _20366_/Y VGND VGND VPWR VPWR _20367_/X sky130_fd_sc_hd__a211o_4
XFILLER_84_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18862__B2 _18835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22106_ _22105_/X _22101_/X _13166_/B _22096_/X VGND VGND VPWR VPWR _23441_/D sky130_fd_sc_hd__o22a_4
X_23086_ _23564_/CLK _22694_/X VGND VGND VPWR VPWR _15762_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20298_ _20297_/Y _20258_/X VGND VGND VPWR VPWR _20298_/X sky130_fd_sc_hd__or2_4
XFILLER_103_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21749__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22037_ _21814_/X _22031_/X _12735_/B _22035_/X VGND VGND VPWR VPWR _23476_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11654__A _14073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13810_ _15429_/A _23591_/Q VGND VGND VPWR VPWR _13812_/B sky130_fd_sc_hd__or2_4
XFILLER_29_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15126__A _12209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14790_ _13694_/A _14790_/B VGND VGND VPWR VPWR _14790_/X sky130_fd_sc_hd__or2_4
X_23988_ _24021_/CLK _21132_/X VGND VGND VPWR VPWR _23988_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22174__A1 _22103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22174__B2 _22169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13741_ _11648_/X _13651_/B VGND VGND VPWR VPWR _13741_/X sky130_fd_sc_hd__or2_4
X_22939_ _22962_/A _22939_/B VGND VGND VPWR VPWR _22939_/Y sky130_fd_sc_hd__nand2_4
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_18_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13672_ _12238_/X _13767_/B VGND VGND VPWR VPWR _13673_/C sky130_fd_sc_hd__or2_4
X_16460_ _16465_/A _16391_/B VGND VGND VPWR VPWR _16460_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12623_ _12622_/X _12623_/B VGND VGND VPWR VPWR _12623_/X sky130_fd_sc_hd__or2_4
X_15411_ _15411_/A _15409_/X _15411_/C VGND VGND VPWR VPWR _15412_/C sky130_fd_sc_hd__and3_4
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16391_ _16002_/A _16391_/B VGND VGND VPWR VPWR _16391_/X sky130_fd_sc_hd__or2_4
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19878__B1 _16919_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12485__A _13659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22477__A2 _22472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15342_ _14000_/A _15269_/B VGND VGND VPWR VPWR _15342_/X sky130_fd_sc_hd__or2_4
X_18130_ _16983_/X VGND VGND VPWR VPWR _18132_/C sky130_fd_sc_hd__inv_2
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ _13046_/A _12661_/B VGND VGND VPWR VPWR _12554_/X sky130_fd_sc_hd__or2_4
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _11505_/A _11504_/Y VGND VGND VPWR VPWR _11506_/A sky130_fd_sc_hd__and2_4
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15273_ _15019_/A _15273_/B VGND VGND VPWR VPWR _15273_/X sky130_fd_sc_hd__or2_4
X_18061_ _18060_/X VGND VGND VPWR VPWR _18061_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15796__A _15823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12485_ _13659_/A VGND VGND VPWR VPWR _13622_/A sky130_fd_sc_hd__buf_2
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14224_ _14020_/A VGND VGND VPWR VPWR _14243_/A sky130_fd_sc_hd__buf_2
X_17012_ _17012_/A VGND VGND VPWR VPWR _17013_/A sky130_fd_sc_hd__buf_2
XFILLER_32_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14155_ _14603_/A VGND VGND VPWR VPWR _14737_/A sky130_fd_sc_hd__buf_2
XANTENNA__18853__A1 _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13106_ _13128_/A _13106_/B _13106_/C VGND VGND VPWR VPWR _13110_/B sky130_fd_sc_hd__and3_4
XANTENNA__20660__A1 _20468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14086_ _13972_/A _14086_/B _14085_/X VGND VGND VPWR VPWR _14086_/X sky130_fd_sc_hd__or3_4
X_18963_ _18956_/X _18962_/X _18956_/X _11530_/A VGND VGND VPWR VPWR _24345_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20660__B2 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22422__A _20590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13037_ _12917_/A _13035_/X _13036_/X VGND VGND VPWR VPWR _13041_/B sky130_fd_sc_hd__and3_4
X_17914_ _17811_/A VGND VGND VPWR VPWR _17914_/X sky130_fd_sc_hd__buf_2
XFILLER_65_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17516__A _13575_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18894_ _12990_/X _18891_/X _24371_/Q _18892_/X VGND VGND VPWR VPWR _24371_/D sky130_fd_sc_hd__o22a_4
XFILLER_26_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17845_ _17845_/A VGND VGND VPWR VPWR _17845_/X sky130_fd_sc_hd__buf_2
XFILLER_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15036__A _15036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17776_ _18203_/A VGND VGND VPWR VPWR _18062_/A sky130_fd_sc_hd__buf_2
X_14988_ _14988_/A VGND VGND VPWR VPWR _14988_/X sky130_fd_sc_hd__buf_2
X_19515_ _19630_/A _19481_/B VGND VGND VPWR VPWR _19516_/A sky130_fd_sc_hd__or2_4
X_16727_ _12086_/A _23483_/Q VGND VGND VPWR VPWR _16729_/B sky130_fd_sc_hd__or2_4
X_13939_ _12472_/X _13939_/B VGND VGND VPWR VPWR _13940_/C sky130_fd_sc_hd__or2_4
XANTENNA__21912__B2 _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19446_ _19449_/A VGND VGND VPWR VPWR _19678_/A sky130_fd_sc_hd__buf_2
X_16658_ _16651_/A _16658_/B VGND VGND VPWR VPWR _16659_/C sky130_fd_sc_hd__or2_4
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15609_ _15633_/A _23531_/Q VGND VGND VPWR VPWR _15610_/C sky130_fd_sc_hd__or2_4
Xclkbuf_5_5_0_HCLK clkbuf_4_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19377_ _19302_/X VGND VGND VPWR VPWR _19377_/X sky130_fd_sc_hd__buf_2
X_16589_ _16586_/A _23708_/Q VGND VGND VPWR VPWR _16591_/B sky130_fd_sc_hd__or2_4
XFILLER_72_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12395__A _15743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18328_ _17794_/X _18425_/B _18076_/X _18327_/X VGND VGND VPWR VPWR _18328_/X sky130_fd_sc_hd__a211o_4
XFILLER_37_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21501__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18259_ _18198_/X _18257_/X _18224_/X _18258_/X VGND VGND VPWR VPWR _18259_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18082__A _18082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21428__B1 _23821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21270_ _21555_/A VGND VGND VPWR VPWR _21270_/X sky130_fd_sc_hd__buf_2
XANTENNA__12842__B _12841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21979__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16314__B _16248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20221_ _20223_/A _20216_/X _20217_/X _20218_/X _20220_/X VGND VGND VPWR VPWR _20618_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11739__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18844__A1 _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14115__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20152_ _20141_/Y _20142_/Y _11556_/X _20151_/X VGND VGND VPWR VPWR _20152_/X sky130_fd_sc_hd__o22a_4
X_20083_ _11625_/X _18626_/X VGND VGND VPWR VPWR _20083_/X sky130_fd_sc_hd__or2_4
XFILLER_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16330__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23911_ _23816_/CLK _21276_/X VGND VGND VPWR VPWR _23911_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20954__A2 _20945_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23842_ _23812_/CLK _21393_/X VGND VGND VPWR VPWR _15307_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22156__B2 _22155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12289__B _12289_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24162__CLK _24162_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23773_ _23707_/CLK _21509_/X VGND VGND VPWR VPWR _23773_/Q sky130_fd_sc_hd__dfxtp_4
X_20985_ _20875_/A _20800_/A VGND VGND VPWR VPWR _20985_/X sky130_fd_sc_hd__or2_4
XFILLER_81_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21903__A1 _21843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21903__B2 _21898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22724_ _19497_/X _22723_/Y HREADY VGND VGND VPWR VPWR _22724_/X sky130_fd_sc_hd__o21a_4
XFILLER_92_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18375__A3 _18371_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22655_ _22446_/X _22650_/X _14308_/B _22654_/X VGND VGND VPWR VPWR _23110_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22459__A2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21606_ _21531_/X _21605_/X _12929_/B _21602_/X VGND VGND VPWR VPWR _21606_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21667__B1 _23691_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22586_ _22586_/A VGND VGND VPWR VPWR _22586_/X sky130_fd_sc_hd__buf_2
XANTENNA__22507__A _22471_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24325_ _24330_/CLK _24325_/D HRESETn VGND VGND VPWR VPWR _24325_/Q sky130_fd_sc_hd__dfstp_4
X_21537_ _21536_/X _21532_/X _13145_/B _21527_/X VGND VGND VPWR VPWR _23761_/D sky130_fd_sc_hd__o22a_4
X_12270_ _12235_/A _12270_/B VGND VGND VPWR VPWR _12270_/X sky130_fd_sc_hd__or2_4
X_24256_ _24321_/CLK _24256_/D HRESETn VGND VGND VPWR VPWR _19205_/A sky130_fd_sc_hd__dfrtp_4
X_21468_ _21241_/X _21463_/X _12658_/B _21467_/X VGND VGND VPWR VPWR _21468_/X sky130_fd_sc_hd__o22a_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23207_ _23847_/CLK _23207_/D VGND VGND VPWR VPWR _13824_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_5_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20419_ _21804_/A VGND VGND VPWR VPWR _20419_/X sky130_fd_sc_hd__buf_2
XANTENNA__11649__A _11648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22092__B1 _16189_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24187_ _24187_/CLK _19548_/Y HRESETn VGND VGND VPWR VPWR _17262_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22631__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21399_ _21398_/X VGND VGND VPWR VPWR _21400_/A sky130_fd_sc_hd__buf_2
XANTENNA__14025__A _11647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23138_ _24065_/CLK _23138_/D VGND VGND VPWR VPWR _15276_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24341__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15960_ _16096_/A _15960_/B VGND VGND VPWR VPWR _15960_/X sky130_fd_sc_hd__or2_4
X_23069_ _16893_/A VGND VGND VPWR VPWR HSIZE[0] sky130_fd_sc_hd__buf_2
XANTENNA__23057__B _23038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16240__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21198__A2 _21197_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22395__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14911_ _15015_/A _14909_/X _14911_/C VGND VGND VPWR VPWR _14911_/X sky130_fd_sc_hd__and3_4
X_15891_ _15879_/A _15835_/B VGND VGND VPWR VPWR _15893_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_60_0_HCLK clkbuf_6_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17630_ _17278_/X _17629_/Y _17902_/B VGND VGND VPWR VPWR _17630_/X sky130_fd_sc_hd__o21a_4
X_14842_ _14811_/A _14770_/B VGND VGND VPWR VPWR _14842_/X sky130_fd_sc_hd__or2_4
XANTENNA__17810__A2 _17805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17561_ _11598_/X _17561_/B VGND VGND VPWR VPWR _17561_/X sky130_fd_sc_hd__and2_4
X_11985_ _11916_/X _11985_/B _11985_/C VGND VGND VPWR VPWR _11989_/B sky130_fd_sc_hd__and3_4
X_14773_ _13645_/A _14773_/B VGND VGND VPWR VPWR _14774_/C sky130_fd_sc_hd__or2_4
XFILLER_17_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22698__A2 _22693_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14695__A _14679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19300_ _23064_/B _24255_/Q _19299_/Y VGND VGND VPWR VPWR _24255_/D sky130_fd_sc_hd__o21a_4
X_16512_ _16231_/A _16496_/X _16512_/C VGND VGND VPWR VPWR _16513_/C sky130_fd_sc_hd__or3_4
X_13724_ _15494_/A _23560_/Q VGND VGND VPWR VPWR _13725_/C sky130_fd_sc_hd__or2_4
XFILLER_32_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17492_ _17194_/X _17517_/B VGND VGND VPWR VPWR _17492_/X sky130_fd_sc_hd__or2_4
XFILLER_44_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21370__A2 _21369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19231_ _19231_/A _19245_/A VGND VGND VPWR VPWR _19231_/X sky130_fd_sc_hd__and2_4
X_16443_ _11843_/X _11618_/X _16412_/X _11597_/X _16442_/X VGND VGND VPWR VPWR _16443_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_32_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13655_ _13794_/A _23592_/Q VGND VGND VPWR VPWR _13655_/X sky130_fd_sc_hd__or2_4
XFILLER_73_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13104__A _13104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12606_ _12652_/A VGND VGND VPWR VPWR _12643_/A sky130_fd_sc_hd__buf_2
X_19162_ _19128_/A _19163_/A _19161_/Y VGND VGND VPWR VPWR _24307_/D sky130_fd_sc_hd__o21a_4
X_13586_ _13586_/A _13585_/Y VGND VGND VPWR VPWR _13586_/Y sky130_fd_sc_hd__nor2_4
X_16374_ _16374_/A VGND VGND VPWR VPWR _16374_/X sky130_fd_sc_hd__buf_2
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18113_ _17975_/A _18111_/X _17797_/X _18112_/X VGND VGND VPWR VPWR _18113_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12537_ _12466_/X _12535_/X _12537_/C VGND VGND VPWR VPWR _12541_/B sky130_fd_sc_hd__and3_4
X_15325_ _14177_/A VGND VGND VPWR VPWR _15325_/X sky130_fd_sc_hd__buf_2
X_19093_ _19092_/Y _11506_/A _11508_/B VGND VGND VPWR VPWR _19093_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16415__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18044_ _17103_/X _18039_/Y _17240_/X _18043_/X VGND VGND VPWR VPWR _18044_/X sky130_fd_sc_hd__a211o_4
X_12468_ _13019_/A VGND VGND VPWR VPWR _12518_/A sky130_fd_sc_hd__buf_2
X_15256_ _14575_/X _15256_/B VGND VGND VPWR VPWR _15256_/X sky130_fd_sc_hd__or2_4
XANTENNA__16134__B _16211_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14207_ _14207_/A VGND VGND VPWR VPWR _14371_/A sky130_fd_sc_hd__buf_2
X_15187_ _11709_/A _15126_/B VGND VGND VPWR VPWR _15188_/C sky130_fd_sc_hd__or2_4
XANTENNA__18826__A1 _16514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12399_ _15882_/A _12399_/B _12398_/X VGND VGND VPWR VPWR _12407_/B sky130_fd_sc_hd__or3_4
XFILLER_99_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14138_ _14121_/A VGND VGND VPWR VPWR _14138_/X sky130_fd_sc_hd__buf_2
XFILLER_99_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21830__B1 _15685_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19995_ _19995_/A VGND VGND VPWR VPWR _19995_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13774__A _13685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14069_ _14046_/A _14069_/B _14068_/X VGND VGND VPWR VPWR _14069_/X sky130_fd_sc_hd__and3_4
X_18946_ _18999_/A VGND VGND VPWR VPWR _18946_/X sky130_fd_sc_hd__buf_2
XFILLER_113_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21189__A2 _21183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24185__CLK _24162_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18877_ _18877_/A VGND VGND VPWR VPWR _18892_/A sky130_fd_sc_hd__buf_2
XFILLER_95_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17828_ _17814_/X _17183_/X _17804_/X _17174_/X VGND VGND VPWR VPWR _17828_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22138__B2 _22132_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17759_ _17680_/A _17479_/X _17680_/X VGND VGND VPWR VPWR _17759_/X sky130_fd_sc_hd__a21bo_4
XANTENNA__22689__A2 _22686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20400__A _20342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21897__B1 _15471_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20770_ _20759_/X _20768_/X _24297_/Q _20769_/X VGND VGND VPWR VPWR _20771_/B sky130_fd_sc_hd__o22a_4
XFILLER_74_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16309__B _16244_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19429_ _19429_/A VGND VGND VPWR VPWR _19485_/A sky130_fd_sc_hd__inv_2
XFILLER_90_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15213__B _15213_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13014__A _13014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22440_ _22384_/X VGND VGND VPWR VPWR _22440_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21649__B1 _23704_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22371_ _22129_/X _22368_/X _13863_/B _22365_/X VGND VGND VPWR VPWR _22371_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12853__A _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24110_ _24202_/CLK _24110_/D HRESETn VGND VGND VPWR VPWR _16996_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21322_ _21251_/X _21319_/X _13171_/B _21316_/X VGND VGND VPWR VPWR _23889_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_2_0_0_HCLK clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_2_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24041_ _23910_/CLK _24041_/D VGND VGND VPWR VPWR _24041_/Q sky130_fd_sc_hd__dfxtp_4
X_21253_ _20591_/A VGND VGND VPWR VPWR _21253_/X sky130_fd_sc_hd__buf_2
XANTENNA__22613__A2 _22586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20204_ _16929_/X VGND VGND VPWR VPWR _20399_/A sky130_fd_sc_hd__buf_2
XFILLER_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20624__B2 _20449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21184_ _20537_/X _21183_/X _23955_/Q _21180_/X VGND VGND VPWR VPWR _23955_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15883__B _15821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20135_ _24432_/Q VGND VGND VPWR VPWR _20135_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17156__A _12430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16060__A _16215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22997__A _22967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14854__A2 _14851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22377__B2 _22372_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20066_ _24455_/Q VGND VGND VPWR VPWR _20066_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_4_0_HCLK_A clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23825_ _23889_/CLK _23825_/D VGND VGND VPWR VPWR _13179_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_113_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15404__A _15404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11932__A _13048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24100__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11770_ _12822_/A VGND VGND VPWR VPWR _11770_/X sky130_fd_sc_hd__buf_2
X_23756_ _23404_/CLK _23756_/D VGND VGND VPWR VPWR _15463_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20968_ _20968_/A VGND VGND VPWR VPWR _20968_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18753__B1 _17737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16219__B _16219_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22707_ _22671_/A VGND VGND VPWR VPWR _22707_/X sky130_fd_sc_hd__buf_2
XANTENNA__11651__B _13991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23687_ _23336_/CLK _21672_/X VGND VGND VPWR VPWR _13831_/B sky130_fd_sc_hd__dfxtp_4
X_20899_ _20214_/Y _20897_/X _20898_/X VGND VGND VPWR VPWR _20899_/X sky130_fd_sc_hd__a21o_4
XFILLER_41_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13440_ _13467_/A _13440_/B _13440_/C VGND VGND VPWR VPWR _13441_/C sky130_fd_sc_hd__and3_4
XFILLER_70_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22638_ _22418_/X _22636_/X _13111_/B _22633_/X VGND VGND VPWR VPWR _22638_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22882__D _19894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21104__A2 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14962__B _14962_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13371_ _12787_/A _13363_/X _13371_/C VGND VGND VPWR VPWR _13391_/B sky130_fd_sc_hd__and3_4
X_22569_ _22576_/A VGND VGND VPWR VPWR _22569_/X sky130_fd_sc_hd__buf_2
XFILLER_107_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12763__A _12754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12322_ _15706_/A VGND VGND VPWR VPWR _12738_/A sky130_fd_sc_hd__buf_2
X_15110_ _15110_/A _24063_/Q VGND VGND VPWR VPWR _15110_/X sky130_fd_sc_hd__or2_4
XANTENNA__20863__A1 _18624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16090_ _16090_/A VGND VGND VPWR VPWR _16091_/A sky130_fd_sc_hd__buf_2
X_24308_ _24301_/CLK _24308_/D HRESETn VGND VGND VPWR VPWR _19129_/A sky130_fd_sc_hd__dfrtp_4
X_15041_ _15041_/A _23775_/Q VGND VGND VPWR VPWR _15042_/C sky130_fd_sc_hd__or2_4
X_12253_ _15448_/A VGND VGND VPWR VPWR _13670_/A sky130_fd_sc_hd__buf_2
X_24239_ _24239_/CLK _24239_/D HRESETn VGND VGND VPWR VPWR _24239_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18808__A1 _15249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22065__B1 _15033_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12184_ _12184_/A VGND VGND VPWR VPWR _12184_/X sky130_fd_sc_hd__buf_2
XANTENNA__23082__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18800_ _13918_/X _18795_/X _24423_/Q _18796_/X VGND VGND VPWR VPWR _18800_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13594__A _11841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19780_ _19667_/A _19779_/X VGND VGND VPWR VPWR _19780_/X sky130_fd_sc_hd__and2_4
X_16992_ _16992_/A VGND VGND VPWR VPWR _16992_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18731_ _17926_/X _18730_/Y _17812_/X _17973_/Y VGND VGND VPWR VPWR _18731_/X sky130_fd_sc_hd__o22a_4
X_15943_ _11933_/X VGND VGND VPWR VPWR _15980_/A sky130_fd_sc_hd__buf_2
XFILLER_95_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22700__A _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18662_ _18662_/A _18662_/B VGND VGND VPWR VPWR _18662_/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21040__B2 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15874_ _13557_/A _15866_/X _15874_/C VGND VGND VPWR VPWR _15875_/C sky130_fd_sc_hd__and3_4
X_17613_ _17612_/X VGND VGND VPWR VPWR _17613_/Y sky130_fd_sc_hd__inv_2
X_14825_ _13706_/A _14821_/X _14824_/X VGND VGND VPWR VPWR _14833_/B sky130_fd_sc_hd__or3_4
XFILLER_97_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21316__A _21316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18593_ _17878_/X _18585_/Y _18586_/X _17998_/X _18592_/X VGND VGND VPWR VPWR _18593_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11842__A _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17544_ _17039_/A _17543_/X _17043_/A VGND VGND VPWR VPWR _17544_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21879__B1 _23577_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14756_ _14756_/A _14820_/B VGND VGND VPWR VPWR _14756_/X sky130_fd_sc_hd__or2_4
X_11968_ _12022_/A VGND VGND VPWR VPWR _12008_/A sky130_fd_sc_hd__buf_2
XANTENNA__21343__A2 _21340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13707_ _13893_/A VGND VGND VPWR VPWR _13747_/A sky130_fd_sc_hd__buf_2
XANTENNA__19736__A2_N _19734_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15033__B _15033_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17475_ _18152_/A VGND VGND VPWR VPWR _18191_/A sky130_fd_sc_hd__inv_2
X_11899_ _13463_/A VGND VGND VPWR VPWR _15956_/A sky130_fd_sc_hd__buf_2
X_14687_ _13886_/A _14670_/X _14686_/X VGND VGND VPWR VPWR _14719_/B sky130_fd_sc_hd__or3_4
XANTENNA__20551__B1 _20550_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_67_0_HCLK clkbuf_7_66_0_HCLK/A VGND VGND VPWR VPWR _24301_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20874__B _20490_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19214_ _24265_/Q _19214_/B VGND VGND VPWR VPWR _19215_/B sky130_fd_sc_hd__and2_4
XFILLER_34_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16426_ _15929_/X _16422_/X _16426_/C VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__or3_4
X_13638_ _15412_/A _13638_/B _13638_/C VGND VGND VPWR VPWR _13638_/X sky130_fd_sc_hd__or3_4
XANTENNA__22147__A _21001_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21051__A _21015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19145_ _19136_/X VGND VGND VPWR VPWR _19145_/Y sky130_fd_sc_hd__inv_2
X_16357_ _16323_/A _16294_/B VGND VGND VPWR VPWR _16358_/C sky130_fd_sc_hd__or2_4
XFILLER_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13569_ _13562_/A _13569_/B VGND VGND VPWR VPWR _13570_/C sky130_fd_sc_hd__or2_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16145__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12673__A _12989_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15308_ _14748_/A _15308_/B _15307_/X VGND VGND VPWR VPWR _15308_/X sky130_fd_sc_hd__and3_4
X_19076_ _24325_/Q VGND VGND VPWR VPWR _19076_/Y sky130_fd_sc_hd__inv_2
X_16288_ _15976_/A _16286_/X _16287_/X VGND VGND VPWR VPWR _16292_/B sky130_fd_sc_hd__and3_4
X_18027_ _18241_/A _17549_/B VGND VGND VPWR VPWR _18027_/Y sky130_fd_sc_hd__nor2_4
XFILLER_103_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15239_ _14190_/A _15235_/X _15238_/X VGND VGND VPWR VPWR _15247_/B sky130_fd_sc_hd__or3_4
XFILLER_99_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18360__A _18242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20606__A1 _20212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16799__B _23707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19978_ _18006_/X _19961_/X _19977_/Y _19972_/X VGND VGND VPWR VPWR _19978_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23575__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22359__B2 _22358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18929_ _24382_/Q _20268_/A _18927_/X _24350_/Q _18928_/Y VGND VGND VPWR VPWR _18929_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_45_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15208__B _23649_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_HCLK HCLK VGND VGND VPWR VPWR clkbuf_0_HCLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_41_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21031__A1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21940_ _21819_/X _21938_/X _23538_/Q _21935_/X VGND VGND VPWR VPWR _21940_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13009__A _13009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21031__B2 _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21871_ _21865_/Y _21870_/X _21789_/X _21870_/X VGND VGND VPWR VPWR _21871_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20130__A _19313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12848__A _12444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23610_ _23699_/CLK _23610_/D VGND VGND VPWR VPWR _23610_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19527__A2 _19829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20822_ _20445_/B _20822_/B VGND VGND VPWR VPWR _20823_/C sky130_fd_sc_hd__or2_4
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21334__A2 _21333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23541_ _23315_/CLK _23541_/D VGND VGND VPWR VPWR _12633_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20753_ HRDATA[10] _20753_/B VGND VGND VPWR VPWR _20753_/X sky130_fd_sc_hd__or2_4
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23472_ _23472_/CLK _22043_/X VGND VGND VPWR VPWR _23472_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20684_ _20681_/X _20683_/X _24364_/Q _20625_/X VGND VGND VPWR VPWR _20684_/X sky130_fd_sc_hd__o22a_4
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22423_ _22423_/A VGND VGND VPWR VPWR _22423_/X sky130_fd_sc_hd__buf_2
XFILLER_52_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21098__A1 _20797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21098__B2 _21093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22354_ _22354_/A VGND VGND VPWR VPWR _22354_/X sky130_fd_sc_hd__buf_2
XFILLER_108_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21305_ _21319_/A VGND VGND VPWR VPWR _21305_/X sky130_fd_sc_hd__buf_2
XANTENNA__22047__B1 _15828_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15894__A _13551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22285_ _22122_/X _22279_/X _23338_/Q _22283_/X VGND VGND VPWR VPWR _22285_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24024_ _23316_/CLK _21076_/X VGND VGND VPWR VPWR _24024_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23918__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22598__B2 _22597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21236_ _21234_/X _21235_/X _23928_/Q _21230_/X VGND VGND VPWR VPWR _23928_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21167_ _21161_/Y _21166_/X _20277_/X _21166_/X VGND VGND VPWR VPWR _21167_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14303__A _12307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20118_ _11544_/X VGND VGND VPWR VPWR _20118_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21098_ _20797_/X _21096_/X _24008_/Q _21093_/X VGND VGND VPWR VPWR _21098_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21022__B2 _21020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12940_ _12964_/A _12934_/X _12940_/C VGND VGND VPWR VPWR _12941_/C sky130_fd_sc_hd__or3_4
X_20049_ _24459_/Q VGND VGND VPWR VPWR _20049_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21573__A2 _21568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12871_ _12920_/A VGND VGND VPWR VPWR _12910_/A sky130_fd_sc_hd__buf_2
XANTENNA__22717__A1_N _19674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ _14725_/A _14691_/B VGND VGND VPWR VPWR _14610_/X sky130_fd_sc_hd__or2_4
XANTENNA__11662__A _14039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11822_ _11780_/X _23870_/Q VGND VGND VPWR VPWR _11822_/X sky130_fd_sc_hd__or2_4
X_23808_ _23840_/CLK _23808_/D VGND VGND VPWR VPWR _23808_/Q sky130_fd_sc_hd__dfxtp_4
X_15590_ _15614_/A _23179_/Q VGND VGND VPWR VPWR _15590_/X sky130_fd_sc_hd__or2_4
XANTENNA__17529__A1 _17156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21325__A2 _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _16023_/A VGND VGND VPWR VPWR _16064_/A sky130_fd_sc_hd__buf_2
X_14541_ _14494_/X _14541_/B _14540_/X VGND VGND VPWR VPWR _14541_/X sky130_fd_sc_hd__and3_4
X_23739_ _23707_/CLK _23739_/D VGND VGND VPWR VPWR _23739_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20533__B1 _20532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14973__A _15072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17103_/X _18716_/B _17240_/X _17259_/X VGND VGND VPWR VPWR _17260_/X sky130_fd_sc_hd__a211o_4
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _16198_/A VGND VGND VPWR VPWR _11684_/X sky130_fd_sc_hd__buf_2
X_14472_ _13019_/A _14472_/B VGND VGND VPWR VPWR _14474_/B sky130_fd_sc_hd__or2_4
XFILLER_14_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _16219_/A _16211_/B VGND VGND VPWR VPWR _16211_/X sky130_fd_sc_hd__or2_4
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _12787_/A _13423_/B _13423_/C VGND VGND VPWR VPWR _13423_/X sky130_fd_sc_hd__and3_4
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17191_ _15517_/X VGND VGND VPWR VPWR _17191_/X sky130_fd_sc_hd__buf_2
XANTENNA__12493__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13354_ _12803_/A VGND VGND VPWR VPWR _13354_/X sky130_fd_sc_hd__buf_2
X_16142_ _16139_/A _23639_/Q VGND VGND VPWR VPWR _16143_/C sky130_fd_sc_hd__or2_4
XFILLER_10_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17701__B2 _17354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12305_ _12713_/A VGND VGND VPWR VPWR _13317_/A sky130_fd_sc_hd__buf_2
XFILLER_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13285_ _13281_/X _13282_/X _13284_/X VGND VGND VPWR VPWR _13285_/X sky130_fd_sc_hd__and3_4
X_16073_ _16063_/A _16071_/X _16072_/X VGND VGND VPWR VPWR _16073_/X sky130_fd_sc_hd__and3_4
XFILLER_115_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22589__B2 _22583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12236_ _12693_/A _12236_/B VGND VGND VPWR VPWR _12236_/X sky130_fd_sc_hd__or2_4
X_15024_ _15028_/A _15024_/B _15024_/C VGND VGND VPWR VPWR _15024_/X sky130_fd_sc_hd__and3_4
X_19901_ _22968_/A VGND VGND VPWR VPWR _19901_/X sky130_fd_sc_hd__buf_2
XFILLER_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_HCLK clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19832_ _19449_/X _19828_/X _19829_/X _21348_/B _19531_/A VGND VGND VPWR VPWR _19832_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11837__A _16077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12167_ _12167_/A _23101_/Q VGND VGND VPWR VPWR _12169_/B sky130_fd_sc_hd__or2_4
XANTENNA__15309__A _14782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19763_ _20576_/B _19496_/X _19762_/X _19616_/X VGND VGND VPWR VPWR _19763_/X sky130_fd_sc_hd__a211o_4
XANTENNA__11556__B IRQ[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12098_ _12098_/A _24093_/Q VGND VGND VPWR VPWR _12099_/C sky130_fd_sc_hd__or2_4
X_16975_ _17699_/A _16975_/B VGND VGND VPWR VPWR _16976_/B sky130_fd_sc_hd__or2_4
XFILLER_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22430__A _20670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18714_ _18714_/A _17330_/A VGND VGND VPWR VPWR _18714_/X sky130_fd_sc_hd__and2_4
XFILLER_77_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17217__B1 _15251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19757__A2 _19789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15926_ _13280_/X _13593_/X _16899_/A _15926_/D VGND VGND VPWR VPWR _15926_/X sky130_fd_sc_hd__or4_4
XANTENNA__17524__A _12990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19694_ _19625_/Y _19687_/X _19663_/A _19692_/X _19693_/X VGND VGND VPWR VPWR _19694_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_20_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21564__A2 _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_30_0_HCLK clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18645_ _18643_/X _18644_/X _18643_/X _18644_/X VGND VGND VPWR VPWR _18645_/X sky130_fd_sc_hd__a2bb2o_4
X_15857_ _13529_/X _15855_/X _15856_/X VGND VGND VPWR VPWR _15858_/C sky130_fd_sc_hd__and3_4
XFILLER_25_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12668__A _12622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14808_ _13706_/A _14804_/X _14807_/X VGND VGND VPWR VPWR _14817_/B sky130_fd_sc_hd__or3_4
XFILLER_24_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24223__CLK _24223_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18576_ _17745_/A _18575_/X _17745_/A _18575_/X VGND VGND VPWR VPWR _18576_/X sky130_fd_sc_hd__a2bb2o_4
X_15788_ _15785_/A _15849_/B VGND VGND VPWR VPWR _15789_/C sky130_fd_sc_hd__or2_4
XFILLER_17_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18717__B1 _18249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12387__B _12263_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22513__B2 _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17527_ _12674_/X _17527_/B VGND VGND VPWR VPWR _17527_/Y sky130_fd_sc_hd__nand2_4
X_14739_ _13606_/A _14739_/B VGND VGND VPWR VPWR _14741_/B sky130_fd_sc_hd__or2_4
XFILLER_90_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17458_ _17039_/A _17457_/X _17043_/A VGND VGND VPWR VPWR _17688_/B sky130_fd_sc_hd__o21a_4
XFILLER_20_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16743__A2 _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16409_ _13442_/X _16409_/B _16409_/C VGND VGND VPWR VPWR _16409_/X sky130_fd_sc_hd__and3_4
XANTENNA__14754__A1 _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13499__A _13550_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22277__B1 _13287_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17389_ _13918_/X _17424_/B VGND VGND VPWR VPWR _17390_/B sky130_fd_sc_hd__or2_4
XFILLER_14_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19128_ _19128_/A _19163_/A VGND VGND VPWR VPWR _19129_/B sky130_fd_sc_hd__and2_4
XFILLER_9_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20827__A1 _20681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20827__B2 _20625_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19693__A1 _19582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22029__B1 _16427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19059_ _19046_/X _19058_/X _19046_/X _24329_/Q VGND VGND VPWR VPWR _24329_/D sky130_fd_sc_hd__a2bb2o_4
X_22070_ _22125_/A VGND VGND VPWR VPWR _22108_/A sky130_fd_sc_hd__inv_2
X_21021_ _20373_/X _21016_/X _16417_/B _21020_/X VGND VGND VPWR VPWR _21021_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11747__A _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21252__B2 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14123__A _14998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22340__A _22354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17434__A _15911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13962__A _13966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19748__A2 HRDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22972_ _22972_/A VGND VGND VPWR VPWR HADDR[15] sky130_fd_sc_hd__inv_2
XFILLER_60_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17759__A1 _17680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13493__A1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21923_ _21919_/A VGND VGND VPWR VPWR _21938_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21854_ _21852_/X _21853_/X _14691_/B _21848_/X VGND VGND VPWR VPWR _23588_/D sky130_fd_sc_hd__o22a_4
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21307__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20805_ _20805_/A _20708_/B VGND VGND VPWR VPWR _20805_/X sky130_fd_sc_hd__or2_4
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15889__A _15889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21785_ _21784_/X VGND VGND VPWR VPWR _21792_/A sky130_fd_sc_hd__buf_2
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18265__A _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19381__B1 _19380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20736_ _20497_/A VGND VGND VPWR VPWR _20736_/X sky130_fd_sc_hd__buf_2
X_23524_ _23107_/CLK _23524_/D VGND VGND VPWR VPWR _14683_/B sky130_fd_sc_hd__dfxtp_4
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_50_0_HCLK clkbuf_7_50_0_HCLK/A VGND VGND VPWR VPWR _23688_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23455_ _23487_/CLK _23455_/D VGND VGND VPWR VPWR _15033_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20667_ _24237_/Q _20639_/X _20666_/X VGND VGND VPWR VPWR _20667_/X sky130_fd_sc_hd__o21a_4
XFILLER_104_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22406_ _20441_/A VGND VGND VPWR VPWR _22406_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23386_ _23354_/CLK _22213_/X VGND VGND VPWR VPWR _16423_/B sky130_fd_sc_hd__dfxtp_4
X_20598_ _20425_/X _20595_/Y _20597_/X _19021_/Y _20473_/X VGND VGND VPWR VPWR _20598_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_100_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22337_ _22344_/A VGND VGND VPWR VPWR _22337_/X sky130_fd_sc_hd__buf_2
XANTENNA__16513__A _11658_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13070_ _13112_/A _23730_/Q VGND VGND VPWR VPWR _13070_/X sky130_fd_sc_hd__or2_4
XFILLER_69_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22268_ _22093_/X _22265_/X _12222_/B _22262_/X VGND VGND VPWR VPWR _23350_/D sky130_fd_sc_hd__o22a_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12021_ _11916_/X VGND VGND VPWR VPWR _12025_/A sky130_fd_sc_hd__buf_2
X_24007_ _24008_/CLK _24007_/D VGND VGND VPWR VPWR _13859_/B sky130_fd_sc_hd__dfxtp_4
X_21219_ _21789_/A VGND VGND VPWR VPWR _21219_/X sky130_fd_sc_hd__buf_2
XANTENNA__11657__A _12989_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19987__A2 _19985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21243__B2 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22199_ _22147_/X _22172_/A _23391_/Q _22162_/A VGND VGND VPWR VPWR _23391_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14033__A _12599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21794__A2 _21793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13872__A _13872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16760_ _16757_/X _16760_/B _16760_/C VGND VGND VPWR VPWR _16761_/C sky130_fd_sc_hd__and3_4
XFILLER_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13972_ _13972_/A _13968_/X _13971_/X VGND VGND VPWR VPWR _13972_/X sky130_fd_sc_hd__or3_4
XFILLER_111_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15711_ _12716_/X _15688_/X _15695_/X _15702_/X _15710_/X VGND VGND VPWR VPWR _15711_/X
+ sky130_fd_sc_hd__a32o_4
X_12923_ _11980_/A _12900_/X _12907_/X _12914_/X _12922_/X VGND VGND VPWR VPWR _12923_/X
+ sky130_fd_sc_hd__a32o_4
X_16691_ _16714_/A _23771_/Q VGND VGND VPWR VPWR _16692_/C sky130_fd_sc_hd__or2_4
XFILLER_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12488__A _13031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18430_ _18418_/X _18423_/Y _18426_/X _18428_/X _18429_/Y VGND VGND VPWR VPWR _18430_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_94_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15642_ _13893_/A _15642_/B _15642_/C VGND VGND VPWR VPWR _15643_/C sky130_fd_sc_hd__or3_4
X_12854_ _12464_/A _12851_/X _12854_/C VGND VGND VPWR VPWR _12855_/C sky130_fd_sc_hd__and3_4
XFILLER_76_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11805_ _11748_/X _11803_/X _11804_/X VGND VGND VPWR VPWR _11805_/X sky130_fd_sc_hd__and3_4
X_18361_ _18297_/A _17484_/A VGND VGND VPWR VPWR _18361_/X sky130_fd_sc_hd__and2_4
XANTENNA__15799__A _12865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15573_ _15576_/A _15573_/B VGND VGND VPWR VPWR _15573_/X sky130_fd_sc_hd__or2_4
X_12785_ _12813_/A _12781_/X _12784_/X VGND VGND VPWR VPWR _12785_/X sky130_fd_sc_hd__and3_4
XFILLER_37_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _14429_/B _17313_/B VGND VGND VPWR VPWR _18587_/B sky130_fd_sc_hd__or2_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14536_/A _14447_/B VGND VGND VPWR VPWR _14524_/X sky130_fd_sc_hd__or2_4
X_11736_ _11685_/X _11719_/X _11735_/X VGND VGND VPWR VPWR _11736_/X sky130_fd_sc_hd__or3_4
X_18292_ _17674_/A _16979_/B _16980_/B VGND VGND VPWR VPWR _22987_/B sky130_fd_sc_hd__a21bo_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16407__B _16407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _17863_/A VGND VGND VPWR VPWR _17837_/A sky130_fd_sc_hd__buf_2
XFILLER_70_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22259__B1 _12123_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _12450_/A _14455_/B _14455_/C VGND VGND VPWR VPWR _14455_/X sky130_fd_sc_hd__and3_4
X_11667_ _11666_/X VGND VGND VPWR VPWR _16045_/A sky130_fd_sc_hd__buf_2
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _13388_/A _13404_/X _13406_/C VGND VGND VPWR VPWR _13407_/C sky130_fd_sc_hd__and3_4
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17174_ _17172_/Y _17173_/X _12992_/X _17145_/X VGND VGND VPWR VPWR _17174_/X sky130_fd_sc_hd__o22a_4
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11598_ _11597_/X VGND VGND VPWR VPWR _11598_/X sky130_fd_sc_hd__buf_2
X_14386_ _15626_/A _14386_/B _14385_/X VGND VGND VPWR VPWR _14387_/C sky130_fd_sc_hd__and3_4
XANTENNA__22425__A _20610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16125_ _16108_/A _23959_/Q VGND VGND VPWR VPWR _16126_/C sky130_fd_sc_hd__or2_4
X_13337_ _13428_/A _13337_/B VGND VGND VPWR VPWR _13338_/C sky130_fd_sc_hd__or2_4
XANTENNA__17519__A _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21482__B2 _21481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_7_0_HCLK_A clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12951__A _12951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20690__C1 _20689_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16056_ _16037_/A _15984_/B VGND VGND VPWR VPWR _16058_/B sky130_fd_sc_hd__or2_4
XANTENNA__24274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19427__A1 HRDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13268_ _12392_/A _13268_/B _13268_/C VGND VGND VPWR VPWR _13268_/X sky130_fd_sc_hd__or3_4
XFILLER_100_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15007_ _15030_/A _23519_/Q VGND VGND VPWR VPWR _15008_/C sky130_fd_sc_hd__or2_4
X_12219_ _13796_/A VGND VGND VPWR VPWR _13054_/A sky130_fd_sc_hd__buf_2
XANTENNA__15039__A _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19978__A2 _19961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22431__B1 _15845_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19734__A HRDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13199_ _13004_/A _13195_/X _13198_/X VGND VGND VPWR VPWR _13200_/B sky130_fd_sc_hd__or3_4
XFILLER_48_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19815_ _19445_/X _19814_/X _19494_/X _19730_/A VGND VGND VPWR VPWR _19815_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15981__B _15981_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13782__A _12450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16958_ _24118_/Q VGND VGND VPWR VPWR _16970_/A sky130_fd_sc_hd__inv_2
X_19746_ _19765_/B _19745_/X _19672_/D VGND VGND VPWR VPWR _19746_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21537__A2 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15909_ _15844_/X _15909_/B VGND VGND VPWR VPWR _15909_/X sky130_fd_sc_hd__or2_4
X_19677_ _19667_/X _19673_/X _19534_/X _19676_/X VGND VGND VPWR VPWR _19677_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23613__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16889_ _16822_/X _16889_/B _16831_/X _16888_/X VGND VGND VPWR VPWR _16890_/B sky130_fd_sc_hd__and4_4
XFILLER_77_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18628_ _18628_/A VGND VGND VPWR VPWR _18628_/Y sky130_fd_sc_hd__inv_2
X_18559_ _18558_/X VGND VGND VPWR VPWR _18559_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22498__B1 _23211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15502__A _15497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21570_ _21855_/A VGND VGND VPWR VPWR _21570_/X sky130_fd_sc_hd__buf_2
XFILLER_36_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16317__B _24025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_37_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_75_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20521_ _20520_/Y _20521_/B VGND VGND VPWR VPWR _20521_/X sky130_fd_sc_hd__or2_4
XFILLER_21_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15221__B _23585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19909__A _19909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14118__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23240_ _23816_/CLK _22443_/X VGND VGND VPWR VPWR _13696_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13022__A _13022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20452_ _20403_/X _20451_/X _24278_/Q _20327_/X VGND VGND VPWR VPWR _20452_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24119__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22335__A _22368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23171_ _23107_/CLK _23171_/D VGND VGND VPWR VPWR _14794_/B sky130_fd_sc_hd__dfxtp_4
X_20383_ _20622_/A _20382_/Y _19230_/A _20301_/X VGND VGND VPWR VPWR _20383_/X sky130_fd_sc_hd__o22a_4
XFILLER_31_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21473__B2 _21467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22122_ _20747_/A VGND VGND VPWR VPWR _22122_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17429__B1 _17422_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22053_ _21840_/X _22052_/X _23465_/Q _22049_/X VGND VGND VPWR VPWR _22053_/X sky130_fd_sc_hd__o22a_4
X_21004_ _24062_/Q VGND VGND VPWR VPWR _21004_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22973__A1 _17893_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15891__B _15835_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22070__A _22125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17164__A _16077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22725__A1 _22898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21528__A2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22725__B2 _19380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22955_ _22985_/A VGND VGND VPWR VPWR _22955_/X sky130_fd_sc_hd__buf_2
XFILLER_56_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21906_ _21847_/X _21901_/X _14293_/B _21905_/X VGND VGND VPWR VPWR _23558_/D sky130_fd_sc_hd__o22a_4
X_22886_ _22985_/A VGND VGND VPWR VPWR _22886_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_119_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR _24021_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21837_ _21835_/X _21829_/X _23595_/Q _21836_/X VGND VGND VPWR VPWR _23595_/D sky130_fd_sc_hd__o22a_4
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16508__A _16159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15412__A _15412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12570_ _15487_/A VGND VGND VPWR VPWR _12959_/A sky130_fd_sc_hd__buf_2
XFILLER_54_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21768_ _21553_/X _21762_/X _23626_/Q _21766_/X VGND VGND VPWR VPWR _23626_/D sky130_fd_sc_hd__o22a_4
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21700__A2 _21698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11521_ _24336_/Q _11521_/B VGND VGND VPWR VPWR _19008_/A sky130_fd_sc_hd__or2_4
X_20719_ _24235_/Q _20639_/X _20718_/X VGND VGND VPWR VPWR _20719_/X sky130_fd_sc_hd__o21a_4
X_23507_ _24082_/CLK _21989_/X VGND VGND VPWR VPWR _23507_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21699_ _21519_/X _21698_/X _23672_/Q _21695_/X VGND VGND VPWR VPWR _23672_/D sky130_fd_sc_hd__o22a_4
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14028__A _14046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240_ _14252_/A _23401_/Q VGND VGND VPWR VPWR _14241_/C sky130_fd_sc_hd__or2_4
X_23438_ _23692_/CLK _23438_/D VGND VGND VPWR VPWR _15677_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14171_ _15032_/A _14171_/B _14170_/X VGND VGND VPWR VPWR _14171_/X sky130_fd_sc_hd__or3_4
XFILLER_10_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23369_ _23910_/CLK _23369_/D VGND VGND VPWR VPWR _23369_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17339__A _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21464__B2 _21460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12771__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13122_ _13098_/A _13122_/B VGND VGND VPWR VPWR _13124_/B sky130_fd_sc_hd__or2_4
XANTENNA__19409__A1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13053_ _12211_/X _13123_/B VGND VGND VPWR VPWR _13054_/C sky130_fd_sc_hd__or2_4
X_17930_ _17798_/X _17923_/X _17823_/X _17929_/X VGND VGND VPWR VPWR _17930_/X sky130_fd_sc_hd__o22a_4
X_12004_ _11971_/A _11814_/B VGND VGND VPWR VPWR _12005_/C sky130_fd_sc_hd__or2_4
XANTENNA__21767__A2 _21762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17861_ _17861_/A VGND VGND VPWR VPWR _17862_/A sky130_fd_sc_hd__buf_2
XFILLER_61_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16812_ _16077_/A _16780_/X _16811_/X VGND VGND VPWR VPWR _16812_/X sky130_fd_sc_hd__and3_4
X_19600_ _19800_/B _19600_/B VGND VGND VPWR VPWR _19600_/X sky130_fd_sc_hd__or2_4
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17074__A _17224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17792_ _17792_/A VGND VGND VPWR VPWR _18082_/A sky130_fd_sc_hd__buf_2
X_19531_ _19531_/A VGND VGND VPWR VPWR _19531_/X sky130_fd_sc_hd__buf_2
X_16743_ _11844_/X _11620_/X _16712_/X _11598_/X _16742_/X VGND VGND VPWR VPWR _16743_/X
+ sky130_fd_sc_hd__a32o_4
X_13955_ _13955_/A _13955_/B _13955_/C VGND VGND VPWR VPWR _13956_/C sky130_fd_sc_hd__and3_4
XFILLER_93_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22192__A2 _22186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12906_ _12910_/A _12904_/X _12905_/X VGND VGND VPWR VPWR _12907_/C sky130_fd_sc_hd__and3_4
X_19462_ _19462_/A VGND VGND VPWR VPWR _19462_/X sky130_fd_sc_hd__buf_2
X_16674_ _16652_/A _16672_/X _16674_/C VGND VGND VPWR VPWR _16674_/X sky130_fd_sc_hd__and3_4
XFILLER_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12011__A _12011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13886_ _13886_/A _13886_/B _13886_/C VGND VGND VPWR VPWR _13886_/X sky130_fd_sc_hd__or3_4
XFILLER_34_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18413_ _17699_/X _18352_/B VGND VGND VPWR VPWR _18413_/Y sky130_fd_sc_hd__nand2_4
X_15625_ _15637_/A _23403_/Q VGND VGND VPWR VPWR _15625_/X sky130_fd_sc_hd__or2_4
X_12837_ _12837_/A _12837_/B _12837_/C VGND VGND VPWR VPWR _12837_/X sky130_fd_sc_hd__and3_4
X_19393_ _19389_/X _18385_/X _19392_/X _24206_/Q VGND VGND VPWR VPWR _19393_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18344_ _16974_/A VGND VGND VPWR VPWR _18344_/X sky130_fd_sc_hd__buf_2
XFILLER_15_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15556_ _15556_/A _15556_/B VGND VGND VPWR VPWR _15557_/C sky130_fd_sc_hd__or2_4
X_12768_ _12816_/A _12768_/B VGND VGND VPWR VPWR _12769_/C sky130_fd_sc_hd__or2_4
XANTENNA__21152__B1 _14379_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14556_/A _14505_/X _14506_/X VGND VGND VPWR VPWR _14507_/X sky130_fd_sc_hd__and3_4
X_11719_ _11692_/X _11705_/X _11718_/X VGND VGND VPWR VPWR _11719_/X sky130_fd_sc_hd__and3_4
X_18275_ _17587_/X _18274_/X VGND VGND VPWR VPWR _18275_/X sky130_fd_sc_hd__and2_4
XFILLER_37_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19729__A _19517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15041__B _23775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15487_ _15487_/A _15487_/B VGND VGND VPWR VPWR _15487_/X sky130_fd_sc_hd__or2_4
X_12699_ _15689_/A _12799_/B VGND VGND VPWR VPWR _12699_/X sky130_fd_sc_hd__or2_4
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17226_ _17160_/X _17219_/X _17825_/A _17225_/X VGND VGND VPWR VPWR _17226_/Y sky130_fd_sc_hd__a22oi_4
X_14438_ _12533_/A _14433_/X _14437_/X VGND VGND VPWR VPWR _14438_/X sky130_fd_sc_hd__or3_4
XANTENNA__24455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22155__A _22162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17157_ _17157_/A VGND VGND VPWR VPWR _17157_/X sky130_fd_sc_hd__buf_2
X_14369_ _15615_/A _14293_/B VGND VGND VPWR VPWR _14370_/C sky130_fd_sc_hd__or2_4
XANTENNA__12681__A _11618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16153__A _11852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16108_ _16108_/A _23991_/Q VGND VGND VPWR VPWR _16108_/X sky130_fd_sc_hd__or2_4
XFILLER_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17088_ _17088_/A _17073_/B VGND VGND VPWR VPWR _17088_/X sky130_fd_sc_hd__or2_4
X_16039_ _16039_/A _16039_/B _16038_/X VGND VGND VPWR VPWR _16043_/B sky130_fd_sc_hd__and3_4
XFILLER_48_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21207__B2 _21201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19464__A _19742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21758__A2 _21755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18084__B1 _18082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20403__A _20403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19729_ _19517_/A _19729_/B _19729_/C VGND VGND VPWR VPWR _19730_/D sky130_fd_sc_hd__or3_4
XFILLER_38_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13017__A _13017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22740_ SYSTICKCLKDIV[6] VGND VGND VPWR VPWR _22740_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21930__A2 _21924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22671_ _22671_/A VGND VGND VPWR VPWR _22686_/A sky130_fd_sc_hd__buf_2
XFILLER_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16328__A _16365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12856__A _11912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21622_ _21560_/X _21619_/X _23719_/Q _21616_/X VGND VGND VPWR VPWR _21622_/X sky130_fd_sc_hd__o22a_4
X_24410_ _24277_/CLK _24410_/D HRESETn VGND VGND VPWR VPWR _24410_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15232__A _14243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21553_ _20748_/A VGND VGND VPWR VPWR _21553_/X sky130_fd_sc_hd__buf_2
X_24341_ _24334_/CLK _24341_/D HRESETn VGND VGND VPWR VPWR _18982_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__21694__B2 _21688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20504_ _24244_/Q VGND VGND VPWR VPWR _20504_/Y sky130_fd_sc_hd__inv_2
X_24272_ _23326_/CLK _19264_/X HRESETn VGND VGND VPWR VPWR _24272_/Q sky130_fd_sc_hd__dfrtp_4
X_21484_ _21455_/A VGND VGND VPWR VPWR _21484_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23223_ _23313_/CLK _22481_/X VGND VGND VPWR VPWR _16226_/B sky130_fd_sc_hd__dfxtp_4
X_20435_ _18124_/X _20424_/X _20290_/X _20434_/Y VGND VGND VPWR VPWR _20436_/A sky130_fd_sc_hd__a211o_4
XFILLER_10_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13923__A2 _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12591__A _12935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21446__B2 _21401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24125__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21997__A2 _21995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23154_ _23826_/CLK _23154_/D VGND VGND VPWR VPWR _13089_/B sky130_fd_sc_hd__dfxtp_4
X_20366_ _20502_/A _20365_/X VGND VGND VPWR VPWR _20366_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__18862__A2 _18834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22105_ _20573_/A VGND VGND VPWR VPWR _22105_/X sky130_fd_sc_hd__buf_2
XANTENNA__19374__A _19370_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23085_ _23922_/CLK _22695_/X VGND VGND VPWR VPWR _15835_/B sky130_fd_sc_hd__dfxtp_4
X_20297_ _20297_/A VGND VGND VPWR VPWR _20297_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21749__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22036_ _21811_/X _22031_/X _12542_/B _22035_/X VGND VGND VPWR VPWR _23477_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21409__A _21401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19811__A1 _19800_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11935__A _16121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15407__A _13630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14311__A _15536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15126__B _15126_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23987_ _23987_/CLK _21134_/X VGND VGND VPWR VPWR _23987_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22174__A2 _22172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13740_ _11664_/A _13722_/X _13740_/C VGND VGND VPWR VPWR _13772_/B sky130_fd_sc_hd__or3_4
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22938_ _22978_/A VGND VGND VPWR VPWR _22962_/A sky130_fd_sc_hd__buf_2
XANTENNA__20185__A1 _18755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20185__B2 _19929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14965__B _14898_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21144__A _21130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13671_ _12233_/X _13766_/B VGND VGND VPWR VPWR _13671_/X sky130_fd_sc_hd__or2_4
XFILLER_38_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22869_ _22872_/A _22869_/B VGND VGND VPWR VPWR HWDATA[27] sky130_fd_sc_hd__nor2_4
XANTENNA__12766__A _12765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15410_ _12211_/A _15410_/B VGND VGND VPWR VPWR _15411_/C sky130_fd_sc_hd__or2_4
XANTENNA__11670__A _11670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12622_ _15512_/A VGND VGND VPWR VPWR _12622_/X sky130_fd_sc_hd__buf_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16390_ _15999_/X _16390_/B VGND VGND VPWR VPWR _16390_/X sky130_fd_sc_hd__or2_4
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24364__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15341_ _15325_/X _15339_/X _15341_/C VGND VGND VPWR VPWR _15345_/B sky130_fd_sc_hd__and3_4
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _12553_/A _12660_/B VGND VGND VPWR VPWR _12555_/B sky130_fd_sc_hd__or2_4
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19549__A _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11504_ _24320_/Q _24319_/Q VGND VGND VPWR VPWR _11504_/Y sky130_fd_sc_hd__nor2_4
X_18060_ _18011_/X _18014_/B _18058_/Y _18016_/X _23027_/B VGND VGND VPWR VPWR _18060_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_20_0_HCLK clkbuf_6_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15272_ _12531_/A _15268_/X _15271_/X VGND VGND VPWR VPWR _15272_/X sky130_fd_sc_hd__or3_4
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12484_ _13643_/A VGND VGND VPWR VPWR _13659_/A sky130_fd_sc_hd__buf_2
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17011_ _17010_/X VGND VGND VPWR VPWR _17012_/A sky130_fd_sc_hd__buf_2
X_14223_ _14039_/A _14202_/X _14222_/X VGND VGND VPWR VPWR _14261_/B sky130_fd_sc_hd__or3_4
XANTENNA__13597__A _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14154_ _15015_/A VGND VGND VPWR VPWR _14603_/A sky130_fd_sc_hd__buf_2
X_13105_ _13112_/A _23954_/Q VGND VGND VPWR VPWR _13106_/C sky130_fd_sc_hd__or2_4
XFILLER_119_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14085_ _12252_/A _14083_/X _14085_/C VGND VGND VPWR VPWR _14085_/X sky130_fd_sc_hd__and3_4
X_18962_ _18941_/X _18960_/X _18961_/Y _18946_/X VGND VGND VPWR VPWR _18962_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12006__A _12112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13036_ _13009_/A _13112_/B VGND VGND VPWR VPWR _13036_/X sky130_fd_sc_hd__or2_4
X_17913_ _17911_/X _17197_/X _17912_/X _17177_/X VGND VGND VPWR VPWR _17913_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__21319__A _21319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18893_ _17181_/X _18891_/X _24372_/Q _18892_/X VGND VGND VPWR VPWR _18893_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19802__A1 _19754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16420__B _16489_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17844_ _17800_/A _17840_/Y _17812_/A _17843_/Y VGND VGND VPWR VPWR _17844_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14221__A _13686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11564__B IRQ[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17775_ _17001_/X _23046_/B _17003_/Y VGND VGND VPWR VPWR _17775_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15036__B _23199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14987_ _14986_/X VGND VGND VPWR VPWR _14988_/A sky130_fd_sc_hd__inv_2
X_16726_ _16689_/A _16726_/B _16726_/C VGND VGND VPWR VPWR _16726_/X sky130_fd_sc_hd__or3_4
X_19514_ _19561_/A VGND VGND VPWR VPWR _19630_/A sky130_fd_sc_hd__inv_2
XANTENNA__17532__A _17531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13938_ _13959_/A _24010_/Q VGND VGND VPWR VPWR _13940_/B sky130_fd_sc_hd__or2_4
XFILLER_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18347__B _16999_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21912__A2 _21908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19445_ _19445_/A VGND VGND VPWR VPWR _19445_/X sky130_fd_sc_hd__buf_2
XFILLER_39_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16657_ _16662_/A _16657_/B VGND VGND VPWR VPWR _16657_/X sky130_fd_sc_hd__or2_4
X_13869_ _13911_/A _13869_/B _13869_/C VGND VGND VPWR VPWR _13869_/X sky130_fd_sc_hd__and3_4
XANTENNA__16148__A _15937_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_102_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR _23383_/CLK sky130_fd_sc_hd__clkbuf_1
X_15608_ _15632_/A _15539_/B VGND VGND VPWR VPWR _15610_/B sky130_fd_sc_hd__or2_4
XFILLER_90_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19376_ _19374_/X _18133_/X _19374_/X _24214_/Q VGND VGND VPWR VPWR _19376_/X sky130_fd_sc_hd__a2bb2o_4
X_16588_ _12020_/A _16586_/X _16588_/C VGND VGND VPWR VPWR _16592_/B sky130_fd_sc_hd__and3_4
XANTENNA__21125__B1 _23993_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18327_ _18327_/A _18326_/Y VGND VGND VPWR VPWR _18327_/X sky130_fd_sc_hd__and2_4
XFILLER_52_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15539_ _14431_/A _15539_/B VGND VGND VPWR VPWR _15541_/B sky130_fd_sc_hd__or2_4
XANTENNA__15987__A _16095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22873__B1 _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18258_ _17668_/Y _18165_/X _17668_/Y _18165_/X VGND VGND VPWR VPWR _18258_/X sky130_fd_sc_hd__a2bb2o_4
X_17209_ _17156_/Y _17173_/X _13920_/X _17145_/X VGND VGND VPWR VPWR _17209_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21428__B2 _21423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18189_ _18189_/A VGND VGND VPWR VPWR _18189_/X sky130_fd_sc_hd__buf_2
X_20220_ _20846_/B HRDATA[7] _19885_/Y VGND VGND VPWR VPWR _20220_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21979__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20151_ _20143_/Y _20144_/Y _11554_/X _20150_/X VGND VGND VPWR VPWR _20151_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16611__A _16616_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23951__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21229__A _21799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20082_ _20090_/D _20071_/X _20076_/X _11626_/Y VGND VGND VPWR VPWR _20082_/X sky130_fd_sc_hd__or4_4
XFILLER_97_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23910_ _23910_/CLK _23910_/D VGND VGND VPWR VPWR _14292_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11755__A _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21600__B2 _21595_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14131__A _11954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23841_ _23487_/CLK _23841_/D VGND VGND VPWR VPWR _15180_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19557__B1 HRDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17442__A _17442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13970__A _12509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20984_ _20844_/A HRDATA[16] VGND VGND VPWR VPWR _20984_/X sky130_fd_sc_hd__or2_4
X_23772_ _23931_/CLK _21511_/X VGND VGND VPWR VPWR _23772_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21903__A2 _21901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22723_ _22723_/A _22723_/B VGND VGND VPWR VPWR _22723_/Y sky130_fd_sc_hd__nor2_4
XFILLER_81_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12586__A _12981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18780__A1 _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24457__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22654_ _22633_/A VGND VGND VPWR VPWR _22654_/X sky130_fd_sc_hd__buf_2
XFILLER_80_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21605_ _21605_/A VGND VGND VPWR VPWR _21605_/X sky130_fd_sc_hd__buf_2
XANTENNA__15897__A _13494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22585_ _22413_/X _22579_/X _23156_/Q _22583_/X VGND VGND VPWR VPWR _22585_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22864__B1 _17411_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21667__B2 _21666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24306__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24324_ _24305_/CLK _24324_/D HRESETn VGND VGND VPWR VPWR _11509_/A sky130_fd_sc_hd__dfstp_4
X_21536_ _20574_/A VGND VGND VPWR VPWR _21536_/X sky130_fd_sc_hd__buf_2
XFILLER_103_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21467_ _21467_/A VGND VGND VPWR VPWR _21467_/X sky130_fd_sc_hd__buf_2
X_24255_ _24290_/CLK _24255_/D HRESETn VGND VGND VPWR VPWR _24255_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20418_ _20418_/A VGND VGND VPWR VPWR _21804_/A sky130_fd_sc_hd__buf_2
X_23206_ _23781_/CLK _23206_/D VGND VGND VPWR VPWR _14417_/B sky130_fd_sc_hd__dfxtp_4
X_21398_ _21348_/A _21784_/B _21348_/C _21734_/B VGND VGND VPWR VPWR _21398_/X sky130_fd_sc_hd__or4_4
X_24186_ _24223_/CLK _19586_/X HRESETn VGND VGND VPWR VPWR _17273_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14025__B _14025_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20349_ _20332_/A _20348_/X VGND VGND VPWR VPWR _20349_/Y sky130_fd_sc_hd__nor2_4
X_23137_ _23233_/CLK _23137_/D VGND VGND VPWR VPWR _15149_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_49_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23068_ VGND VGND VPWR VPWR _23068_/HI HTRANS[0] sky130_fd_sc_hd__conb_1
XFILLER_1_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18599__A1 _16919_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22395__A2 _22392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16240__B _16240_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14910_ _14880_/A _23776_/Q VGND VGND VPWR VPWR _14911_/C sky130_fd_sc_hd__or2_4
X_22019_ _22052_/A VGND VGND VPWR VPWR _22035_/A sky130_fd_sc_hd__inv_2
XFILLER_118_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11665__A _12957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18599__B2 _18598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15137__A _14098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15890_ _13557_/A _15882_/X _15889_/X VGND VGND VPWR VPWR _15890_/X sky130_fd_sc_hd__and3_4
XFILLER_114_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14041__A _14813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14841_ _14841_/A _14769_/B VGND VGND VPWR VPWR _14841_/X sky130_fd_sc_hd__or2_4
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17560_ _16155_/X VGND VGND VPWR VPWR _17560_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14772_ _15443_/A _14772_/B VGND VGND VPWR VPWR _14774_/B sky130_fd_sc_hd__or2_4
X_11984_ _11901_/X _23582_/Q VGND VGND VPWR VPWR _11985_/C sky130_fd_sc_hd__or2_4
XFILLER_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16511_ _11673_/X _16503_/X _16511_/C VGND VGND VPWR VPWR _16512_/C sky130_fd_sc_hd__and3_4
X_13723_ _15486_/A _13723_/B VGND VGND VPWR VPWR _13723_/X sky130_fd_sc_hd__or2_4
X_17491_ _17488_/X VGND VGND VPWR VPWR _17517_/B sky130_fd_sc_hd__inv_2
XANTENNA__12496__A _12496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18771__A1 _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19230_ _19230_/A _19247_/A VGND VGND VPWR VPWR _19245_/A sky130_fd_sc_hd__and2_4
XFILLER_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16442_ _11982_/A _16419_/X _16426_/X _16433_/X _16441_/X VGND VGND VPWR VPWR _16442_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13654_ _13654_/A VGND VGND VPWR VPWR _15431_/A sky130_fd_sc_hd__buf_2
XFILLER_32_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12605_ _12605_/A VGND VGND VPWR VPWR _12652_/A sky130_fd_sc_hd__buf_2
X_19161_ _19129_/B VGND VGND VPWR VPWR _19161_/Y sky130_fd_sc_hd__inv_2
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21602__A _21602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21658__A1 _21536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16373_ _11658_/X _16373_/B _16373_/C VGND VGND VPWR VPWR _16374_/A sky130_fd_sc_hd__and3_4
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21658__B2 _21652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13585_ _12842_/X _12994_/Y _12843_/X VGND VGND VPWR VPWR _13585_/Y sky130_fd_sc_hd__o21ai_4
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18112_ _17800_/A _17922_/Y _17914_/X _17928_/Y VGND VGND VPWR VPWR _18112_/X sky130_fd_sc_hd__o22a_4
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15324_ _15334_/A _15324_/B _15324_/C VGND VGND VPWR VPWR _15330_/B sky130_fd_sc_hd__and3_4
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12536_ _12905_/A _12648_/B VGND VGND VPWR VPWR _12537_/C sky130_fd_sc_hd__or2_4
X_19092_ _19092_/A VGND VGND VPWR VPWR _19092_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18043_ _17259_/A _18042_/Y VGND VGND VPWR VPWR _18043_/X sky130_fd_sc_hd__and2_4
X_15255_ _14315_/A _15255_/B VGND VGND VPWR VPWR _15255_/X sky130_fd_sc_hd__or2_4
X_12467_ _13651_/A VGND VGND VPWR VPWR _13019_/A sky130_fd_sc_hd__buf_2
X_14206_ _14206_/A _14206_/B _14205_/X VGND VGND VPWR VPWR _14212_/B sky130_fd_sc_hd__and3_4
X_15186_ _14644_/A _15125_/B VGND VGND VPWR VPWR _15186_/X sky130_fd_sc_hd__or2_4
X_12398_ _12398_/A _12396_/X _12398_/C VGND VGND VPWR VPWR _12398_/X sky130_fd_sc_hd__and3_4
XFILLER_119_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14137_ _14995_/A VGND VGND VPWR VPWR _14145_/A sky130_fd_sc_hd__buf_2
XFILLER_10_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17527__A _12674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20633__A2 _20621_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21830__B2 _21824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19994_ _19994_/A VGND VGND VPWR VPWR _19994_/X sky130_fd_sc_hd__buf_2
XFILLER_99_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_27_0_HCLK clkbuf_6_13_0_HCLK/X VGND VGND VPWR VPWR _23233_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14068_ _14068_/A _23626_/Q VGND VGND VPWR VPWR _14068_/X sky130_fd_sc_hd__or2_4
X_18945_ _19027_/A VGND VGND VPWR VPWR _18999_/A sky130_fd_sc_hd__buf_2
XANTENNA__23204__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13774__B _13772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13019_ _13019_/A _23922_/Q VGND VGND VPWR VPWR _13021_/B sky130_fd_sc_hd__or2_4
XANTENNA__19742__A _19742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18876_ _18898_/A VGND VGND VPWR VPWR _18877_/A sky130_fd_sc_hd__inv_2
XFILLER_80_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20888__A _20888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17827_ _17826_/X _17176_/X _17815_/X _17193_/X VGND VGND VPWR VPWR _17827_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18358__A _18418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22138__A2 _22137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13790__A _13813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17758_ _17758_/A _17758_/B VGND VGND VPWR VPWR _17758_/X sky130_fd_sc_hd__or2_4
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21346__B1 _23871_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20400__B _20400_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16709_ _11875_/X _16709_/B _16709_/C VGND VGND VPWR VPWR _16709_/X sky130_fd_sc_hd__and3_4
X_17689_ _16945_/Y _17469_/Y VGND VGND VPWR VPWR _17690_/A sky130_fd_sc_hd__or2_4
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21897__B2 _21891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19428_ _19428_/A VGND VGND VPWR VPWR _19429_/A sky130_fd_sc_hd__buf_2
XANTENNA__24470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19359_ _19370_/A VGND VGND VPWR VPWR _19359_/X sky130_fd_sc_hd__buf_2
XANTENNA__21649__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16606__A _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15510__A _13737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22370_ _22127_/X _22368_/X _23272_/Q _22365_/X VGND VGND VPWR VPWR _23272_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16525__B1 _16524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21321_ _21249_/X _21319_/X _13104_/B _21316_/X VGND VGND VPWR VPWR _21321_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19917__A _22723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18821__A _18835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21252_ _21251_/X _21247_/X _13162_/B _21242_/X VGND VGND VPWR VPWR _21252_/X sky130_fd_sc_hd__o22a_4
X_24040_ _23591_/CLK _24040_/D VGND VGND VPWR VPWR _13745_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_11_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22074__B2 _22072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20203_ _20202_/X VGND VGND VPWR VPWR _20203_/X sky130_fd_sc_hd__buf_2
XANTENNA__20085__B1 _19303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13965__A _12302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21183_ _21183_/A VGND VGND VPWR VPWR _21183_/X sky130_fd_sc_hd__buf_2
XFILLER_116_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16341__A _16188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20134_ _20134_/A VGND VGND VPWR VPWR _20134_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22377__A2 _22375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20065_ _20065_/A VGND VGND VPWR VPWR _24118_/D sky130_fd_sc_hd__inv_2
XANTENNA__18450__B1 _18398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14796__A _13710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17172__A _17171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23824_ _23920_/CLK _23824_/D VGND VGND VPWR VPWR _13326_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_57_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21888__A1 _21816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23755_ _24011_/CLK _23755_/D VGND VGND VPWR VPWR _15530_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21888__B2 _21884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20967_ _20966_/Y _20471_/A VGND VGND VPWR VPWR _20967_/X sky130_fd_sc_hd__or2_4
XFILLER_14_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19950__B1 _17874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22706_ _20870_/A _22700_/X _14547_/B _22704_/X VGND VGND VPWR VPWR _22706_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23686_ _23845_/CLK _23686_/D VGND VGND VPWR VPWR _14330_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20560__A1 _20425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20898_ _19734_/Y _20850_/Y _20895_/B _20821_/B VGND VGND VPWR VPWR _20898_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22518__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20560__B2 _20473_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22637_ _22415_/X _22636_/X _12965_/B _22633_/X VGND VGND VPWR VPWR _23123_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24140__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16516__A _16444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15420__A _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13370_ _13370_/A _13370_/B _13370_/C VGND VGND VPWR VPWR _13371_/C sky130_fd_sc_hd__or3_4
XFILLER_35_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22568_ _22583_/A VGND VGND VPWR VPWR _22576_/A sky130_fd_sc_hd__buf_2
XFILLER_16_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12321_ _12435_/A VGND VGND VPWR VPWR _12740_/A sky130_fd_sc_hd__buf_2
X_24307_ _24301_/CLK _24307_/D HRESETn VGND VGND VPWR VPWR _19128_/A sky130_fd_sc_hd__dfrtp_4
X_21519_ _21804_/A VGND VGND VPWR VPWR _21519_/X sky130_fd_sc_hd__buf_2
X_22499_ _22437_/X _22493_/X _14066_/B _22497_/X VGND VGND VPWR VPWR _23210_/D sky130_fd_sc_hd__o22a_4
X_15040_ _15013_/A _23071_/Q VGND VGND VPWR VPWR _15040_/X sky130_fd_sc_hd__or2_4
X_12252_ _12252_/A VGND VGND VPWR VPWR _15448_/A sky130_fd_sc_hd__buf_2
X_24238_ _24239_/CLK _24238_/D HRESETn VGND VGND VPWR VPWR _24238_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22065__B2 _22020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22253__A _22286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16819__A1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13875__A _13910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12183_ _16077_/A _12183_/B _12183_/C VGND VGND VPWR VPWR _12184_/A sky130_fd_sc_hd__and3_4
X_24169_ _23584_/CLK _24169_/D HRESETn VGND VGND VPWR VPWR _19823_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_1_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16991_ _16991_/A _16991_/B VGND VGND VPWR VPWR _16992_/A sky130_fd_sc_hd__or2_4
X_15942_ _16095_/A _15942_/B _15942_/C VGND VGND VPWR VPWR _15942_/X sky130_fd_sc_hd__or3_4
X_18730_ _17912_/X _18729_/X _17801_/X _17809_/X VGND VGND VPWR VPWR _18730_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_77_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19562__A _19784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18661_ _17966_/X _17334_/X _18107_/A _17616_/X VGND VGND VPWR VPWR _18662_/B sky130_fd_sc_hd__o22a_4
XFILLER_23_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21040__A2 _21037_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15873_ _13494_/X _15869_/X _15873_/C VGND VGND VPWR VPWR _15874_/C sky130_fd_sc_hd__or3_4
XFILLER_37_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18178__A _18242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14824_ _14050_/A _14822_/X _14824_/C VGND VGND VPWR VPWR _14824_/X sky130_fd_sc_hd__and3_4
X_17612_ _17221_/Y _17135_/A VGND VGND VPWR VPWR _17612_/X sky130_fd_sc_hd__or2_4
X_18592_ _18697_/A _17619_/A _18588_/X _18591_/Y VGND VGND VPWR VPWR _18592_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21328__B1 _23885_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17543_ _17543_/A _17457_/B VGND VGND VPWR VPWR _17543_/X sky130_fd_sc_hd__and2_4
XFILLER_75_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14755_ _12439_/A _14819_/B VGND VGND VPWR VPWR _14757_/B sky130_fd_sc_hd__or2_4
XANTENNA__15314__B _15253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11967_ _11886_/X VGND VGND VPWR VPWR _12022_/A sky130_fd_sc_hd__buf_2
XANTENNA__21879__B2 _21877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18906__A _18877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13706_ _13706_/A VGND VGND VPWR VPWR _13893_/A sky130_fd_sc_hd__buf_2
X_17474_ _17472_/Y _17473_/X VGND VGND VPWR VPWR _18152_/A sky130_fd_sc_hd__or2_4
X_14686_ _15628_/A _14678_/X _14685_/X VGND VGND VPWR VPWR _14686_/X sky130_fd_sc_hd__and3_4
X_11898_ _12444_/A VGND VGND VPWR VPWR _13463_/A sky130_fd_sc_hd__buf_2
XANTENNA__22428__A _22416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16425_ _16087_/X _16423_/X _16424_/X VGND VGND VPWR VPWR _16426_/C sky130_fd_sc_hd__and3_4
X_19213_ _19213_/A _19213_/B VGND VGND VPWR VPWR _19214_/B sky130_fd_sc_hd__and2_4
XFILLER_60_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13637_ _15411_/A _13634_/X _13637_/C VGND VGND VPWR VPWR _13638_/C sky130_fd_sc_hd__and3_4
XFILLER_44_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16426__A _15929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12954__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19144_ _19137_/A _19136_/X _19143_/Y VGND VGND VPWR VPWR _19144_/X sky130_fd_sc_hd__o21a_4
X_16356_ _16322_/A _16293_/B VGND VGND VPWR VPWR _16356_/X sky130_fd_sc_hd__or2_4
XFILLER_13_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13568_ _13561_/A _13568_/B VGND VGND VPWR VPWR _13568_/X sky130_fd_sc_hd__or2_4
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15307_ _13927_/A _15307_/B VGND VGND VPWR VPWR _15307_/X sky130_fd_sc_hd__or2_4
X_12519_ _12518_/X _12639_/B VGND VGND VPWR VPWR _12519_/X sky130_fd_sc_hd__or2_4
X_19075_ _19060_/X _19073_/X _19074_/X _11511_/A VGND VGND VPWR VPWR _24326_/D sky130_fd_sc_hd__a2bb2o_4
X_16287_ _15934_/X _16365_/B VGND VGND VPWR VPWR _16287_/X sky130_fd_sc_hd__or2_4
X_13499_ _13550_/A _13496_/X _13498_/X VGND VGND VPWR VPWR _13499_/X sky130_fd_sc_hd__and3_4
XANTENNA__17180__B1 _12676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18641__A _18640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18026_ _18295_/A VGND VGND VPWR VPWR _18241_/A sky130_fd_sc_hd__buf_2
X_15238_ _14345_/A _15238_/B _15237_/X VGND VGND VPWR VPWR _15238_/X sky130_fd_sc_hd__and3_4
XANTENNA__15984__B _15984_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24152__CLK _24223_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15169_ _14113_/A _15240_/B VGND VGND VPWR VPWR _15169_/X sky130_fd_sc_hd__or2_4
XANTENNA__21803__B2 _21800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16161__A _16194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19977_ _19977_/A VGND VGND VPWR VPWR _19977_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22359__A2 _22354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18928_ _18927_/X VGND VGND VPWR VPWR _18928_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21031__A2 _21030_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21507__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18859_ _14851_/X _18855_/X _24387_/Q _18856_/X VGND VGND VPWR VPWR _18859_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17704__B _17404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21870_ _21869_/X VGND VGND VPWR VPWR _21870_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20821_ HRDATA[7] _20821_/B VGND VGND VPWR VPWR _20823_/B sky130_fd_sc_hd__or2_4
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18735__A1 _18424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13025__A _13025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22531__A2 _22529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19932__B1 _23064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23540_ _24084_/CLK _21937_/X VGND VGND VPWR VPWR _12803_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_93_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20752_ _18577_/Y VGND VGND VPWR VPWR _20913_/A sky130_fd_sc_hd__buf_2
XANTENNA__20542__A1 _20448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21242__A _21242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20683_ _24396_/Q _20623_/X _24428_/Q _20682_/X VGND VGND VPWR VPWR _20683_/X sky130_fd_sc_hd__o22a_4
X_23471_ _23311_/CLK _22044_/X VGND VGND VPWR VPWR _23471_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12864__A _12518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16336__A _11727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22422_ _20590_/A VGND VGND VPWR VPWR _22422_/X sky130_fd_sc_hd__buf_2
XANTENNA__21098__A2 _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22295__B2 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19696__C1 _19695_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22353_ _22098_/X _22347_/X _12784_/B _22351_/X VGND VGND VPWR VPWR _23284_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17710__A2 _17413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21304_ _21300_/A VGND VGND VPWR VPWR _21319_/A sky130_fd_sc_hd__buf_2
X_22284_ _22119_/X _22279_/X _23339_/Q _22283_/X VGND VGND VPWR VPWR _22284_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22047__B2 _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15894__B _15838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22073__A _20276_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22598__A2 _22593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21235_ _21247_/A VGND VGND VPWR VPWR _21235_/X sky130_fd_sc_hd__buf_2
X_24023_ _23316_/CLK _21077_/X VGND VGND VPWR VPWR _16175_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_30_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13695__A _13890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16071__A _16071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21166_ _21165_/X VGND VGND VPWR VPWR _21166_/X sky130_fd_sc_hd__buf_2
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20117_ _20086_/A _20116_/X _20087_/Y VGND VGND VPWR VPWR _20117_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19382__A _19382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_10_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR _23363_/CLK sky130_fd_sc_hd__clkbuf_1
X_21097_ _20779_/X _21096_/X _24009_/Q _21093_/X VGND VGND VPWR VPWR _21097_/X sky130_fd_sc_hd__o22a_4
XFILLER_63_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12104__A _12100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_73_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR _23100_/CLK sky130_fd_sc_hd__clkbuf_1
X_20048_ _20000_/A VGND VGND VPWR VPWR _20048_/X sky130_fd_sc_hd__buf_2
XFILLER_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20321__A _20493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11943__A _11943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15415__A _13632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12870_ _12870_/A _12870_/B _12869_/X VGND VGND VPWR VPWR _12870_/X sky130_fd_sc_hd__and3_4
XANTENNA__24392__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12758__B _12758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11821_ _11821_/A _23710_/Q VGND VGND VPWR VPWR _11821_/X sky130_fd_sc_hd__or2_4
X_23807_ _23130_/CLK _23807_/D VGND VGND VPWR VPWR _23807_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21999_ _21985_/A VGND VGND VPWR VPWR _21999_/X sky130_fd_sc_hd__buf_2
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19923__B1 _22723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14533_/A _14470_/B VGND VGND VPWR VPWR _14540_/X sky130_fd_sc_hd__or2_4
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11691_/X VGND VGND VPWR VPWR _11820_/A sky130_fd_sc_hd__buf_2
X_23738_ _23706_/CLK _21596_/X VGND VGND VPWR VPWR _16384_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21730__B1 _23649_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _12862_/A _14469_/X _14470_/X VGND VGND VPWR VPWR _14471_/X sky130_fd_sc_hd__and3_4
XFILLER_14_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _13415_/A VGND VGND VPWR VPWR _16198_/A sky130_fd_sc_hd__buf_2
X_23669_ _24021_/CLK _21703_/X VGND VGND VPWR VPWR _12627_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16194_/A _16208_/X _16209_/X VGND VGND VPWR VPWR _16210_/X sky130_fd_sc_hd__and3_4
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _13422_/A _13422_/B _13422_/C VGND VGND VPWR VPWR _13423_/C sky130_fd_sc_hd__or3_4
XANTENNA__15150__A _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17190_ _17160_/A VGND VGND VPWR VPWR _17817_/A sky130_fd_sc_hd__buf_2
XFILLER_35_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16141_ _16107_/A _16226_/B VGND VGND VPWR VPWR _16143_/B sky130_fd_sc_hd__or2_4
X_13353_ _13352_/X _13282_/B VGND VGND VPWR VPWR _13353_/X sky130_fd_sc_hd__or2_4
XFILLER_6_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17162__B1 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12304_ _15558_/A VGND VGND VPWR VPWR _12713_/A sky130_fd_sc_hd__buf_2
X_16072_ _16072_/A _23640_/Q VGND VGND VPWR VPWR _16072_/X sky130_fd_sc_hd__or2_4
X_13284_ _13283_/X _23504_/Q VGND VGND VPWR VPWR _13284_/X sky130_fd_sc_hd__or2_4
X_15023_ _15023_/A _15023_/B VGND VGND VPWR VPWR _15024_/C sky130_fd_sc_hd__or2_4
X_19900_ _22978_/A VGND VGND VPWR VPWR _22968_/A sky130_fd_sc_hd__inv_2
XANTENNA__22589__A2 _22586_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12235_ _12235_/A VGND VGND VPWR VPWR _12693_/A sky130_fd_sc_hd__buf_2
XFILLER_83_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19831_ _21582_/A VGND VGND VPWR VPWR _21348_/B sky130_fd_sc_hd__buf_2
X_12166_ _11772_/X _12158_/X _12166_/C VGND VGND VPWR VPWR _12166_/X sky130_fd_sc_hd__and3_4
XFILLER_29_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19762_ _19712_/A HRDATA[1] VGND VGND VPWR VPWR _19762_/X sky130_fd_sc_hd__and2_4
X_12097_ _12093_/A _23485_/Q VGND VGND VPWR VPWR _12099_/B sky130_fd_sc_hd__or2_4
X_16974_ _16974_/A _16974_/B VGND VGND VPWR VPWR _16975_/B sky130_fd_sc_hd__or2_4
XFILLER_49_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21549__B1 _15463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17217__A1 _17132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18713_ _18713_/A _17808_/X _18711_/X VGND VGND VPWR VPWR _18713_/X sky130_fd_sc_hd__or3_4
X_15925_ _15391_/X _15914_/X _15782_/X _15924_/Y VGND VGND VPWR VPWR _15926_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22210__B2 _22205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19693_ _19582_/A _19668_/X _19625_/Y VGND VGND VPWR VPWR _19693_/X sky130_fd_sc_hd__a21o_4
XANTENNA__20231__A _20421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11853__A _11852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15325__A _14177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15856_ _13548_/X _15795_/B VGND VGND VPWR VPWR _15856_/X sky130_fd_sc_hd__or2_4
X_18644_ _18644_/A _18609_/Y VGND VGND VPWR VPWR _18644_/X sky130_fd_sc_hd__and2_4
XFILLER_76_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20772__A1 _18528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14807_ _12599_/A _14807_/B _14806_/X VGND VGND VPWR VPWR _14807_/X sky130_fd_sc_hd__and3_4
XFILLER_80_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15044__B _23839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15787_ _12443_/A _15848_/B VGND VGND VPWR VPWR _15787_/X sky130_fd_sc_hd__or2_4
X_18575_ _17745_/C _17745_/B _17720_/X VGND VGND VPWR VPWR _18575_/X sky130_fd_sc_hd__o21a_4
X_12999_ _12852_/A _23506_/Q VGND VGND VPWR VPWR _12999_/X sky130_fd_sc_hd__or2_4
XFILLER_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18636__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14738_ _11929_/A _14734_/X _14738_/C VGND VGND VPWR VPWR _14738_/X sky130_fd_sc_hd__or3_4
X_17526_ _17456_/Y _17524_/Y _17525_/X VGND VGND VPWR VPWR _17526_/X sky130_fd_sc_hd__o21a_4
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20524__A1 _20468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22158__A _22172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14883__B _14883_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19390__B2 _24208_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17457_ _11853_/X _17457_/B VGND VGND VPWR VPWR _17457_/X sky130_fd_sc_hd__and2_4
X_14669_ _15115_/A _14663_/X _14668_/X VGND VGND VPWR VPWR _14669_/X sky130_fd_sc_hd__or3_4
XANTENNA__12684__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16408_ _16100_/X _16408_/B VGND VGND VPWR VPWR _16409_/C sky130_fd_sc_hd__or2_4
X_17388_ _17388_/A VGND VGND VPWR VPWR _17424_/B sky130_fd_sc_hd__inv_2
XANTENNA__22277__B2 _22276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16339_ _11666_/X _16321_/X _16338_/X VGND VGND VPWR VPWR _16373_/B sky130_fd_sc_hd__or3_4
X_19127_ _24306_/Q _19165_/A VGND VGND VPWR VPWR _19163_/A sky130_fd_sc_hd__and2_4
XANTENNA__19467__A _19517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17153__B1 _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23542__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19058_ _19052_/X _19055_/X _19056_/Y _19057_/X VGND VGND VPWR VPWR _19058_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22029__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12517__A1 _13491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18009_ _18198_/A VGND VGND VPWR VPWR _18009_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21020_ _21012_/X VGND VGND VPWR VPWR _21020_/X sky130_fd_sc_hd__buf_2
XFILLER_114_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21252__A2 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22621__A _22621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21237__A _20442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22971_ _22955_/X _18383_/A _22967_/X _22970_/X VGND VGND VPWR VPWR _22972_/A sky130_fd_sc_hd__a211o_4
XFILLER_68_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12859__A _12859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17759__A2 _17479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13493__A2 _11618_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15235__A _14215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11763__A _11675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21922_ _21915_/Y _21921_/X _21789_/X _21921_/X VGND VGND VPWR VPWR _23550_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19930__A _19929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22670__A2_N _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21853_ _21792_/A VGND VGND VPWR VPWR _21853_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20804_ _24423_/Q VGND VGND VPWR VPWR _20805_/A sky130_fd_sc_hd__inv_2
XFILLER_93_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21784_ _21784_/A _21784_/B _21784_/C _21784_/D VGND VGND VPWR VPWR _21784_/X sky130_fd_sc_hd__or4_4
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19381__A1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23523_ _23270_/CLK _23523_/D VGND VGND VPWR VPWR _14743_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20735_ _20681_/X _20734_/X _24362_/Q _20625_/X VGND VGND VPWR VPWR _20735_/X sky130_fd_sc_hd__o22a_4
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12594__A _12937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23454_ _23358_/CLK _23454_/D VGND VGND VPWR VPWR _11781_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20666_ _20640_/X _20652_/X _20515_/X _20665_/Y VGND VGND VPWR VPWR _20666_/X sky130_fd_sc_hd__a211o_4
XFILLER_91_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22405_ _22403_/X _22404_/X _23256_/Q _22399_/X VGND VGND VPWR VPWR _23256_/D sky130_fd_sc_hd__o22a_4
X_20597_ _20596_/Y _20521_/B VGND VGND VPWR VPWR _20597_/X sky130_fd_sc_hd__or2_4
X_23385_ _23354_/CLK _23385_/D VGND VGND VPWR VPWR _16282_/B sky130_fd_sc_hd__dfxtp_4
X_22336_ _22351_/A VGND VGND VPWR VPWR _22344_/A sky130_fd_sc_hd__buf_2
XANTENNA__11938__A _11993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22267_ _22091_/X _22265_/X _16092_/B _22262_/X VGND VGND VPWR VPWR _22267_/X sky130_fd_sc_hd__o22a_4
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _12020_/A _12020_/B _12020_/C VGND VGND VPWR VPWR _12026_/B sky130_fd_sc_hd__and3_4
X_24006_ _23845_/CLK _24006_/D VGND VGND VPWR VPWR _14278_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_117_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21218_ _21230_/A VGND VGND VPWR VPWR _21218_/X sky130_fd_sc_hd__buf_2
XANTENNA__21243__A2 _21235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22198_ _22145_/X _22193_/X _14899_/B _22162_/A VGND VGND VPWR VPWR _22198_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21149_ _20797_/X _21147_/X _13630_/B _21144_/X VGND VGND VPWR VPWR _23976_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21147__A _21118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13971_ _12217_/A _13971_/B _13971_/C VGND VGND VPWR VPWR _13971_/X sky130_fd_sc_hd__and3_4
XFILLER_47_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12769__A _12769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15710_ _11850_/A _15709_/X VGND VGND VPWR VPWR _15710_/X sky130_fd_sc_hd__and2_4
XANTENNA__11673__A _12787_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12922_ _12922_/A _12921_/X VGND VGND VPWR VPWR _12922_/X sky130_fd_sc_hd__and2_4
XFILLER_24_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15145__A _14145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16690_ _16686_/A _16754_/B VGND VGND VPWR VPWR _16692_/B sky130_fd_sc_hd__or2_4
XFILLER_73_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15641_ _13896_/A _15641_/B _15641_/C VGND VGND VPWR VPWR _15642_/C sky130_fd_sc_hd__and3_4
XFILLER_94_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12853_ _12895_/A _12929_/B VGND VGND VPWR VPWR _12854_/C sky130_fd_sc_hd__or2_4
XFILLER_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_3_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR _24208_/CLK sky130_fd_sc_hd__clkbuf_1
X_11804_ _11717_/X _21161_/A VGND VGND VPWR VPWR _11804_/X sky130_fd_sc_hd__or2_4
X_18360_ _18242_/A _17483_/X VGND VGND VPWR VPWR _18360_/Y sky130_fd_sc_hd__nor2_4
X_15572_ _12460_/A _15568_/X _15571_/X VGND VGND VPWR VPWR _15572_/X sky130_fd_sc_hd__or3_4
X_12784_ _12800_/A _12784_/B VGND VGND VPWR VPWR _12784_/X sky130_fd_sc_hd__or2_4
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15799__B _15799_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17336_/B _17310_/X VGND VGND VPWR VPWR _17311_/X sky130_fd_sc_hd__or2_4
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14554_/A _14523_/B VGND VGND VPWR VPWR _14523_/X sky130_fd_sc_hd__or2_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12995__A1 _12924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11730_/X _11732_/X _11734_/X VGND VGND VPWR VPWR _11735_/X sky130_fd_sc_hd__and3_4
X_18291_ _18129_/A VGND VGND VPWR VPWR _18291_/X sky130_fd_sc_hd__buf_2
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17242_/A VGND VGND VPWR VPWR _17259_/A sky130_fd_sc_hd__buf_2
XFILLER_70_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _15393_/A _14516_/B VGND VGND VPWR VPWR _14455_/C sky130_fd_sc_hd__or2_4
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11665_/X VGND VGND VPWR VPWR _11666_/X sky130_fd_sc_hd__buf_2
XFILLER_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22259__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13397_/X _13329_/B VGND VGND VPWR VPWR _13406_/C sky130_fd_sc_hd__or2_4
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17173_ _17173_/A VGND VGND VPWR VPWR _17173_/X sky130_fd_sc_hd__buf_2
X_14385_ _15633_/A _14289_/B VGND VGND VPWR VPWR _14385_/X sky130_fd_sc_hd__or2_4
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11597_ _11596_/X VGND VGND VPWR VPWR _11597_/X sky130_fd_sc_hd__buf_2
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16704__A _11888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16124_ _16127_/A _16124_/B VGND VGND VPWR VPWR _16126_/B sky130_fd_sc_hd__or2_4
X_13336_ _13300_/A _13336_/B VGND VGND VPWR VPWR _13336_/X sky130_fd_sc_hd__or2_4
XFILLER_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21482__A2 _21477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16423__B _16423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16055_ _16039_/A _16053_/X _16054_/X VGND VGND VPWR VPWR _16055_/X sky130_fd_sc_hd__and3_4
XANTENNA__11848__A _13682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13267_ _11671_/A _13259_/X _13266_/X VGND VGND VPWR VPWR _13268_/C sky130_fd_sc_hd__and3_4
XANTENNA__14224__A _14020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19427__A2 _19545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15006_ _15006_/A _15081_/B VGND VGND VPWR VPWR _15006_/X sky130_fd_sc_hd__or2_4
XANTENNA__17438__A1 _17338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12218_ _13632_/A VGND VGND VPWR VPWR _13796_/A sky130_fd_sc_hd__buf_2
X_13198_ _11912_/A _13196_/X _13197_/X VGND VGND VPWR VPWR _13198_/X sky130_fd_sc_hd__and3_4
XANTENNA__22431__B2 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19814_ _19442_/B _19500_/X _19740_/A _19813_/X VGND VGND VPWR VPWR _19814_/X sky130_fd_sc_hd__o22a_4
XFILLER_97_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12149_ _11824_/A _12145_/X _12148_/X VGND VGND VPWR VPWR _12149_/X sky130_fd_sc_hd__or3_4
XANTENNA__17535__A _17535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20993__A1 _20494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20993__B2 _20453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19745_ _19429_/A _19873_/B VGND VGND VPWR VPWR _19745_/X sky130_fd_sc_hd__and2_4
XFILLER_81_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16957_ _16957_/A VGND VGND VPWR VPWR _17708_/A sky130_fd_sc_hd__inv_2
XANTENNA__24243__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15055__A _15072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15908_ _15907_/X VGND VGND VPWR VPWR _15909_/B sky130_fd_sc_hd__inv_2
XFILLER_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19676_ _16997_/X _19674_/X _20800_/A _19553_/A HRDATA[8] VGND VGND VPWR VPWR _19676_/X
+ sky130_fd_sc_hd__a32o_4
X_16888_ _16834_/X _16845_/X _16879_/X _16887_/X VGND VGND VPWR VPWR _16888_/X sky130_fd_sc_hd__and4_4
XANTENNA__23095__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18627_ _18602_/Y _18604_/X _18605_/X _18626_/X VGND VGND VPWR VPWR _18628_/A sky130_fd_sc_hd__o22a_4
X_15839_ _13009_/A _15839_/B VGND VGND VPWR VPWR _15839_/X sky130_fd_sc_hd__or2_4
X_18558_ _18558_/A _18557_/X VGND VGND VPWR VPWR _18558_/X sky130_fd_sc_hd__or2_4
XANTENNA__23908__CLK _23107_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22498__B2 _22497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17509_ _17508_/X VGND VGND VPWR VPWR _18297_/B sky130_fd_sc_hd__inv_2
XANTENNA__15502__B _23788_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18489_ _17421_/A _18488_/X VGND VGND VPWR VPWR _18489_/X sky130_fd_sc_hd__or2_4
XFILLER_33_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21170__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13303__A _12255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20520_ _20520_/A VGND VGND VPWR VPWR _20520_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20451_ _20448_/X _20450_/X _24374_/Q _20407_/X VGND VGND VPWR VPWR _20451_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21520__A _21532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17126__B1 _15784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20382_ _20381_/X VGND VGND VPWR VPWR _20382_/Y sky130_fd_sc_hd__inv_2
X_23170_ _24065_/CLK _23170_/D VGND VGND VPWR VPWR _15259_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21473__A2 _21470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22670__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20136__A IRQ[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22121_ _22119_/X _22113_/X _23435_/Q _22120_/X VGND VGND VPWR VPWR _22121_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19925__A _22985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14134__A _14318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22052_ _22052_/A VGND VGND VPWR VPWR _22052_/X sky130_fd_sc_hd__buf_2
XFILLER_115_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22351__A _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21003_ _20511_/A _21002_/X _24063_/Q _20202_/X VGND VGND VPWR VPWR _24063_/D sky130_fd_sc_hd__o22a_4
XFILLER_114_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22973__A2 _16977_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13973__A _13643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12589__A _11740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22954_ _22954_/A VGND VGND VPWR VPWR HADDR[12] sky130_fd_sc_hd__inv_2
XFILLER_99_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21905_ _21884_/A VGND VGND VPWR VPWR _21905_/X sky130_fd_sc_hd__buf_2
X_22885_ _22885_/A VGND VGND VPWR VPWR HADDR[1] sky130_fd_sc_hd__inv_2
XFILLER_3_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21836_ _21812_/A VGND VGND VPWR VPWR _21836_/X sky130_fd_sc_hd__buf_2
XFILLER_110_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22489__B2 _22483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21767_ _21550_/X _21762_/X _15570_/B _21766_/X VGND VGND VPWR VPWR _23627_/D sky130_fd_sc_hd__o22a_4
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _24335_/Q _11520_/B VGND VGND VPWR VPWR _11521_/B sky130_fd_sc_hd__or2_4
X_23506_ _23986_/CLK _23506_/D VGND VGND VPWR VPWR _23506_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13213__A _12794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20718_ _20640_/X _20702_/X _20515_/X _20717_/Y VGND VGND VPWR VPWR _20718_/X sky130_fd_sc_hd__a211o_4
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21698_ _21705_/A VGND VGND VPWR VPWR _21698_/X sky130_fd_sc_hd__buf_2
XANTENNA__22526__A _22518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19106__A1 _18934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21430__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23437_ _23122_/CLK _23437_/D VGND VGND VPWR VPWR _15864_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20649_ _20754_/B VGND VGND VPWR VPWR _20822_/B sky130_fd_sc_hd__buf_2
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19657__A2 _19872_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14170_ _14617_/A _14170_/B _14169_/X VGND VGND VPWR VPWR _14170_/X sky130_fd_sc_hd__and3_4
XANTENNA__21464__A2 _21463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23368_ _23368_/CLK _23368_/D VGND VGND VPWR VPWR _13664_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22661__B2 _22626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13121_ _13096_/A _13119_/X _13121_/C VGND VGND VPWR VPWR _13121_/X sky130_fd_sc_hd__and3_4
XANTENNA__11668__A _13991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20672__B1 _15829_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22319_ _15539_/B VGND VGND VPWR VPWR _23307_/D sky130_fd_sc_hd__buf_2
XFILLER_3_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19835__A _19877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23299_ _23494_/CLK _23299_/D VGND VGND VPWR VPWR _14742_/B sky130_fd_sc_hd__dfxtp_4
X_13052_ _12496_/A _13122_/B VGND VGND VPWR VPWR _13054_/B sky130_fd_sc_hd__or2_4
XFILLER_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24324__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12003_ _11996_/A _11813_/B VGND VGND VPWR VPWR _12005_/B sky130_fd_sc_hd__or2_4
XFILLER_105_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13883__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17860_ _17860_/A VGND VGND VPWR VPWR _17861_/A sky130_fd_sc_hd__buf_2
XANTENNA__20975__A1 _22824_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14698__B _14698_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16811_ _16677_/A _16795_/X _16811_/C VGND VGND VPWR VPWR _16811_/X sky130_fd_sc_hd__or3_4
XFILLER_93_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17791_ _17101_/X VGND VGND VPWR VPWR _17792_/A sky130_fd_sc_hd__buf_2
XANTENNA__12499__A _12211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19530_ _19419_/A VGND VGND VPWR VPWR _19531_/A sky130_fd_sc_hd__buf_2
X_13954_ _12472_/A _14027_/B VGND VGND VPWR VPWR _13955_/C sky130_fd_sc_hd__or2_4
X_16742_ _11992_/X _16719_/X _16726_/X _16733_/X _16741_/X VGND VGND VPWR VPWR _16742_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_6_43_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12905_ _12905_/A _23411_/Q VGND VGND VPWR VPWR _12905_/X sky130_fd_sc_hd__or2_4
XFILLER_4_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16673_ _16670_/A _23644_/Q VGND VGND VPWR VPWR _16674_/C sky130_fd_sc_hd__or2_4
X_19461_ _24154_/Q _19459_/X HRDATA[28] _19460_/X VGND VGND VPWR VPWR _19461_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21605__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13885_ _13901_/A _13885_/B _13885_/C VGND VGND VPWR VPWR _13886_/C sky130_fd_sc_hd__and3_4
XFILLER_28_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18412_ _18381_/X _18411_/X _24462_/Q _18381_/X VGND VGND VPWR VPWR _24462_/D sky130_fd_sc_hd__a2bb2o_4
X_12836_ _12829_/A _12836_/B VGND VGND VPWR VPWR _12837_/C sky130_fd_sc_hd__or2_4
X_15624_ _15601_/A _23371_/Q VGND VGND VPWR VPWR _15624_/X sky130_fd_sc_hd__or2_4
X_19392_ _19385_/A VGND VGND VPWR VPWR _19392_/X sky130_fd_sc_hd__buf_2
XFILLER_62_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12946__B _23443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19345__B2 _20792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15555_ _15536_/A _23595_/Q VGND VGND VPWR VPWR _15555_/X sky130_fd_sc_hd__or2_4
X_18343_ _17694_/A VGND VGND VPWR VPWR _18383_/A sky130_fd_sc_hd__buf_2
XFILLER_37_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12767_ _12808_/A _12767_/B VGND VGND VPWR VPWR _12769_/B sky130_fd_sc_hd__or2_4
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21152__B2 _21151_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14533_/A _14506_/B VGND VGND VPWR VPWR _14506_/X sky130_fd_sc_hd__or2_4
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _11717_/X _23518_/Q VGND VGND VPWR VPWR _11718_/X sky130_fd_sc_hd__or2_4
X_18274_ _18274_/A _17495_/A _18274_/C VGND VGND VPWR VPWR _18274_/X sky130_fd_sc_hd__or3_4
X_15486_ _15486_/A _23884_/Q VGND VGND VPWR VPWR _15486_/X sky130_fd_sc_hd__or2_4
X_12698_ _12710_/A VGND VGND VPWR VPWR _15689_/A sky130_fd_sc_hd__buf_2
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14437_ _14464_/A _14435_/X _14436_/X VGND VGND VPWR VPWR _14437_/X sky130_fd_sc_hd__and3_4
X_17225_ _17222_/X _17826_/A _17224_/X VGND VGND VPWR VPWR _17225_/X sky130_fd_sc_hd__o21a_4
XFILLER_52_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11649_ _11648_/X VGND VGND VPWR VPWR _12965_/A sky130_fd_sc_hd__buf_2
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17156_ _12430_/X VGND VGND VPWR VPWR _17156_/Y sky130_fd_sc_hd__inv_2
X_14368_ _15586_/A _14292_/B VGND VGND VPWR VPWR _14368_/X sky130_fd_sc_hd__or2_4
XANTENNA__22652__B2 _22647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16107_ _16107_/A _23671_/Q VGND VGND VPWR VPWR _16109_/B sky130_fd_sc_hd__or2_4
X_13319_ _13283_/X _23952_/Q VGND VGND VPWR VPWR _13319_/X sky130_fd_sc_hd__or2_4
XANTENNA__11578__A _16893_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17087_ _18240_/A VGND VGND VPWR VPWR _18180_/A sky130_fd_sc_hd__buf_2
XANTENNA__19745__A _19429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14299_ _12269_/A _14298_/X VGND VGND VPWR VPWR _14299_/X sky130_fd_sc_hd__and2_4
XFILLER_6_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16038_ _16050_/A _23992_/Q VGND VGND VPWR VPWR _16038_/X sky130_fd_sc_hd__or2_4
XFILLER_118_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21207__A2 _21204_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15992__B _15992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_125_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR _23472_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18084__A1 _17989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17989_ _18216_/A VGND VGND VPWR VPWR _17989_/X sky130_fd_sc_hd__buf_2
XFILLER_22_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19728_ _19570_/A _19597_/A _19645_/A _19522_/X VGND VGND VPWR VPWR _19818_/A sky130_fd_sc_hd__or4_4
XANTENNA__19480__A _19742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12202__A _12202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20718__A1 _20640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23730__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21515__A _21515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19659_ _19659_/A _19573_/A VGND VGND VPWR VPWR _19718_/B sky130_fd_sc_hd__or2_4
XFILLER_77_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17712__B _17393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18096__A _16999_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21391__A1 _21282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16609__A _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21391__B2 _21387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15513__A _13087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22670_ _22664_/Y _22669_/X _21789_/A _22669_/X VGND VGND VPWR VPWR _22670_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16328__B _16267_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21621_ _21558_/X _21619_/X _13703_/B _21616_/X VGND VGND VPWR VPWR _21621_/X sky130_fd_sc_hd__o22a_4
XFILLER_34_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21143__B2 _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13033__A _12917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24340_ _23358_/CLK _18993_/X HRESETn VGND VGND VPWR VPWR _24340_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__17898__A1 _17766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21552_ _21550_/X _21544_/X _15530_/B _21551_/X VGND VGND VPWR VPWR _23755_/D sky130_fd_sc_hd__o22a_4
XFILLER_90_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21694__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20503_ _18222_/X _20447_/X _20492_/X _20502_/Y VGND VGND VPWR VPWR _20503_/X sky130_fd_sc_hd__a211o_4
X_24271_ _24092_/CLK _24271_/D HRESETn VGND VGND VPWR VPWR _19220_/A sky130_fd_sc_hd__dfrtp_4
X_21483_ _21268_/X _21477_/X _23786_/Q _21481_/X VGND VGND VPWR VPWR _21483_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12872__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23110__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16344__A _16365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23222_ _23313_/CLK _22482_/X VGND VGND VPWR VPWR _12323_/B sky130_fd_sc_hd__dfxtp_4
X_20434_ _20291_/X _20433_/X VGND VGND VPWR VPWR _20434_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21739__A2_N _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21446__A2 _21419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23153_ _23889_/CLK _23153_/D VGND VGND VPWR VPWR _13165_/B sky130_fd_sc_hd__dfxtp_4
X_20365_ _20321_/X _20364_/X _24314_/Q _20330_/X VGND VGND VPWR VPWR _20365_/X sky130_fd_sc_hd__o22a_4
X_22104_ _22103_/X _22101_/X _13091_/B _22096_/X VGND VGND VPWR VPWR _23442_/D sky130_fd_sc_hd__o22a_4
X_20296_ _20296_/A _20519_/B VGND VGND VPWR VPWR _20296_/Y sky130_fd_sc_hd__nand2_4
X_23084_ _23698_/CLK _22696_/X VGND VGND VPWR VPWR _23084_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14799__A _14050_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22081__A _20355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22035_ _22035_/A VGND VGND VPWR VPWR _22035_/X sky130_fd_sc_hd__buf_2
XFILLER_118_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17175__A _13274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22159__B1 _23421_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17903__A _18443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23986_ _23986_/CLK _21135_/X VGND VGND VPWR VPWR _23986_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12112__A _12112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21906__B1 _14293_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22937_ _22967_/A VGND VGND VPWR VPWR _22937_/X sky130_fd_sc_hd__buf_2
XFILLER_99_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21382__B2 _21380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15423__A _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13670_ _13670_/A _13670_/B _13669_/X VGND VGND VPWR VPWR _13674_/B sky130_fd_sc_hd__and3_4
X_22868_ _16444_/Y _22863_/X _22853_/X _22867_/X VGND VGND VPWR VPWR _22869_/B sky130_fd_sc_hd__o22a_4
XFILLER_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12621_ _12605_/A VGND VGND VPWR VPWR _15512_/A sky130_fd_sc_hd__buf_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21819_ _21249_/A VGND VGND VPWR VPWR _21819_/X sky130_fd_sc_hd__buf_2
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21134__A1 _20537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22799_ _17383_/Y _22794_/X _22796_/X _22798_/X VGND VGND VPWR VPWR _22800_/B sky130_fd_sc_hd__o22a_4
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18734__A _18713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14039__A _14039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21134__B2 _21130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15340_ _15333_/A _15267_/B VGND VGND VPWR VPWR _15341_/C sky130_fd_sc_hd__or2_4
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12552_ _13014_/A _12550_/X _12552_/C VGND VGND VPWR VPWR _12556_/B sky130_fd_sc_hd__and3_4
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _11503_/A VGND VGND VPWR VPWR _11505_/A sky130_fd_sc_hd__inv_2
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15271_ _14734_/A _15269_/X _15271_/C VGND VGND VPWR VPWR _15271_/X sky130_fd_sc_hd__and3_4
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _13953_/A VGND VGND VPWR VPWR _13643_/A sky130_fd_sc_hd__buf_2
X_24469_ _23522_/CLK _24469_/D HRESETn VGND VGND VPWR VPWR _24469_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16254__A _16147_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17010_ _17010_/A VGND VGND VPWR VPWR _17010_/X sky130_fd_sc_hd__buf_2
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ _11766_/A _14212_/X _14221_/X VGND VGND VPWR VPWR _14222_/X sky130_fd_sc_hd__and3_4
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22634__A1 _22410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22634__B2 _22633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14153_ _14117_/A _14149_/X _14153_/C VGND VGND VPWR VPWR _14153_/X sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_5_27_0_HCLK_A clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13104_ _13104_/A _13104_/B VGND VGND VPWR VPWR _13106_/B sky130_fd_sc_hd__or2_4
XFILLER_98_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14084_ _14089_/A _23721_/Q VGND VGND VPWR VPWR _14085_/C sky130_fd_sc_hd__or2_4
X_18961_ _18961_/A VGND VGND VPWR VPWR _18961_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11548__D _20071_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13035_ _12915_/A _13111_/B VGND VGND VPWR VPWR _13035_/X sky130_fd_sc_hd__or2_4
X_17912_ _17817_/X VGND VGND VPWR VPWR _17912_/X sky130_fd_sc_hd__buf_2
XFILLER_79_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18892_ _18892_/A VGND VGND VPWR VPWR _18892_/X sky130_fd_sc_hd__buf_2
XANTENNA__20948__A1 _20403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20948__B2 _20497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20223__B HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17843_ _17825_/X _17841_/X _17806_/X _17842_/X VGND VGND VPWR VPWR _17843_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_39_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15317__B _15255_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13118__A _13118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17774_ _17002_/A _17001_/C _16991_/B VGND VGND VPWR VPWR _23046_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__12022__A _12022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14986_ _11652_/X _14986_/B _14986_/C VGND VGND VPWR VPWR _14986_/X sky130_fd_sc_hd__and3_4
XFILLER_82_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19513_ _19523_/B VGND VGND VPWR VPWR _19829_/A sky130_fd_sc_hd__buf_2
XANTENNA__24109__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16725_ _12044_/X _16725_/B _16725_/C VGND VGND VPWR VPWR _16726_/C sky130_fd_sc_hd__and3_4
X_13937_ _13611_/A _13934_/X _13937_/C VGND VGND VPWR VPWR _13937_/X sky130_fd_sc_hd__and3_4
XANTENNA__12957__A _12957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11861__A _12458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19444_ _19839_/A VGND VGND VPWR VPWR _19445_/A sky130_fd_sc_hd__buf_2
X_13868_ _13895_/A _23559_/Q VGND VGND VPWR VPWR _13869_/C sky130_fd_sc_hd__or2_4
X_16656_ _16621_/A _16654_/X _16656_/C VGND VGND VPWR VPWR _16660_/B sky130_fd_sc_hd__and3_4
XFILLER_56_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12819_ _12803_/A _12819_/B VGND VGND VPWR VPWR _12820_/C sky130_fd_sc_hd__or2_4
X_15607_ _15607_/A _15607_/B _15607_/C VGND VGND VPWR VPWR _15611_/B sky130_fd_sc_hd__and3_4
XFILLER_72_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19375_ _19374_/X _18098_/X _19374_/X _24215_/Q VGND VGND VPWR VPWR _19375_/X sky130_fd_sc_hd__a2bb2o_4
X_13799_ _13799_/A _23559_/Q VGND VGND VPWR VPWR _13800_/C sky130_fd_sc_hd__or2_4
X_16587_ _12024_/A _23804_/Q VGND VGND VPWR VPWR _16588_/C sky130_fd_sc_hd__or2_4
XFILLER_17_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23133__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21125__B2 _21123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18326_ _17962_/X _17236_/X _17964_/X VGND VGND VPWR VPWR _18326_/Y sky130_fd_sc_hd__o21ai_4
X_15538_ _15571_/A _15536_/X _15537_/X VGND VGND VPWR VPWR _15538_/X sky130_fd_sc_hd__and3_4
XANTENNA__14891__B _23584_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13788__A _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15469_ _13770_/A _15461_/X _15469_/C VGND VGND VPWR VPWR _15469_/X sky130_fd_sc_hd__and3_4
X_18257_ _18171_/X _18238_/X _18202_/X _18256_/X VGND VGND VPWR VPWR _18257_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12692__A _12688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17208_ _17151_/X _17204_/X _17160_/X _17207_/X VGND VGND VPWR VPWR _17208_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_102_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21428__A2 _21426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18188_ _18107_/X _18185_/Y _17240_/X _18187_/X VGND VGND VPWR VPWR _18188_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22625__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17139_ _14988_/X _17137_/X _17007_/X _17138_/X VGND VGND VPWR VPWR _17139_/X sky130_fd_sc_hd__o22a_4
X_20150_ _20145_/Y _20146_/Y _11536_/X _20149_/Y VGND VGND VPWR VPWR _20150_/X sky130_fd_sc_hd__o22a_4
XFILLER_48_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20414__A _20414_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20081_ _19411_/X _20080_/X _19411_/X _16960_/A VGND VGND VPWR VPWR _20081_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15508__A _13735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14412__A _15611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21600__A2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24370__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14131__B _23945_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23840_ _23840_/CLK _23840_/D VGND VGND VPWR VPWR _23840_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13028__A _12518_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23771_ _23707_/CLK _23771_/D VGND VGND VPWR VPWR _23771_/Q sky130_fd_sc_hd__dfxtp_4
X_20983_ _20872_/X _20982_/X _14903_/B _20202_/X VGND VGND VPWR VPWR _24064_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12867__A _12528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20167__A2 IRQ[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16339__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21364__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11771__A _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22722_ _22898_/A _19303_/X _23064_/B _22721_/Y VGND VGND VPWR VPWR _22722_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12586__B _12586_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22653_ _22444_/X _22650_/X _13814_/B _22647_/X VGND VGND VPWR VPWR _23111_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18554__A _18381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21604_ _21529_/X _21598_/X _12768_/B _21602_/X VGND VGND VPWR VPWR _23732_/D sky130_fd_sc_hd__o22a_4
XFILLER_70_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21667__A2 _21662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22584_ _22410_/X _22579_/X _12620_/B _22583_/X VGND VGND VPWR VPWR _22584_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22076__A _22125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24323_ _24330_/CLK _19091_/X HRESETn VGND VGND VPWR VPWR _24323_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__23626__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13698__A _13697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21535_ _21534_/X _21532_/X _13075_/B _21527_/X VGND VGND VPWR VPWR _21535_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24254_ _24250_/CLK _19310_/X HRESETn VGND VGND VPWR VPWR _20210_/A sky130_fd_sc_hd__dfrtp_4
X_21466_ _21239_/X _21463_/X _12329_/B _21460_/X VGND VGND VPWR VPWR _23798_/D sky130_fd_sc_hd__o22a_4
XFILLER_33_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_7_0_HCLK clkbuf_6_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23205_ _23557_/CLK _22506_/X VGND VGND VPWR VPWR _14479_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_68_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20417_ _24216_/Q _20398_/X _20416_/Y VGND VGND VPWR VPWR _20418_/A sky130_fd_sc_hd__o21a_4
X_24185_ _24162_/CLK _19613_/X HRESETn VGND VGND VPWR VPWR _17533_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22092__A2 _22089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21397_ _23838_/Q VGND VGND VPWR VPWR _21397_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23776__CLK _23840_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23136_ _23233_/CLK _23136_/D VGND VGND VPWR VPWR _14882_/B sky130_fd_sc_hd__dfxtp_4
X_20348_ _20321_/X _20347_/X _24315_/Q _20330_/X VGND VGND VPWR VPWR _20348_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15418__A _13654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23067_ VGND VGND VPWR VPWR _23067_/HI HSIZE[2] sky130_fd_sc_hd__conb_1
XFILLER_66_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20279_ _20279_/A VGND VGND VPWR VPWR _20511_/A sky130_fd_sc_hd__buf_2
XANTENNA__14322__A _14322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19796__A1 _19706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18599__A2 _18577_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22018_ _22017_/X VGND VGND VPWR VPWR _22052_/A sky130_fd_sc_hd__buf_2
XFILLER_49_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14840_ _14816_/A _14836_/X _14839_/X VGND VGND VPWR VPWR _14840_/X sky130_fd_sc_hd__or3_4
XFILLER_79_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14771_ _13800_/A _14769_/X _14771_/C VGND VGND VPWR VPWR _14771_/X sky130_fd_sc_hd__and3_4
XFILLER_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11983_ _11983_/A _23934_/Q VGND VGND VPWR VPWR _11985_/B sky130_fd_sc_hd__or2_4
X_23969_ _24032_/CLK _21158_/X VGND VGND VPWR VPWR _15210_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12777__A _13087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11681__A _11680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13722_ _13770_/A _13705_/X _13721_/X VGND VGND VPWR VPWR _13722_/X sky130_fd_sc_hd__and3_4
X_16510_ _16363_/X _16506_/X _16510_/C VGND VGND VPWR VPWR _16511_/C sky130_fd_sc_hd__or3_4
X_17490_ _17489_/X VGND VGND VPWR VPWR _17490_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13653_ _13796_/A _13651_/X _13652_/X VGND VGND VPWR VPWR _13658_/B sky130_fd_sc_hd__and3_4
X_16441_ _11851_/X _16440_/X VGND VGND VPWR VPWR _16441_/X sky130_fd_sc_hd__and2_4
XANTENNA__18464__A _18418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14992__A _14992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21107__B2 _21072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12604_ _12604_/A _24021_/Q VGND VGND VPWR VPWR _12604_/X sky130_fd_sc_hd__or2_4
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16372_ _11800_/X _16372_/B _16372_/C VGND VGND VPWR VPWR _16373_/C sky130_fd_sc_hd__or3_4
X_19160_ _19129_/A _19129_/B _19159_/Y VGND VGND VPWR VPWR _24308_/D sky130_fd_sc_hd__o21a_4
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13584_ _16899_/A _13583_/Y VGND VGND VPWR VPWR _15927_/A sky130_fd_sc_hd__or2_4
XANTENNA__21658__A2 _21655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15323_ _15314_/A _15260_/B VGND VGND VPWR VPWR _15324_/C sky130_fd_sc_hd__or2_4
X_18111_ _17910_/X _17925_/X _17252_/X VGND VGND VPWR VPWR _18111_/X sky130_fd_sc_hd__o21a_4
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20866__B1 _20865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12535_ _12904_/A _12647_/B VGND VGND VPWR VPWR _12535_/X sky130_fd_sc_hd__or2_4
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19091_ _19087_/X _19090_/X _19087_/X _24323_/Q VGND VGND VPWR VPWR _19091_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13348__A1 _11980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20218__B HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15254_ _14098_/A _15254_/B _15254_/C VGND VGND VPWR VPWR _15254_/X sky130_fd_sc_hd__and3_4
X_18042_ _18040_/X _18041_/X _17868_/X VGND VGND VPWR VPWR _18042_/Y sky130_fd_sc_hd__o21ai_4
X_12466_ _12917_/A VGND VGND VPWR VPWR _12466_/X sky130_fd_sc_hd__buf_2
XANTENNA__22714__A _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14205_ _14205_/A _23561_/Q VGND VGND VPWR VPWR _14205_/X sky130_fd_sc_hd__or2_4
X_15185_ _11839_/X _11615_/X _15154_/X _11592_/X _15184_/X VGND VGND VPWR VPWR _15185_/X
+ sky130_fd_sc_hd__a32o_4
X_12397_ _12419_/A _24054_/Q VGND VGND VPWR VPWR _12398_/C sky130_fd_sc_hd__or2_4
X_14136_ _14136_/A _14136_/B _14136_/C VGND VGND VPWR VPWR _14136_/X sky130_fd_sc_hd__or3_4
X_19993_ _19992_/X VGND VGND VPWR VPWR _19993_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21830__A2 _21829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14067_ _14026_/A VGND VGND VPWR VPWR _14068_/A sky130_fd_sc_hd__buf_2
X_18944_ _24380_/Q VGND VGND VPWR VPWR _18944_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14232__A _14246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13018_ _13041_/A _13014_/X _13018_/C VGND VGND VPWR VPWR _13018_/X sky130_fd_sc_hd__or3_4
XFILLER_67_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18875_ _18891_/A VGND VGND VPWR VPWR _18875_/X sky130_fd_sc_hd__buf_2
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21594__B2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17826_ _17826_/A VGND VGND VPWR VPWR _17826_/X sky130_fd_sc_hd__buf_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21065__A _21072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17757_ _17757_/A VGND VGND VPWR VPWR _17758_/B sky130_fd_sc_hd__inv_2
X_14969_ _14243_/A _14969_/B _14968_/X VGND VGND VPWR VPWR _14985_/B sky130_fd_sc_hd__and3_4
XANTENNA__12687__A _12286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20149__A2 IRQ[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_13_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21346__B2 _21301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15063__A _15063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16708_ _11921_/X _16708_/B VGND VGND VPWR VPWR _16709_/C sky130_fd_sc_hd__or2_4
XFILLER_78_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24081__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21897__A2 _21894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17688_ _24132_/Q _17688_/B VGND VGND VPWR VPWR _17755_/B sky130_fd_sc_hd__and2_4
XFILLER_1_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19427_ HRDATA[0] _19545_/A _19426_/X VGND VGND VPWR VPWR _19428_/A sky130_fd_sc_hd__a21o_4
XANTENNA__15998__A _15948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16639_ _16621_/A _16637_/X _16639_/C VGND VGND VPWR VPWR _16639_/X sky130_fd_sc_hd__and3_4
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19358_ _19355_/X _18723_/X _19355_/X _24224_/Q VGND VGND VPWR VPWR _24224_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21649__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18309_ _18294_/X _18299_/Y _18305_/X _18307_/X _18308_/Y VGND VGND VPWR VPWR _18309_/X
+ sky130_fd_sc_hd__a32o_4
X_19289_ _19209_/B VGND VGND VPWR VPWR _19289_/Y sky130_fd_sc_hd__inv_2
X_21320_ _21246_/X _21319_/X _23891_/Q _21316_/X VGND VGND VPWR VPWR _21320_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13311__A _15696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21251_ _20574_/A VGND VGND VPWR VPWR _21251_/X sky130_fd_sc_hd__buf_2
XFILLER_11_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19475__B1 HRDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16622__A _16622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20085__A1 _19884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20202_ _20488_/A VGND VGND VPWR VPWR _20202_/X sky130_fd_sc_hd__buf_2
X_21182_ _20509_/X _21176_/X _23956_/Q _21180_/X VGND VGND VPWR VPWR _21182_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20144__A IRQ[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11766__A _11766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20133_ _18708_/X VGND VGND VPWR VPWR _20133_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15238__A _14345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19933__A _19933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14142__A _14113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20064_ _20042_/X _18533_/A _20048_/X _20063_/X VGND VGND VPWR VPWR _20065_/A sky130_fd_sc_hd__o22a_4
XFILLER_28_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18450__A1 _18216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17453__A _12841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23823_ _23859_/CLK _21425_/X VGND VGND VPWR VPWR _23823_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12597__A _14177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23754_ _23978_/CLK _21554_/X VGND VGND VPWR VPWR _23754_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20966_ _20966_/A VGND VGND VPWR VPWR _20966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21888__A2 _21887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22705_ _20838_/A _22700_/X _14327_/B _22704_/X VGND VGND VPWR VPWR _23078_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19950__A1 _17989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18753__A2 _18752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23685_ _23845_/CLK _23685_/D VGND VGND VPWR VPWR _14486_/B sky130_fd_sc_hd__dfxtp_4
X_20897_ _20223_/A _20895_/X _20896_/X HRDATA[12] _20846_/X VGND VGND VPWR VPWR _20897_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_13_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15701__A _12849_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22636_ _22636_/A VGND VGND VPWR VPWR _22636_/X sky130_fd_sc_hd__buf_2
XANTENNA__16516__B _16513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20848__B1 HRDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22567_ _22600_/A VGND VGND VPWR VPWR _22583_/A sky130_fd_sc_hd__inv_2
Xclkbuf_7_33_0_HCLK clkbuf_7_33_0_HCLK/A VGND VGND VPWR VPWR _23494_/CLK sky130_fd_sc_hd__clkbuf_1
X_12320_ _12320_/A VGND VGND VPWR VPWR _12435_/A sky130_fd_sc_hd__buf_2
X_24306_ _24305_/CLK _24306_/D HRESETn VGND VGND VPWR VPWR _24306_/Q sky130_fd_sc_hd__dfrtp_4
X_21518_ _21517_/X _21508_/X _16249_/B _21515_/X VGND VGND VPWR VPWR _23769_/D sky130_fd_sc_hd__o22a_4
XFILLER_103_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_96_0_HCLK clkbuf_6_48_0_HCLK/X VGND VGND VPWR VPWR _23487_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22498_ _22434_/X _22493_/X _23211_/Q _22497_/X VGND VGND VPWR VPWR _22498_/X sky130_fd_sc_hd__o22a_4
X_12251_ _13985_/A VGND VGND VPWR VPWR _12252_/A sky130_fd_sc_hd__buf_2
X_24237_ _24239_/CLK _24237_/D HRESETn VGND VGND VPWR VPWR _24237_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21449_ _21784_/A _21348_/B _21348_/C _21734_/B VGND VGND VPWR VPWR _21449_/X sky130_fd_sc_hd__or4_4
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22065__A2 _22031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19466__B1 HRDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16532__A _12011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12182_ _16677_/A _12166_/X _12182_/C VGND VGND VPWR VPWR _12183_/C sky130_fd_sc_hd__or3_4
X_24168_ _23584_/CLK _19833_/Y HRESETn VGND VGND VPWR VPWR _21296_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24171__D _24171_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16251__B _24025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23119_ _23827_/CLK _23119_/D VGND VGND VPWR VPWR _13547_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15148__A _14998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_16990_ _17769_/A _17000_/A VGND VGND VPWR VPWR _16991_/B sky130_fd_sc_hd__or2_4
X_24099_ _24321_/CLK _24099_/D HRESETn VGND VGND VPWR VPWR _24099_/Q sky130_fd_sc_hd__dfrtp_4
X_15941_ _15976_/A _15941_/B _15941_/C VGND VGND VPWR VPWR _15942_/C sky130_fd_sc_hd__and3_4
XFILLER_110_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13891__A _13879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18660_ _18424_/X _17965_/Y _17854_/X _18659_/Y VGND VGND VPWR VPWR _18660_/X sky130_fd_sc_hd__a211o_4
XFILLER_27_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15872_ _13500_/X _15870_/X _15871_/X VGND VGND VPWR VPWR _15873_/C sky130_fd_sc_hd__and3_4
XFILLER_77_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17611_ _17330_/A VGND VGND VPWR VPWR _17611_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14823_ _14811_/A _14759_/B VGND VGND VPWR VPWR _14824_/C sky130_fd_sc_hd__or2_4
X_18591_ _18591_/A VGND VGND VPWR VPWR _18591_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21328__B2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17542_ _16302_/X VGND VGND VPWR VPWR _17542_/Y sky130_fd_sc_hd__inv_2
X_11966_ _11916_/X VGND VGND VPWR VPWR _11966_/X sky130_fd_sc_hd__buf_2
X_14754_ _15450_/A _14731_/X _14738_/X _14745_/X _14753_/X VGND VGND VPWR VPWR _14754_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_79_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12300__A _12706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13705_ _13754_/A _13699_/X _13705_/C VGND VGND VPWR VPWR _13705_/X sky130_fd_sc_hd__or3_4
X_14685_ _15589_/A _14681_/X _14684_/X VGND VGND VPWR VPWR _14685_/X sky130_fd_sc_hd__or3_4
X_17473_ _12676_/X _17527_/B VGND VGND VPWR VPWR _17473_/X sky130_fd_sc_hd__and2_4
X_11897_ _12852_/A VGND VGND VPWR VPWR _12444_/A sky130_fd_sc_hd__buf_2
XFILLER_32_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16707__A _11888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19212_ _19212_/A _19212_/B VGND VGND VPWR VPWR _19213_/B sky130_fd_sc_hd__and2_4
X_13636_ _13636_/A _13636_/B VGND VGND VPWR VPWR _13637_/C sky130_fd_sc_hd__or2_4
X_16424_ _16397_/X _16424_/B VGND VGND VPWR VPWR _16424_/X sky130_fd_sc_hd__or2_4
XFILLER_38_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15611__A _15611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22828__A1 _15051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20229__A _20229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19143_ _19137_/X VGND VGND VPWR VPWR _19143_/Y sky130_fd_sc_hd__inv_2
X_13567_ _13500_/X _13565_/X _13567_/C VGND VGND VPWR VPWR _13571_/B sky130_fd_sc_hd__and3_4
X_16355_ _11681_/X VGND VGND VPWR VPWR _16355_/X sky130_fd_sc_hd__buf_2
XFILLER_12_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14227__A _14195_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12518_ _12518_/A VGND VGND VPWR VPWR _12518_/X sky130_fd_sc_hd__buf_2
X_15306_ _13925_/A _15306_/B VGND VGND VPWR VPWR _15308_/B sky130_fd_sc_hd__or2_4
X_16286_ _16286_/A _23481_/Q VGND VGND VPWR VPWR _16286_/X sky130_fd_sc_hd__or2_4
X_19074_ _18935_/X VGND VGND VPWR VPWR _19074_/X sky130_fd_sc_hd__buf_2
XFILLER_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13498_ _15884_/A _23503_/Q VGND VGND VPWR VPWR _13498_/X sky130_fd_sc_hd__or2_4
XFILLER_69_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22444__A _22129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18025_ _18025_/A VGND VGND VPWR VPWR _18295_/A sky130_fd_sc_hd__buf_2
XFILLER_51_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12449_ _12449_/A VGND VGND VPWR VPWR _12450_/A sky130_fd_sc_hd__buf_2
X_15237_ _14210_/A _15180_/B VGND VGND VPWR VPWR _15237_/X sky130_fd_sc_hd__or2_4
XANTENNA__12970__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20067__B2 _19929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21264__B1 _23916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15168_ _14145_/A _15164_/X _15167_/X VGND VGND VPWR VPWR _15168_/X sky130_fd_sc_hd__or3_4
XANTENNA__21803__A2 _21793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13785__B _23751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14119_ _12301_/A VGND VGND VPWR VPWR _14119_/X sky130_fd_sc_hd__buf_2
X_15099_ _15107_/A _15099_/B _15099_/C VGND VGND VPWR VPWR _15100_/C sky130_fd_sc_hd__and3_4
X_19976_ _20000_/A VGND VGND VPWR VPWR _19976_/X sky130_fd_sc_hd__buf_2
XANTENNA__24447__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18927_ _18927_/A _18926_/X VGND VGND VPWR VPWR _18927_/X sky130_fd_sc_hd__and2_4
XFILLER_68_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19472__B _19754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18858_ _17297_/X _18855_/X _24388_/Q _18856_/X VGND VGND VPWR VPWR _24388_/D sky130_fd_sc_hd__o22a_4
X_17809_ _17802_/X _17134_/X _17808_/X _17142_/X VGND VGND VPWR VPWR _17809_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15505__B _23852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18789_ _18789_/A VGND VGND VPWR VPWR _18789_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20820_ _20750_/X _20819_/X _24071_/Q _20724_/X VGND VGND VPWR VPWR _20820_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22619__A _22626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20751_ _20512_/A VGND VGND VPWR VPWR _20751_/X sky130_fd_sc_hd__buf_2
XANTENNA__17720__B _17290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17943__B1 _17878_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23470_ _23692_/CLK _23470_/D VGND VGND VPWR VPWR _15769_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22819__A1 _15910_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20682_ _20258_/X VGND VGND VPWR VPWR _20682_/X sky130_fd_sc_hd__buf_2
XFILLER_50_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22421_ _22420_/X _22416_/X _13137_/B _22411_/X VGND VGND VPWR VPWR _23249_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15240__B _15240_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22295__A2 _22293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19928__A _19927_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13041__A _13041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22352_ _22095_/X _22347_/X _12607_/B _22351_/X VGND VGND VPWR VPWR _22352_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22354__A _22354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21303_ _21295_/Y _21302_/X _21219_/X _21302_/X VGND VGND VPWR VPWR _21303_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13976__A _12202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22047__A2 _22045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22283_ _22269_/A VGND VGND VPWR VPWR _22283_/X sky130_fd_sc_hd__buf_2
XANTENNA__19448__B1 _18016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16352__A _11727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24022_ _23316_/CLK _21078_/X VGND VGND VPWR VPWR _12236_/B sky130_fd_sc_hd__dfxtp_4
X_21234_ _21804_/A VGND VGND VPWR VPWR _21234_/X sky130_fd_sc_hd__buf_2
XFILLER_2_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16071__B _15992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21165_ _21180_/A VGND VGND VPWR VPWR _21165_/X sky130_fd_sc_hd__buf_2
XFILLER_85_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22801__B _15120_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20116_ _11550_/X _20114_/X _20115_/Y VGND VGND VPWR VPWR _20116_/X sky130_fd_sc_hd__o21a_4
X_21096_ _21067_/A VGND VGND VPWR VPWR _21096_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20047_ _20047_/A VGND VGND VPWR VPWR _20047_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14600__A _14617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20230__A1 _18759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11820_ _11820_/A _11820_/B _11820_/C VGND VGND VPWR VPWR _11820_/X sky130_fd_sc_hd__and3_4
X_23806_ _23320_/CLK _23806_/D VGND VGND VPWR VPWR _23806_/Q sky130_fd_sc_hd__dfxtp_4
X_21998_ _21833_/X _21995_/X _15455_/B _21992_/X VGND VGND VPWR VPWR _23500_/D sky130_fd_sc_hd__o22a_4
XFILLER_42_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22529__A _22536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19923__A1 _19909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11748_/X _11749_/X _11750_/X VGND VGND VPWR VPWR _11751_/X sky130_fd_sc_hd__and3_4
X_23737_ _23770_/CLK _21597_/X VGND VGND VPWR VPWR _16245_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_82_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19923__B2 _19770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20949_ _20494_/A _20948_/X _11503_/A _20453_/A VGND VGND VPWR VPWR _20949_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20533__A2 _20421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21730__B2 _21687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15431__A _15431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _12885_/A _14470_/B VGND VGND VPWR VPWR _14470_/X sky130_fd_sc_hd__or2_4
XFILLER_92_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11681_/X VGND VGND VPWR VPWR _13415_/A sky130_fd_sc_hd__buf_2
X_23668_ _23316_/CLK _21704_/X VGND VGND VPWR VPWR _12799_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24166__D _19850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12774__B _12774_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13399_/A _13419_/X _13421_/C VGND VGND VPWR VPWR _13422_/C sky130_fd_sc_hd__and3_4
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22619_ _22626_/A VGND VGND VPWR VPWR _22619_/X sky130_fd_sc_hd__buf_2
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23599_ _23311_/CLK _21827_/X VGND VGND VPWR VPWR _23599_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14047__A _14847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18742__A _18728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16140_ _16140_/A _16140_/B _16139_/X VGND VGND VPWR VPWR _16144_/B sky130_fd_sc_hd__and3_4
X_13352_ _12802_/A VGND VGND VPWR VPWR _13352_/X sky130_fd_sc_hd__buf_2
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17162__A1 _14723_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12303_ _12459_/A VGND VGND VPWR VPWR _15558_/A sky130_fd_sc_hd__buf_2
X_16071_ _16071_/A _15992_/B VGND VGND VPWR VPWR _16071_/X sky130_fd_sc_hd__or2_4
XANTENNA__13886__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13283_ _13046_/A VGND VGND VPWR VPWR _13283_/X sky130_fd_sc_hd__buf_2
XANTENNA__16262__A _16095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15022_ _14588_/X _23583_/Q VGND VGND VPWR VPWR _15024_/B sky130_fd_sc_hd__or2_4
X_12234_ _12233_/X VGND VGND VPWR VPWR _12235_/A sky130_fd_sc_hd__buf_2
XANTENNA__17077__B _18203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19830_ _19830_/A VGND VGND VPWR VPWR _21582_/A sky130_fd_sc_hd__buf_2
X_12165_ _11685_/X _12161_/X _12164_/X VGND VGND VPWR VPWR _12166_/C sky130_fd_sc_hd__or3_4
X_19761_ HRDATA[17] VGND VGND VPWR VPWR _20576_/B sky130_fd_sc_hd__buf_2
X_12096_ _12096_/A _12096_/B _12096_/C VGND VGND VPWR VPWR _12096_/X sky130_fd_sc_hd__or3_4
X_16973_ _16973_/A _16973_/B VGND VGND VPWR VPWR _16974_/B sky130_fd_sc_hd__or2_4
XANTENNA__23494__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20512__A _20512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18189__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21549__B2 _21539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18712_ _18082_/A _17808_/X _18711_/X VGND VGND VPWR VPWR _18712_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_42_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17093__A _18656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15924_ _15923_/X VGND VGND VPWR VPWR _15924_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19692_ _19661_/B _19690_/X _19877_/A VGND VGND VPWR VPWR _19692_/X sky130_fd_sc_hd__a21o_4
XANTENNA__14510__A _13895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18643_ _17726_/X _18642_/A _22907_/B _18644_/A VGND VGND VPWR VPWR _18643_/X sky130_fd_sc_hd__o22a_4
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15855_ _13546_/X _15855_/B VGND VGND VPWR VPWR _15855_/X sky130_fd_sc_hd__or2_4
XFILLER_92_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14806_ _14845_/A _14806_/B VGND VGND VPWR VPWR _14806_/X sky130_fd_sc_hd__or2_4
X_18574_ _18554_/X _18573_/X _24455_/Q _18554_/X VGND VGND VPWR VPWR _24455_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15786_ _12849_/A _15784_/X _15785_/X VGND VGND VPWR VPWR _15786_/X sky130_fd_sc_hd__and3_4
XANTENNA__24449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12998_ _12850_/A _13064_/B VGND VGND VPWR VPWR _12998_/X sky130_fd_sc_hd__or2_4
XANTENNA__22439__A _20778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17525_ _17182_/Y _17525_/B VGND VGND VPWR VPWR _17525_/X sky130_fd_sc_hd__or2_4
XANTENNA__19914__B2 _20445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14737_ _14737_/A _14737_/B _14737_/C VGND VGND VPWR VPWR _14738_/C sky130_fd_sc_hd__and3_4
XFILLER_45_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11949_ _11983_/A VGND VGND VPWR VPWR _11996_/A sky130_fd_sc_hd__buf_2
XANTENNA__12965__A _12965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21721__B2 _21716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18193__A3 _18188_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17456_ _17455_/X VGND VGND VPWR VPWR _17456_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14668_ _14664_/X _14665_/X _14667_/X VGND VGND VPWR VPWR _14668_/X sky130_fd_sc_hd__and3_4
X_16407_ _16394_/X _16407_/B VGND VGND VPWR VPWR _16409_/B sky130_fd_sc_hd__or2_4
XFILLER_53_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13619_ _12883_/A VGND VGND VPWR VPWR _13620_/A sky130_fd_sc_hd__buf_2
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22277__A2 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17387_ _13920_/X _17388_/A VGND VGND VPWR VPWR _17387_/X sky130_fd_sc_hd__or2_4
X_14599_ _14151_/A _23556_/Q VGND VGND VPWR VPWR _14600_/C sky130_fd_sc_hd__or2_4
XFILLER_53_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19126_ _24305_/Q _19167_/A VGND VGND VPWR VPWR _19165_/A sky130_fd_sc_hd__and2_4
X_16338_ _11770_/X _16338_/B _16338_/C VGND VGND VPWR VPWR _16338_/X sky130_fd_sc_hd__and3_4
XANTENNA__17153__A1 _14429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19057_ _19027_/A VGND VGND VPWR VPWR _19057_/X sky130_fd_sc_hd__buf_2
XANTENNA__17268__A _17266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16269_ _11933_/X _16265_/X _16268_/X VGND VGND VPWR VPWR _16269_/X sky130_fd_sc_hd__or3_4
XANTENNA__16172__A _16203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18008_ _16925_/Y VGND VGND VPWR VPWR _18198_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22902__A _23051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12205__A _12496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20996__C1 _20995_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19959_ _18653_/X _19306_/Y _19934_/X _19958_/X VGND VGND VPWR VPWR _19960_/A sky130_fd_sc_hd__o22a_4
XFILLER_101_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15516__A _12392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22970_ _22982_/A _22968_/X _22970_/C VGND VGND VPWR VPWR _22970_/X sky130_fd_sc_hd__and3_4
XFILLER_60_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20212__A1 _16907_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21921_ _21920_/X VGND VGND VPWR VPWR _21921_/X sky130_fd_sc_hd__buf_2
XFILLER_56_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21960__A1 _21852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21960__B2 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18827__A _18834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13036__A _13009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21852_ _21282_/A VGND VGND VPWR VPWR _21852_/X sky130_fd_sc_hd__buf_2
XFILLER_42_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20803_ _24391_/Q _20556_/A VGND VGND VPWR VPWR _20803_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__19905__B2 _20650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21783_ _23614_/Q VGND VGND VPWR VPWR _21783_/Y sky130_fd_sc_hd__inv_2
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24119__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16347__A _16185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23522_ _23522_/CLK _23522_/D VGND VGND VPWR VPWR _15343_/B sky130_fd_sc_hd__dfxtp_4
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20734_ _24394_/Q _20623_/X _24426_/Q _20682_/X VGND VGND VPWR VPWR _20734_/X sky130_fd_sc_hd__o22a_4
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23453_ _23293_/CLK _23453_/D VGND VGND VPWR VPWR _12140_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_50_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20665_ _20665_/A VGND VGND VPWR VPWR _20665_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22268__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22404_ _22416_/A VGND VGND VPWR VPWR _22404_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23384_ _23383_/CLK _23384_/D VGND VGND VPWR VPWR _15984_/B sky130_fd_sc_hd__dfxtp_4
X_20596_ _24431_/Q VGND VGND VPWR VPWR _20596_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22084__A _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22335_ _22368_/A VGND VGND VPWR VPWR _22351_/A sky130_fd_sc_hd__inv_2
XANTENNA__17178__A _13772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16082__A _13442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21228__B1 _23931_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22266_ _22088_/X _22265_/X _23352_/Q _22262_/X VGND VGND VPWR VPWR _23352_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24005_ _23973_/CLK _21102_/X VGND VGND VPWR VPWR _14442_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21779__B2 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21217_ _21242_/A VGND VGND VPWR VPWR _21230_/A sky130_fd_sc_hd__buf_2
X_22197_ _22143_/X _22193_/X _15166_/B _22162_/A VGND VGND VPWR VPWR _23393_/D sky130_fd_sc_hd__o22a_4
XFILLER_78_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16810__A _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20451__A1 _20448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21148_ _20779_/X _21147_/X _23977_/Q _21144_/X VGND VGND VPWR VPWR _23977_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11954__A _11954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15426__A _15430_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13970_ _12509_/A _13970_/B VGND VGND VPWR VPWR _13971_/C sky130_fd_sc_hd__or2_4
X_21079_ _21079_/A VGND VGND VPWR VPWR _21079_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12921_ _13041_/A _12921_/B _12921_/C VGND VGND VPWR VPWR _12921_/X sky130_fd_sc_hd__or3_4
XFILLER_101_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21951__B2 _21949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15640_ _13845_/A _15570_/B VGND VGND VPWR VPWR _15641_/C sky130_fd_sc_hd__or2_4
XFILLER_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17641__A _17769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12852_ _12852_/A VGND VGND VPWR VPWR _12895_/A sky130_fd_sc_hd__buf_2
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11803_ _11803_/A _23902_/Q VGND VGND VPWR VPWR _11803_/X sky130_fd_sc_hd__or2_4
X_12783_ _15725_/A VGND VGND VPWR VPWR _12800_/A sky130_fd_sc_hd__buf_2
X_15571_ _15571_/A _15571_/B _15571_/C VGND VGND VPWR VPWR _15571_/X sky130_fd_sc_hd__and3_4
XFILLER_37_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12785__A _12813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21703__B2 _21702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17307_/Y _17308_/X _17309_/X VGND VGND VPWR VPWR _17310_/X sky130_fd_sc_hd__o21a_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15161__A _14136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11734_/A _23742_/Q VGND VGND VPWR VPWR _11734_/X sky130_fd_sc_hd__or2_4
X_14522_ _13747_/A _14517_/X _14521_/X VGND VGND VPWR VPWR _14522_/X sky130_fd_sc_hd__or3_4
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12995__A2 _12992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18290_ _18228_/X _18289_/X _24466_/Q _18228_/X VGND VGND VPWR VPWR _18290_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24347__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _18728_/B VGND VGND VPWR VPWR _17242_/A sky130_fd_sc_hd__buf_2
XFILLER_42_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _12957_/A VGND VGND VPWR VPWR _11665_/X sky130_fd_sc_hd__buf_2
X_14453_ _15392_/A _14453_/B VGND VGND VPWR VPWR _14455_/B sky130_fd_sc_hd__or2_4
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24292__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _13395_/X _13328_/B VGND VGND VPWR VPWR _13404_/X sky130_fd_sc_hd__or2_4
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _13844_/A VGND VGND VPWR VPWR _15633_/A sky130_fd_sc_hd__buf_2
X_17172_ _17171_/X VGND VGND VPWR VPWR _17172_/Y sky130_fd_sc_hd__inv_2
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ _11596_/A VGND VGND VPWR VPWR _11596_/X sky130_fd_sc_hd__buf_2
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16704__B _23931_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13335_ _12849_/A VGND VGND VPWR VPWR _13467_/A sky130_fd_sc_hd__buf_2
X_16123_ _11853_/X _16095_/X _16105_/X _16113_/X _16122_/X VGND VGND VPWR VPWR _16123_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18883__A1 _16514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20690__A1 _18453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13266_ _12367_/A _13266_/B _13265_/X VGND VGND VPWR VPWR _13266_/X sky130_fd_sc_hd__or3_4
X_16054_ _16047_/A _23832_/Q VGND VGND VPWR VPWR _16054_/X sky130_fd_sc_hd__or2_4
X_12217_ _12217_/A VGND VGND VPWR VPWR _13632_/A sky130_fd_sc_hd__buf_2
X_15005_ _15028_/A _15005_/B _15004_/X VGND VGND VPWR VPWR _15009_/B sky130_fd_sc_hd__and3_4
XFILLER_83_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18635__A1 _18500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13197_ _15707_/A _13257_/B VGND VGND VPWR VPWR _13197_/X sky130_fd_sc_hd__or2_4
XANTENNA__12025__A _12025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22431__A2 _22428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19832__B1 _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19813_ _19813_/A _19808_/X _19812_/X VGND VGND VPWR VPWR _19813_/X sky130_fd_sc_hd__and3_4
X_12148_ _11730_/X _12146_/X _12147_/X VGND VGND VPWR VPWR _12148_/X sky130_fd_sc_hd__and3_4
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11864__A _16113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19744_ _19744_/A _19744_/B _19793_/B _19743_/X VGND VGND VPWR VPWR _19765_/B sky130_fd_sc_hd__and4_4
XANTENNA__15336__A _12567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12079_ _11998_/A _12077_/X _12079_/C VGND VGND VPWR VPWR _12080_/C sky130_fd_sc_hd__and3_4
X_16956_ _16956_/A VGND VGND VPWR VPWR _16972_/A sky130_fd_sc_hd__inv_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14240__A _14252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22195__B2 _22190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15907_ _11657_/X _15907_/B _15907_/C VGND VGND VPWR VPWR _15907_/X sky130_fd_sc_hd__and3_4
X_19675_ HRDATA[24] VGND VGND VPWR VPWR _20800_/A sky130_fd_sc_hd__buf_2
XFILLER_38_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16887_ _16887_/A _16887_/B _16887_/C _16886_/X VGND VGND VPWR VPWR _16887_/X sky130_fd_sc_hd__and4_4
XANTENNA__20896__B _20342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18626_ _17639_/A _18606_/X _16927_/A _18625_/X VGND VGND VPWR VPWR _18626_/X sky130_fd_sc_hd__o22a_4
X_15838_ _12915_/A _15838_/B VGND VGND VPWR VPWR _15838_/X sky130_fd_sc_hd__or2_4
XFILLER_64_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22169__A _22169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18557_ _18557_/A _18556_/X VGND VGND VPWR VPWR _18557_/X sky130_fd_sc_hd__or2_4
X_15769_ _15750_/A _15769_/B VGND VGND VPWR VPWR _15771_/B sky130_fd_sc_hd__or2_4
XFILLER_55_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12695__A _12695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22498__A2 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17508_ _13278_/X _17510_/B VGND VGND VPWR VPWR _17508_/X sky130_fd_sc_hd__or2_4
XFILLER_94_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18488_ _17621_/D _17621_/C _17599_/Y VGND VGND VPWR VPWR _18488_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21170__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _12924_/X VGND VGND VPWR VPWR _17439_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19478__A _19598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20450_ _24406_/Q _20405_/X _24438_/Q _20449_/X VGND VGND VPWR VPWR _20450_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19109_ _24288_/Q _19108_/X VGND VGND VPWR VPWR _19110_/B sky130_fd_sc_hd__and2_4
XFILLER_118_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20381_ _20407_/A _20378_/Y _20380_/X _18961_/Y _20253_/X VGND VGND VPWR VPWR _20381_/X
+ sky130_fd_sc_hd__a32o_4
X_22120_ _22108_/A VGND VGND VPWR VPWR _22120_/X sky130_fd_sc_hd__buf_2
XFILLER_115_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22051_ _21838_/X _22045_/X _23466_/Q _22049_/X VGND VGND VPWR VPWR _22051_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21002_ _21293_/A VGND VGND VPWR VPWR _21002_/X sky130_fd_sc_hd__buf_2
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15246__A _14367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22953_ _22924_/X _18459_/A _22937_/X _22952_/X VGND VGND VPWR VPWR _22954_/A sky130_fd_sc_hd__a211o_4
XFILLER_60_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21933__B2 _21928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21904_ _21845_/X _21901_/X _23559_/Q _21898_/X VGND VGND VPWR VPWR _23559_/D sky130_fd_sc_hd__o22a_4
XFILLER_99_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17461__A _17156_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22884_ _22719_/X _22924_/A _22932_/A _19888_/X VGND VGND VPWR VPWR _22885_/A sky130_fd_sc_hd__or4_4
XANTENNA__22079__A _20338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21835_ _21265_/A VGND VGND VPWR VPWR _21835_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22489__A2 _22486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16077__A _16077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21697__B1 _16256_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21766_ _21752_/A VGND VGND VPWR VPWR _21766_/X sky130_fd_sc_hd__buf_2
XFILLER_52_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20717_ _20717_/A VGND VGND VPWR VPWR _20717_/Y sky130_fd_sc_hd__inv_2
X_23505_ _24082_/CLK _21991_/X VGND VGND VPWR VPWR _13138_/B sky130_fd_sc_hd__dfxtp_4
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21697_ _21517_/X _21691_/X _16256_/B _21695_/X VGND VGND VPWR VPWR _23673_/D sky130_fd_sc_hd__o22a_4
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16805__A _16747_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23436_ _23698_/CLK _22118_/X VGND VGND VPWR VPWR _15474_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20648_ _20644_/X VGND VGND VPWR VPWR _20754_/B sky130_fd_sc_hd__buf_2
XANTENNA__17117__A1 _13048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17117__B2 _17032_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20327__A _20497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23367_ _23591_/CLK _22239_/X VGND VGND VPWR VPWR _23367_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17668__A2 _17442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20579_ _24400_/Q _20405_/X _24432_/Q _20449_/X VGND VGND VPWR VPWR _20579_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14325__A _15571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22661__A2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13120_ _13080_/A _13120_/B VGND VGND VPWR VPWR _13121_/C sky130_fd_sc_hd__or2_4
X_22318_ _23308_/Q VGND VGND VPWR VPWR _22318_/X sky130_fd_sc_hd__buf_2
XANTENNA__20672__A1 _20613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20672__B2 _20592_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23298_ _23812_/CLK _22328_/X VGND VGND VPWR VPWR _15269_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13051_ _12465_/A _13051_/B _13051_/C VGND VGND VPWR VPWR _13051_/X sky130_fd_sc_hd__and3_4
X_22249_ _22147_/X _22222_/A _15097_/B _22212_/A VGND VGND VPWR VPWR _22249_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12002_ _11998_/A _12000_/X _12002_/C VGND VGND VPWR VPWR _12006_/B sky130_fd_sc_hd__and3_4
XFILLER_87_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16810_ _16597_/X _16802_/X _16810_/C VGND VGND VPWR VPWR _16811_/C sky130_fd_sc_hd__and3_4
XANTENNA__15156__A _11954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11684__A _16198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17790_ _17790_/A VGND VGND VPWR VPWR _17790_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22177__B2 _22176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16741_ _16741_/A _16741_/B VGND VGND VPWR VPWR _16741_/X sky130_fd_sc_hd__and2_4
X_13953_ _13953_/A _14025_/B VGND VGND VPWR VPWR _13955_/B sky130_fd_sc_hd__or2_4
XFILLER_78_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18467__A _18421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12904_ _12904_/A _23379_/Q VGND VGND VPWR VPWR _12904_/X sky130_fd_sc_hd__or2_4
X_19460_ _19433_/A VGND VGND VPWR VPWR _19460_/X sky130_fd_sc_hd__buf_2
XANTENNA__17371__A _15782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16672_ _16630_/X _16672_/B VGND VGND VPWR VPWR _16672_/X sky130_fd_sc_hd__or2_4
XFILLER_62_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23532__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13884_ _13884_/A _13884_/B _13884_/C VGND VGND VPWR VPWR _13885_/C sky130_fd_sc_hd__or3_4
XFILLER_61_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18411_ _18340_/X _18408_/X _18377_/X _18410_/X VGND VGND VPWR VPWR _18411_/X sky130_fd_sc_hd__o22a_4
X_15623_ _15623_/A _15621_/X _15623_/C VGND VGND VPWR VPWR _15623_/X sky130_fd_sc_hd__and3_4
X_12835_ _12827_/A _23220_/Q VGND VGND VPWR VPWR _12837_/B sky130_fd_sc_hd__or2_4
X_19391_ _19389_/X _18356_/X _19389_/X _24207_/Q VGND VGND VPWR VPWR _24207_/D sky130_fd_sc_hd__a2bb2o_4
X_18342_ _18342_/A _18341_/Y VGND VGND VPWR VPWR _18354_/A sky130_fd_sc_hd__or2_4
X_15554_ _12307_/A _15554_/B _15553_/X VGND VGND VPWR VPWR _15554_/X sky130_fd_sc_hd__and3_4
XFILLER_76_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12766_ _12765_/X VGND VGND VPWR VPWR _12769_/A sky130_fd_sc_hd__buf_2
XFILLER_72_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21152__A2 _21147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14500_/X _14505_/B VGND VGND VPWR VPWR _14505_/X sky130_fd_sc_hd__or2_4
X_11717_ _16072_/A VGND VGND VPWR VPWR _11717_/X sky130_fd_sc_hd__buf_2
X_18273_ _17961_/X _18269_/Y _18076_/X _18272_/Y VGND VGND VPWR VPWR _18273_/X sky130_fd_sc_hd__a211o_4
XANTENNA__19298__A _22924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12198_/X VGND VGND VPWR VPWR _15664_/A sky130_fd_sc_hd__buf_2
X_15485_ _11664_/A _15469_/X _15484_/X VGND VGND VPWR VPWR _15485_/X sky130_fd_sc_hd__or3_4
XFILLER_15_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17224_ _17224_/A _17222_/X VGND VGND VPWR VPWR _17224_/X sky130_fd_sc_hd__or2_4
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _12578_/A VGND VGND VPWR VPWR _11648_/X sky130_fd_sc_hd__buf_2
X_14436_ _14463_/A _14502_/B VGND VGND VPWR VPWR _14436_/X sky130_fd_sc_hd__or2_4
XFILLER_54_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17155_ _17173_/A VGND VGND VPWR VPWR _17155_/X sky130_fd_sc_hd__buf_2
X_11579_ _17052_/A _16909_/B VGND VGND VPWR VPWR _11579_/X sky130_fd_sc_hd__or2_4
X_14367_ _14367_/A VGND VGND VPWR VPWR _15604_/A sky130_fd_sc_hd__buf_2
XANTENNA__22652__A2 _22650_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14235__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16106_ _16091_/A VGND VGND VPWR VPWR _16107_/A sky130_fd_sc_hd__buf_2
X_13318_ _13286_/X _13318_/B VGND VGND VPWR VPWR _13318_/X sky130_fd_sc_hd__or2_4
XANTENNA__21860__B1 _23585_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14298_ _12459_/A _14298_/B _14298_/C VGND VGND VPWR VPWR _14298_/X sky130_fd_sc_hd__or3_4
X_17086_ _18048_/A VGND VGND VPWR VPWR _18240_/A sky130_fd_sc_hd__inv_2
XANTENNA__19745__B _19873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22452__A _22384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16037_ _16037_/A _23672_/Q VGND VGND VPWR VPWR _16039_/B sky130_fd_sc_hd__or2_4
X_13249_ _13242_/A _13249_/B VGND VGND VPWR VPWR _13250_/C sky130_fd_sc_hd__or2_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14889__B _14889_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21068__A _21075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11594__A _11594_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19761__A HRDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17988_ _18189_/A VGND VGND VPWR VPWR _18216_/A sky130_fd_sc_hd__buf_2
XANTENNA__24464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19727_ _19719_/A VGND VGND VPWR VPWR _19730_/A sky130_fd_sc_hd__buf_2
XFILLER_111_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16939_ _16939_/A VGND VGND VPWR VPWR _16989_/A sky130_fd_sc_hd__inv_2
XANTENNA__20700__A _20342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18377__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19658_ _19483_/X VGND VGND VPWR VPWR _19661_/A sky130_fd_sc_hd__inv_2
XFILLER_80_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21391__A2 _21390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18609_ _18556_/X VGND VGND VPWR VPWR _18609_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19589_ _20358_/B _19551_/X _19588_/X _19554_/X VGND VGND VPWR VPWR _19589_/X sky130_fd_sc_hd__a211o_4
XFILLER_53_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21620_ _21555_/X _21619_/X _23721_/Q _21616_/X VGND VGND VPWR VPWR _23721_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13314__A _13317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17347__A1 _17339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18544__B1 _18500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17347__B2 _17346_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21143__A2 _21140_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21551_ _21527_/A VGND VGND VPWR VPWR _21551_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20502_ _20502_/A _20502_/B VGND VGND VPWR VPWR _20502_/Y sky130_fd_sc_hd__nor2_4
X_24270_ _24092_/CLK _24270_/D HRESETn VGND VGND VPWR VPWR _19219_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_53_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24330__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21482_ _21265_/X _21477_/X _23787_/Q _21481_/X VGND VGND VPWR VPWR _21482_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23221_ _23983_/CLK _23221_/D VGND VGND VPWR VPWR _12667_/B sky130_fd_sc_hd__dfxtp_4
X_20433_ _20292_/X _20432_/X _19132_/A _20305_/X VGND VGND VPWR VPWR _20433_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11769__A _13102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18847__A1 _15646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14145__A _14145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23152_ _23473_/CLK _23152_/D VGND VGND VPWR VPWR _13311_/B sky130_fd_sc_hd__dfxtp_4
X_20364_ _20322_/X _20363_/X _24346_/Q _20247_/X VGND VGND VPWR VPWR _20364_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23405__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22103_ _20552_/A VGND VGND VPWR VPWR _22103_/X sky130_fd_sc_hd__buf_2
XANTENNA__16998__C _16997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23083_ _24044_/CLK _23083_/D VGND VGND VPWR VPWR _15573_/B sky130_fd_sc_hd__dfxtp_4
X_20295_ _20556_/A VGND VGND VPWR VPWR _20519_/B sky130_fd_sc_hd__buf_2
XANTENNA__16360__A _11715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22034_ _21809_/X _22031_/X _12312_/B _22028_/X VGND VGND VPWR VPWR _22034_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21603__B1 _12586_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19671__A _19722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22159__B2 _22155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23985_ _24082_/CLK _21136_/X VGND VGND VPWR VPWR _23985_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20610__A _20610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21906__B2 _21905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17191__A _15517_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19575__A2 _19706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15704__A _12743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22936_ _22936_/A VGND VGND VPWR VPWR HADDR[9] sky130_fd_sc_hd__inv_2
XFILLER_112_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21382__A2 _21376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22867_ _22854_/X _22807_/X _14074_/A _22855_/X VGND VGND VPWR VPWR _22867_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13224__A _13260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12620_ _12660_/A _12620_/B VGND VGND VPWR VPWR _12620_/X sky130_fd_sc_hd__or2_4
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21818_ _21816_/X _21817_/X _23603_/Q _21812_/X VGND VGND VPWR VPWR _21818_/X sky130_fd_sc_hd__o22a_4
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22798_ _22807_/A _15051_/X VGND VGND VPWR VPWR _22798_/X sky130_fd_sc_hd__or2_4
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17338__A1 _14425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21134__A2 _21133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ _13032_/A _12658_/B VGND VGND VPWR VPWR _12552_/C sky130_fd_sc_hd__or2_4
X_21749_ _21519_/X _21748_/X _23640_/Q _21745_/X VGND VGND VPWR VPWR _21749_/X sky130_fd_sc_hd__o22a_4
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11502_ _24384_/Q VGND VGND VPWR VPWR _20965_/A sky130_fd_sc_hd__inv_2
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _11610_/A VGND VGND VPWR VPWR _13953_/A sky130_fd_sc_hd__buf_2
X_15270_ _14161_/A _15343_/B VGND VGND VPWR VPWR _15271_/C sky130_fd_sc_hd__or2_4
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24174__D _19783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24468_ _23522_/CLK _18229_/X HRESETn VGND VGND VPWR VPWR _24468_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ _13686_/A _14221_/B _14220_/X VGND VGND VPWR VPWR _14221_/X sky130_fd_sc_hd__or3_4
XANTENNA__11679__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23419_ _23293_/CLK _23419_/D VGND VGND VPWR VPWR _16792_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18838__A1 _13274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19846__A _19872_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24399_ _24334_/CLK _24399_/D HRESETn VGND VGND VPWR VPWR _20595_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14055__A _14055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22634__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14152_ _14152_/A _24073_/Q VGND VGND VPWR VPWR _14153_/C sky130_fd_sc_hd__or2_4
XANTENNA__23085__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22272__A _22272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13103_ _12957_/A _13103_/B _13103_/C VGND VGND VPWR VPWR _13135_/B sky130_fd_sc_hd__or3_4
X_14083_ _14083_/A _23337_/Q VGND VGND VPWR VPWR _14083_/X sky130_fd_sc_hd__or2_4
X_18960_ _18958_/Y _18959_/Y _11530_/X VGND VGND VPWR VPWR _18960_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16270__A _11980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13034_ _12891_/A _13030_/X _13034_/C VGND VGND VPWR VPWR _13034_/X sky130_fd_sc_hd__or3_4
X_17911_ _17911_/A VGND VGND VPWR VPWR _17911_/X sky130_fd_sc_hd__buf_2
X_18891_ _18891_/A VGND VGND VPWR VPWR _18891_/X sky130_fd_sc_hd__buf_2
X_17842_ _17814_/X _17213_/X _17815_/X _17209_/X VGND VGND VPWR VPWR _17842_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21070__B2 _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12303__A _12459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21616__A _21602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17773_ _11629_/X _17772_/X _24477_/Q _11629_/X VGND VGND VPWR VPWR _24477_/D sky130_fd_sc_hd__a2bb2o_4
X_14985_ _11798_/A _14985_/B _14985_/C VGND VGND VPWR VPWR _14986_/C sky130_fd_sc_hd__or3_4
X_19512_ _19754_/A VGND VGND VPWR VPWR _19523_/B sky130_fd_sc_hd__inv_2
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16724_ _12091_/A _16792_/B VGND VGND VPWR VPWR _16725_/C sky130_fd_sc_hd__or2_4
X_13936_ _15037_/A _23754_/Q VGND VGND VPWR VPWR _13937_/C sky130_fd_sc_hd__or2_4
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12957__B _12957_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19443_ _19450_/A VGND VGND VPWR VPWR _19839_/A sky130_fd_sc_hd__inv_2
XANTENNA__22570__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16655_ _16610_/A _23836_/Q VGND VGND VPWR VPWR _16656_/C sky130_fd_sc_hd__or2_4
XANTENNA__15333__B _15274_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13867_ _13878_/A _23911_/Q VGND VGND VPWR VPWR _13869_/B sky130_fd_sc_hd__or2_4
XFILLER_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15606_ _15618_/A _23979_/Q VGND VGND VPWR VPWR _15607_/C sky130_fd_sc_hd__or2_4
XFILLER_50_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13134__A _12672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12818_ _12802_/A _23380_/Q VGND VGND VPWR VPWR _12818_/X sky130_fd_sc_hd__or2_4
X_19374_ _19370_/A VGND VGND VPWR VPWR _19374_/X sky130_fd_sc_hd__buf_2
X_16586_ _16586_/A _23100_/Q VGND VGND VPWR VPWR _16586_/X sky130_fd_sc_hd__or2_4
X_13798_ _15413_/A _23911_/Q VGND VGND VPWR VPWR _13798_/X sky130_fd_sc_hd__or2_4
XANTENNA__18526__B1 _18063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22447__A _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18325_ _18324_/X VGND VGND VPWR VPWR _18425_/B sky130_fd_sc_hd__inv_2
XANTENNA__21351__A _21373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15537_ _15556_/A _23979_/Q VGND VGND VPWR VPWR _15537_/X sky130_fd_sc_hd__or2_4
X_12749_ _11850_/A _12748_/X VGND VGND VPWR VPWR _12749_/X sky130_fd_sc_hd__and2_4
XANTENNA__16445__A _11702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18256_ _18239_/X _18245_/Y _18252_/X _18254_/X _18255_/Y VGND VGND VPWR VPWR _18256_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20884__B2 _20686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15468_ _13731_/A _15464_/X _15468_/C VGND VGND VPWR VPWR _15469_/C sky130_fd_sc_hd__or3_4
XFILLER_50_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23428__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16164__B _16092_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17207_ _17152_/X _17205_/X _17154_/X _17206_/X VGND VGND VPWR VPWR _17207_/X sky130_fd_sc_hd__o22a_4
X_14419_ _13896_/A _14417_/X _14419_/C VGND VGND VPWR VPWR _14420_/C sky130_fd_sc_hd__and3_4
XANTENNA__18829__A1 _16374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18187_ _17259_/A _18186_/Y VGND VGND VPWR VPWR _18187_/X sky130_fd_sc_hd__and2_4
XANTENNA__22625__A2 _22622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15399_ _15399_/A _15462_/B VGND VGND VPWR VPWR _15401_/B sky130_fd_sc_hd__or2_4
X_17138_ _17157_/A VGND VGND VPWR VPWR _17138_/X sky130_fd_sc_hd__buf_2
XFILLER_102_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17069_ _17069_/A _17068_/A _11591_/D _18866_/B VGND VGND VPWR VPWR _17069_/X sky130_fd_sc_hd__or4_4
XANTENNA__23578__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16180__A _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22389__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20080_ _20176_/A _20078_/X _20079_/Y _19936_/X VGND VGND VPWR VPWR _20080_/X sky130_fd_sc_hd__o22a_4
XFILLER_48_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13309__A _15667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12213__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15524__A _12320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23770_ _23770_/CLK _23770_/D VGND VGND VPWR VPWR _16388_/B sky130_fd_sc_hd__dfxtp_4
X_20982_ _21291_/A VGND VGND VPWR VPWR _20982_/X sky130_fd_sc_hd__buf_2
XFILLER_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21364__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22561__B2 _22518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22721_ _22714_/X VGND VGND VPWR VPWR _22721_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18835__A _18835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13044__A _13017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22652_ _22442_/X _22650_/X _13660_/B _22647_/X VGND VGND VPWR VPWR _22652_/X sky130_fd_sc_hd__o22a_4
XFILLER_13_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24203__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21603_ _21526_/X _21598_/X _12586_/B _21602_/X VGND VGND VPWR VPWR _21603_/X sky130_fd_sc_hd__o22a_4
XFILLER_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13979__A _12302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22583_ _22583_/A VGND VGND VPWR VPWR _22583_/X sky130_fd_sc_hd__buf_2
XANTENNA__12883__A _12883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21534_ _21249_/A VGND VGND VPWR VPWR _21534_/X sky130_fd_sc_hd__buf_2
X_24322_ _24321_/CLK _19096_/X HRESETn VGND VGND VPWR VPWR _19092_/A sky130_fd_sc_hd__dfstp_4
XFILLER_90_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24253_ _24250_/CLK _24253_/D HRESETn VGND VGND VPWR VPWR _24253_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21465_ _21237_/X _21463_/X _16217_/B _21460_/X VGND VGND VPWR VPWR _23799_/D sky130_fd_sc_hd__o22a_4
X_23204_ _23812_/CLK _23204_/D VGND VGND VPWR VPWR _14627_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22804__B _17115_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20627__A1 _20622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20416_ _20588_/A _20415_/X VGND VGND VPWR VPWR _20416_/Y sky130_fd_sc_hd__nand2_4
XFILLER_88_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20627__B2 _20497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24184_ _24162_/CLK _19636_/X HRESETn VGND VGND VPWR VPWR _17543_/A sky130_fd_sc_hd__dfrtp_4
X_21396_ _21293_/X _21369_/A _23839_/Q _21359_/A VGND VGND VPWR VPWR _21396_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12107__B _23805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23135_ _23889_/CLK _23135_/D VGND VGND VPWR VPWR _23135_/Q sky130_fd_sc_hd__dfxtp_4
X_20347_ _20322_/X _20346_/X _11532_/A _20247_/X VGND VGND VPWR VPWR _20347_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24386__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23066_ VGND VGND VPWR VPWR _24108_/D _23066_/LO sky130_fd_sc_hd__conb_1
X_20278_ _20188_/Y _20203_/X _20203_/X _20277_/X VGND VGND VPWR VPWR _24094_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22017_ _22017_/A _22017_/B _20199_/A _21212_/B VGND VGND VPWR VPWR _22017_/X sky130_fd_sc_hd__or4_4
XFILLER_88_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13219__A _11671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21052__B2 _21048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18599__A3 _18594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_56_0_HCLK clkbuf_6_28_0_HCLK/X VGND VGND VPWR VPWR _23692_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__11962__A _16139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15434__A _15411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14770_ _13799_/A _14770_/B VGND VGND VPWR VPWR _14771_/C sky130_fd_sc_hd__or2_4
XFILLER_99_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24169__D _24169_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11982_ _11982_/A VGND VGND VPWR VPWR _11982_/X sky130_fd_sc_hd__buf_2
X_23968_ _24032_/CLK _21159_/X VGND VGND VPWR VPWR _14873_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_112_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22552__B2 _22547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13721_ _13747_/A _13714_/X _13721_/C VGND VGND VPWR VPWR _13721_/X sky130_fd_sc_hd__or3_4
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22919_ _22919_/A VGND VGND VPWR VPWR HADDR[6] sky130_fd_sc_hd__inv_2
X_23899_ _23515_/CLK _23899_/D VGND VGND VPWR VPWR _23899_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16440_ _11861_/X _16436_/X _16440_/C VGND VGND VPWR VPWR _16440_/X sky130_fd_sc_hd__or3_4
X_13652_ _12475_/A _13652_/B VGND VGND VPWR VPWR _13652_/X sky130_fd_sc_hd__or2_4
XANTENNA__21107__A2 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14992__B _15056_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12603_ _12650_/A VGND VGND VPWR VPWR _12604_/A sky130_fd_sc_hd__buf_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16371_ _11673_/X _16362_/X _16371_/C VGND VGND VPWR VPWR _16372_/C sky130_fd_sc_hd__and3_4
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13583_ _13582_/X VGND VGND VPWR VPWR _13583_/Y sky130_fd_sc_hd__inv_2
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12793__A _12802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16265__A _15937_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18110_ _17797_/X _18108_/X _17846_/X _18109_/X VGND VGND VPWR VPWR _18110_/X sky130_fd_sc_hd__o22a_4
X_15322_ _13871_/A _15259_/B VGND VGND VPWR VPWR _15324_/B sky130_fd_sc_hd__or2_4
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12534_ _13041_/A VGND VGND VPWR VPWR _12876_/A sky130_fd_sc_hd__buf_2
X_19090_ _18965_/A _19088_/Y _19089_/Y _19084_/X VGND VGND VPWR VPWR _19090_/X sky130_fd_sc_hd__o22a_4
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18041_ _17797_/X _17850_/X _17254_/X VGND VGND VPWR VPWR _18041_/X sky130_fd_sc_hd__o21a_4
X_15253_ _11954_/A _15253_/B VGND VGND VPWR VPWR _15254_/C sky130_fd_sc_hd__or2_4
XANTENNA__13401__B _13325_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12465_ _12465_/A VGND VGND VPWR VPWR _12917_/A sky130_fd_sc_hd__buf_2
XANTENNA__18480__A _18198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14204_ _14204_/A _23913_/Q VGND VGND VPWR VPWR _14206_/B sky130_fd_sc_hd__or2_4
XANTENNA__23720__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22714__B HREADY VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12396_ _12418_/A _12289_/B VGND VGND VPWR VPWR _12396_/X sky130_fd_sc_hd__or2_4
X_15184_ _12267_/X _15161_/X _15168_/X _15175_/X _15183_/X VGND VGND VPWR VPWR _15184_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_67_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14135_ _14108_/A _14135_/B _14134_/X VGND VGND VPWR VPWR _14136_/C sky130_fd_sc_hd__and3_4
XFILLER_4_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19992_ _19970_/X _16985_/A _19976_/X _19991_/X VGND VGND VPWR VPWR _19992_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14513__A _11740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14066_ _11647_/A _14066_/B VGND VGND VPWR VPWR _14069_/B sky130_fd_sc_hd__or2_4
X_18943_ _24348_/Q _11532_/X _18926_/C _18942_/Y VGND VGND VPWR VPWR _18943_/X sky130_fd_sc_hd__o22a_4
XFILLER_45_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13017_ _13017_/A _13017_/B _13017_/C VGND VGND VPWR VPWR _13018_/C sky130_fd_sc_hd__and3_4
XANTENNA__13129__A _13129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21043__B2 _21041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18874_ _18898_/A VGND VGND VPWR VPWR _18891_/A sky130_fd_sc_hd__buf_2
XFILLER_80_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12033__A _18728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17825_ _17825_/A VGND VGND VPWR VPWR _17825_/X sky130_fd_sc_hd__buf_2
XANTENNA__12968__A _12980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11872__A _12493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15344__A _14009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17756_ _17662_/X _17690_/A VGND VGND VPWR VPWR _17756_/Y sky130_fd_sc_hd__nand2_4
X_14968_ _14642_/A _14968_/B _14967_/X VGND VGND VPWR VPWR _14968_/X sky130_fd_sc_hd__or3_4
XFILLER_78_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21346__A2 _21319_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12687__B _12768_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16707_ _11888_/A _16767_/B VGND VGND VPWR VPWR _16709_/B sky130_fd_sc_hd__or2_4
XFILLER_75_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13919_ _13918_/X VGND VGND VPWR VPWR _13921_/B sky130_fd_sc_hd__inv_2
XFILLER_63_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17687_ _17669_/X _17684_/X _17686_/X VGND VGND VPWR VPWR _17687_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20554__B1 _24082_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14899_ _14867_/X _14899_/B VGND VGND VPWR VPWR _14899_/X sky130_fd_sc_hd__or2_4
XFILLER_78_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18655__A _18498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19426_ HRDATA[16] _16996_/A _19425_/Y _24142_/Q _19416_/B VGND VGND VPWR VPWR _19426_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_62_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16638_ _16651_/A _23996_/Q VGND VGND VPWR VPWR _16639_/C sky130_fd_sc_hd__or2_4
XFILLER_91_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23250__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17970__B2 _17816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19357_ _19355_/X _19356_/Y _19355_/X _24225_/Q VGND VGND VPWR VPWR _19357_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13799__A _13799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14784__A1 _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16569_ _16569_/A _16569_/B _16569_/C VGND VGND VPWR VPWR _16570_/C sky130_fd_sc_hd__and3_4
XFILLER_17_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18308_ _18307_/A _18307_/B _18048_/X VGND VGND VPWR VPWR _18308_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_91_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19288_ _19209_/A _19209_/B _19287_/Y VGND VGND VPWR VPWR _24260_/D sky130_fd_sc_hd__o21a_4
XFILLER_108_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18239_ _18239_/A _17447_/X VGND VGND VPWR VPWR _18239_/X sky130_fd_sc_hd__or2_4
XANTENNA__18390__A _18390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20609__A1 _24207_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21250_ _21249_/X _21247_/X _23922_/Q _21242_/X VGND VGND VPWR VPWR _21250_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19475__A1 _24156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17718__B _17287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20201_ _20279_/A VGND VGND VPWR VPWR _20488_/A sky130_fd_sc_hd__inv_2
X_21181_ _20487_/X _21176_/X _12640_/B _21180_/X VGND VGND VPWR VPWR _21181_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15519__A _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14423__A _13918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20132_ _24449_/Q VGND VGND VPWR VPWR _20132_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22640__A _22633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13039__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20063_ _18552_/X _20057_/X _20062_/Y _20044_/X VGND VGND VPWR VPWR _20063_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15254__A _14098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11782__A _11782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23822_ _23922_/CLK _21427_/X VGND VGND VPWR VPWR _15690_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22534__A1 _22410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22534__B2 _22533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20965_ _20965_/A _18813_/X VGND VGND VPWR VPWR _20965_/X sky130_fd_sc_hd__or2_4
X_23753_ _24011_/CLK _21557_/X VGND VGND VPWR VPWR _23753_/Q sky130_fd_sc_hd__dfxtp_4
X_22704_ _22683_/A VGND VGND VPWR VPWR _22704_/X sky130_fd_sc_hd__buf_2
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13027__A1 _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20896_ _20849_/B _20342_/B VGND VGND VPWR VPWR _20896_/X sky130_fd_sc_hd__or2_4
X_23684_ _23363_/CLK _21677_/X VGND VGND VPWR VPWR _14706_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22635_ _22413_/X _22629_/X _23124_/Q _22633_/X VGND VGND VPWR VPWR _22635_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22566_ _22566_/A VGND VGND VPWR VPWR _22600_/A sky130_fd_sc_hd__buf_2
XFILLER_22_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21517_ _21802_/A VGND VGND VPWR VPWR _21517_/X sky130_fd_sc_hd__buf_2
X_24305_ _24305_/CLK _24305_/D HRESETn VGND VGND VPWR VPWR _24305_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13221__B _23569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22497_ _22483_/A VGND VGND VPWR VPWR _22497_/X sky130_fd_sc_hd__buf_2
XFILLER_6_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12250_ _12250_/A VGND VGND VPWR VPWR _13985_/A sky130_fd_sc_hd__buf_2
X_21448_ _21005_/A VGND VGND VPWR VPWR _21784_/A sky130_fd_sc_hd__buf_2
X_24236_ _24239_/CLK _19339_/X HRESETn VGND VGND VPWR VPWR _24236_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11957__A _15707_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12181_ _11675_/X _12181_/B _12180_/X VGND VGND VPWR VPWR _12182_/C sky130_fd_sc_hd__and3_4
X_24167_ _23584_/CLK _19844_/Y HRESETn VGND VGND VPWR VPWR _21583_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15429__A _15429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21379_ _21263_/X _21376_/X _23852_/Q _21373_/X VGND VGND VPWR VPWR _21379_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14333__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17554__A1_N _16008_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23118_ _23564_/CLK _22644_/X VGND VGND VPWR VPWR _15689_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_1_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24098_ _24290_/CLK _24098_/D HRESETn VGND VGND VPWR VPWR _22731_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22550__A _22521_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17229__B1 _15381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15940_ _15952_/A _23736_/Q VGND VGND VPWR VPWR _15941_/C sky130_fd_sc_hd__or2_4
X_23049_ _19925_/X _17769_/A _23026_/X _23048_/X VGND VGND VPWR VPWR _23050_/A sky130_fd_sc_hd__a211o_4
XANTENNA__23123__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21025__B2 _21020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21166__A _21165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15871_ _13554_/A _15802_/B VGND VGND VPWR VPWR _15871_/X sky130_fd_sc_hd__or2_4
XFILLER_95_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17610_ _17325_/X VGND VGND VPWR VPWR _17610_/Y sky130_fd_sc_hd__inv_2
X_14822_ _14841_/A _14758_/B VGND VGND VPWR VPWR _14822_/X sky130_fd_sc_hd__or2_4
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15164__A _14098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18590_ _17858_/X _18115_/Y _17854_/X _18589_/Y VGND VGND VPWR VPWR _18591_/A sky130_fd_sc_hd__a211o_4
XFILLER_40_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21328__A2 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22525__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17541_ _17627_/A VGND VGND VPWR VPWR _17569_/A sky130_fd_sc_hd__inv_2
X_14753_ _11976_/A _14752_/X VGND VGND VPWR VPWR _14753_/X sky130_fd_sc_hd__and2_4
X_11965_ _11998_/A _11965_/B _11965_/C VGND VGND VPWR VPWR _11973_/B sky130_fd_sc_hd__and3_4
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13704_ _13765_/A _13702_/X _13704_/C VGND VGND VPWR VPWR _13705_/C sky130_fd_sc_hd__and3_4
X_17472_ _17471_/X VGND VGND VPWR VPWR _17472_/Y sky130_fd_sc_hd__inv_2
X_14684_ _15592_/A _14682_/X _14683_/X VGND VGND VPWR VPWR _14684_/X sky130_fd_sc_hd__and3_4
XFILLER_60_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11896_ _14463_/A VGND VGND VPWR VPWR _12852_/A sky130_fd_sc_hd__buf_2
XFILLER_71_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19211_ _19211_/A _19211_/B VGND VGND VPWR VPWR _19212_/B sky130_fd_sc_hd__and2_4
X_16423_ _16400_/A _16423_/B VGND VGND VPWR VPWR _16423_/X sky130_fd_sc_hd__or2_4
X_13635_ _13635_/A VGND VGND VPWR VPWR _13636_/A sky130_fd_sc_hd__buf_2
XANTENNA__14508__A _13890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19142_ _19138_/A _19137_/X _19140_/Y VGND VGND VPWR VPWR _24317_/D sky130_fd_sc_hd__o21a_4
X_16354_ _11770_/X _16354_/B _16353_/X VGND VGND VPWR VPWR _16372_/B sky130_fd_sc_hd__and3_4
X_13566_ _13554_/A _13566_/B VGND VGND VPWR VPWR _13567_/C sky130_fd_sc_hd__or2_4
XFILLER_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15305_ _14603_/A _15303_/X _15305_/C VGND VGND VPWR VPWR _15305_/X sky130_fd_sc_hd__and3_4
XFILLER_34_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12517_ _13491_/A _12458_/X _12480_/X _12503_/X _12516_/X VGND VGND VPWR VPWR _12517_/X
+ sky130_fd_sc_hd__a32o_4
X_19073_ _19052_/X _19071_/Y _19072_/Y _19057_/X VGND VGND VPWR VPWR _19073_/X sky130_fd_sc_hd__o22a_4
XFILLER_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16285_ _16152_/A _16281_/X _16285_/C VGND VGND VPWR VPWR _16285_/X sky130_fd_sc_hd__or3_4
X_13497_ _12926_/A VGND VGND VPWR VPWR _15884_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18024_ _18239_/A _18024_/B VGND VGND VPWR VPWR _18024_/X sky130_fd_sc_hd__or2_4
X_15236_ _14251_/A _23681_/Q VGND VGND VPWR VPWR _15238_/B sky130_fd_sc_hd__or2_4
X_12448_ _14748_/A VGND VGND VPWR VPWR _12449_/A sky130_fd_sc_hd__buf_2
XFILLER_8_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20245__A _20248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_11_0_HCLK_A clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15167_ _15144_/A _15165_/X _15166_/X VGND VGND VPWR VPWR _15167_/X sky130_fd_sc_hd__and3_4
XANTENNA__21264__B2 _21254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12379_ _13211_/A VGND VGND VPWR VPWR _15889_/A sky130_fd_sc_hd__buf_2
XANTENNA__14243__A _14243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14118_ _12531_/A _14118_/B _14117_/X VGND VGND VPWR VPWR _14118_/X sky130_fd_sc_hd__or3_4
XFILLER_4_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15098_ _15110_/A _23391_/Q VGND VGND VPWR VPWR _15099_/C sky130_fd_sc_hd__or2_4
X_19975_ _19974_/X VGND VGND VPWR VPWR _24137_/D sky130_fd_sc_hd__inv_2
XANTENNA__22460__A _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22213__B1 _16423_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14049_ _12568_/A _23818_/Q VGND VGND VPWR VPWR _14050_/C sky130_fd_sc_hd__or2_4
X_18926_ _18923_/Y _18924_/Y _18926_/C _18934_/A VGND VGND VPWR VPWR _18926_/X sky130_fd_sc_hd__and4_4
XFILLER_45_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18857_ _14564_/X _18855_/X _20854_/A _18856_/X VGND VGND VPWR VPWR _24389_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20775__B1 _20774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12698__A _12710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15074__A _15074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17808_ _17804_/A VGND VGND VPWR VPWR _17808_/X sky130_fd_sc_hd__buf_2
X_18788_ _18788_/A VGND VGND VPWR VPWR _18788_/X sky130_fd_sc_hd__buf_2
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17739_ _16997_/A _17122_/X _16997_/A _17122_/X VGND VGND VPWR VPWR _17739_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20750_ _20279_/A VGND VGND VPWR VPWR _20750_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15802__A _12477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19409_ _19377_/X _18682_/X _19380_/X _24194_/Q VGND VGND VPWR VPWR _19409_/X sky130_fd_sc_hd__o22a_4
X_20681_ _20253_/X VGND VGND VPWR VPWR _20681_/X sky130_fd_sc_hd__buf_2
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22420_ _20573_/A VGND VGND VPWR VPWR _22420_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22351_ _22351_/A VGND VGND VPWR VPWR _22351_/X sky130_fd_sc_hd__buf_2
X_21302_ _21301_/X VGND VGND VPWR VPWR _21302_/X sky130_fd_sc_hd__buf_2
XFILLER_40_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11991__A1 _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22282_ _22117_/X _22279_/X _15458_/B _22276_/X VGND VGND VPWR VPWR _22282_/X sky130_fd_sc_hd__o22a_4
X_24021_ _24021_/CLK _21080_/X VGND VGND VPWR VPWR _24021_/Q sky130_fd_sc_hd__dfxtp_4
X_21233_ _21232_/X _21223_/X _16263_/B _21230_/X VGND VGND VPWR VPWR _21233_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19944__A _17779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15249__A _11652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21255__B2 _21254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21164_ _21168_/A VGND VGND VPWR VPWR _21180_/A sky130_fd_sc_hd__inv_2
XFILLER_104_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20115_ _11552_/X VGND VGND VPWR VPWR _20115_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13992__A _13992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21095_ _20748_/X _21089_/X _24010_/Q _21093_/X VGND VGND VPWR VPWR _24010_/D sky130_fd_sc_hd__o22a_4
X_20046_ _20042_/X _18344_/X _20024_/X _20045_/X VGND VGND VPWR VPWR _20047_/A sky130_fd_sc_hd__o22a_4
XFILLER_115_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20230__A2 _20224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12401__A _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23805_ _23867_/CLK _21457_/X VGND VGND VPWR VPWR _23805_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12120__B _23517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21997_ _21831_/X _21995_/X _23501_/Q _21992_/X VGND VGND VPWR VPWR _21997_/X sky130_fd_sc_hd__o22a_4
XFILLER_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18295__A _18295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16808__A _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11717_/X _21498_/A VGND VGND VPWR VPWR _11750_/X sky130_fd_sc_hd__or2_4
X_23736_ _24084_/CLK _23736_/D VGND VGND VPWR VPWR _23736_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20403_/A _20947_/X _24257_/Q _20497_/A VGND VGND VPWR VPWR _20948_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21191__B1 _15748_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17934__B2 _17847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21730__A2 _21726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11680_/X VGND VGND VPWR VPWR _11681_/X sky130_fd_sc_hd__buf_2
X_23667_ _23987_/CLK _21706_/X VGND VGND VPWR VPWR _23667_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _20878_/Y _20851_/X _20490_/B _20675_/X VGND VGND VPWR VPWR _20879_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13378_/X _13337_/B VGND VGND VPWR VPWR _13421_/C sky130_fd_sc_hd__or2_4
XANTENNA__13232__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22618_ _22633_/A VGND VGND VPWR VPWR _22626_/A sky130_fd_sc_hd__buf_2
XFILLER_70_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23598_ _23692_/CLK _23598_/D VGND VGND VPWR VPWR _15685_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13351_ _12813_/A VGND VGND VPWR VPWR _13351_/X sky130_fd_sc_hd__buf_2
X_22549_ _22437_/X _22543_/X _14011_/B _22547_/X VGND VGND VPWR VPWR _23178_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21494__B2 _21488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16543__A _12020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12302_ _12302_/A VGND VGND VPWR VPWR _12459_/A sky130_fd_sc_hd__buf_2
X_16070_ _16058_/A _16070_/B _16070_/C VGND VGND VPWR VPWR _16070_/X sky130_fd_sc_hd__and3_4
XANTENNA__24182__D _19679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13282_ _12546_/A _13282_/B VGND VGND VPWR VPWR _13282_/X sky130_fd_sc_hd__or2_4
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15021_ _14994_/A _15021_/B _15021_/C VGND VGND VPWR VPWR _15021_/X sky130_fd_sc_hd__and3_4
X_12233_ _13678_/A VGND VGND VPWR VPWR _12233_/X sky130_fd_sc_hd__buf_2
X_24219_ _24216_/CLK _24219_/D HRESETn VGND VGND VPWR VPWR _24219_/Q sky130_fd_sc_hd__dfrtp_4
X_12164_ _11773_/X _12162_/X _12163_/X VGND VGND VPWR VPWR _12164_/X sky130_fd_sc_hd__and3_4
XFILLER_68_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14998__A _14998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12095_ _12068_/X _12095_/B _12095_/C VGND VGND VPWR VPWR _12096_/C sky130_fd_sc_hd__and3_4
X_16972_ _16972_/A _16972_/B VGND VGND VPWR VPWR _16973_/B sky130_fd_sc_hd__or2_4
X_19760_ _19710_/X _19753_/X _19759_/X _16597_/X _19697_/X VGND VGND VPWR VPWR _19760_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_46_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21549__A2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15923_ _15913_/B _15921_/Y _15783_/A _15922_/Y VGND VGND VPWR VPWR _15923_/X sky130_fd_sc_hd__a211o_4
X_18711_ _17330_/X _17331_/X _17330_/X _17331_/X VGND VGND VPWR VPWR _18711_/X sky130_fd_sc_hd__a2bb2o_4
X_19691_ _19691_/A VGND VGND VPWR VPWR _19877_/A sky130_fd_sc_hd__buf_2
XANTENNA__15606__B _23979_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18642_ _18642_/A VGND VGND VPWR VPWR _18644_/A sky130_fd_sc_hd__inv_2
X_15854_ _12413_/X _15852_/X _15853_/X VGND VGND VPWR VPWR _15854_/X sky130_fd_sc_hd__and3_4
XANTENNA__23789__CLK _23794_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12311__A _12745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_26_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_26_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14805_ _14813_/A _23139_/Q VGND VGND VPWR VPWR _14807_/B sky130_fd_sc_hd__or2_4
X_18573_ _18480_/X _18571_/X _18508_/X _18572_/X VGND VGND VPWR VPWR _18573_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13126__B _23474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15785_ _15785_/A _23501_/Q VGND VGND VPWR VPWR _15785_/X sky130_fd_sc_hd__or2_4
X_12997_ _13586_/A _12996_/X VGND VGND VPWR VPWR _16899_/A sky130_fd_sc_hd__or2_4
XANTENNA__19375__B1 _19374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17524_ _12990_/X _17524_/B VGND VGND VPWR VPWR _17524_/Y sky130_fd_sc_hd__nand2_4
XFILLER_73_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14736_ _14763_/A _14798_/B VGND VGND VPWR VPWR _14737_/C sky130_fd_sc_hd__or2_4
X_11948_ _16113_/A VGND VGND VPWR VPWR _12112_/A sky130_fd_sc_hd__buf_2
XANTENNA__21182__B1 _23956_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21721__A2 _21719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17455_ _17452_/X _17455_/B VGND VGND VPWR VPWR _17455_/X sky130_fd_sc_hd__or2_4
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14667_ _14666_/X _14667_/B VGND VGND VPWR VPWR _14667_/X sky130_fd_sc_hd__or2_4
XFILLER_92_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11879_ _11879_/A VGND VGND VPWR VPWR _15543_/A sky130_fd_sc_hd__buf_2
XANTENNA__14238__A _13839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16406_ _13447_/X _16404_/X _16406_/C VGND VGND VPWR VPWR _16406_/X sky130_fd_sc_hd__and3_4
XANTENNA__13142__A _12720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13618_ _13614_/A _13712_/B VGND VGND VPWR VPWR _13618_/X sky130_fd_sc_hd__or2_4
XFILLER_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17386_ _17383_/Y _17012_/A _17020_/A _17385_/X VGND VGND VPWR VPWR _17388_/A sky130_fd_sc_hd__o22a_4
X_14598_ _15026_/A _23908_/Q VGND VGND VPWR VPWR _14598_/X sky130_fd_sc_hd__or2_4
XFILLER_53_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19125_ _24304_/Q _19169_/A VGND VGND VPWR VPWR _19167_/A sky130_fd_sc_hd__and2_4
X_16337_ _13415_/A _16333_/X _16337_/C VGND VGND VPWR VPWR _16338_/C sky130_fd_sc_hd__or3_4
XFILLER_105_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13549_ _13548_/X _23823_/Q VGND VGND VPWR VPWR _13549_/X sky130_fd_sc_hd__or2_4
XANTENNA__17549__A _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21485__B2 _21481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12981__A _12981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19056_ _24361_/Q VGND VGND VPWR VPWR _19056_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16268_ _11872_/X _16266_/X _16267_/X VGND VGND VPWR VPWR _16268_/X sky130_fd_sc_hd__and3_4
X_18007_ _17888_/X _18006_/X _19977_/A _17888_/X VGND VGND VPWR VPWR _24474_/D sky130_fd_sc_hd__a2bb2o_4
X_15219_ _14182_/A _15156_/B VGND VGND VPWR VPWR _15219_/X sky130_fd_sc_hd__or2_4
XANTENNA__11597__A _11596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16199_ _16215_/A _16199_/B _16199_/C VGND VGND VPWR VPWR _16200_/C sky130_fd_sc_hd__and3_4
XANTENNA__22190__A _22169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20996__B1 _20640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19958_ _19985_/A _19955_/X _19956_/Y _19957_/X VGND VGND VPWR VPWR _19958_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_108_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR _23473_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__14701__A _15108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18909_ _17178_/X _18905_/X _19062_/A _18906_/X VGND VGND VPWR VPWR _24360_/D sky130_fd_sc_hd__o22a_4
X_19889_ _19884_/X _20644_/A _19888_/X VGND VGND VPWR VPWR _19889_/Y sky130_fd_sc_hd__o21ai_4
X_21920_ _21935_/A VGND VGND VPWR VPWR _21920_/X sky130_fd_sc_hd__buf_2
XANTENNA__13317__A _13317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12221__A _12496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21960__A2 _21959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18651__A2_N _18649_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21534__A _21249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21851_ _21850_/X _21841_/X _14535_/B _21848_/X VGND VGND VPWR VPWR _21851_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18169__B2 _18168_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16628__A _11782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20802_ _20802_/A _20801_/X VGND VGND VPWR VPWR _20802_/X sky130_fd_sc_hd__or2_4
XFILLER_97_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15532__A _14283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19905__A2 _24156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21782_ _21578_/X _21755_/A _23615_/Q _21737_/X VGND VGND VPWR VPWR _21782_/X sky130_fd_sc_hd__o22a_4
XFILLER_70_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16347__B _16279_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23521_ _23391_/CLK _23521_/D VGND VGND VPWR VPWR _15213_/B sky130_fd_sc_hd__dfxtp_4
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20733_ _20293_/X VGND VGND VPWR VPWR _20733_/X sky130_fd_sc_hd__buf_2
XFILLER_36_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20920__B1 HRDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14148__A _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13052__A _12496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20664_ _18430_/X _20653_/X _20516_/X _20663_/Y VGND VGND VPWR VPWR _20665_/A sky130_fd_sc_hd__a211o_4
X_23452_ _23293_/CLK _23452_/D VGND VGND VPWR VPWR _16559_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22365__A _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22403_ _20418_/A VGND VGND VPWR VPWR _22403_/X sky130_fd_sc_hd__buf_2
X_23383_ _23383_/CLK _23383_/D VGND VGND VPWR VPWR _16211_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17459__A _17688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21476__B2 _21474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20595_ _20595_/A _20595_/B VGND VGND VPWR VPWR _20595_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12891__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24094__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22334_ _22333_/X VGND VGND VPWR VPWR _22368_/A sky130_fd_sc_hd__buf_2
XFILLER_104_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21228__A1 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22265_ _22272_/A VGND VGND VPWR VPWR _22265_/X sky130_fd_sc_hd__buf_2
XANTENNA__21228__B2 _21218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21779__A2 _21776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21216_ _21271_/A VGND VGND VPWR VPWR _21242_/A sky130_fd_sc_hd__inv_2
X_24004_ _23363_/CLK _24004_/D VGND VGND VPWR VPWR _24004_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21709__A _21702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22196_ _22141_/X _22193_/X _15293_/B _22190_/X VGND VGND VPWR VPWR _23394_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20613__A _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21147_ _21118_/A VGND VGND VPWR VPWR _21147_/X sky130_fd_sc_hd__buf_2
XFILLER_117_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17194__A _13425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15707__A _15707_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17625__C _18274_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14611__A _11894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20332__B _20331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21078_ _20464_/X _21075_/X _12236_/B _21072_/X VGND VGND VPWR VPWR _21078_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14330__B _14330_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12920_ _12920_/A _12920_/B _12920_/C VGND VGND VPWR VPWR _12921_/C sky130_fd_sc_hd__and3_4
X_20029_ _20029_/A VGND VGND VPWR VPWR _20029_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13227__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21951__A2 _21945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12851_ _12851_/A _12928_/B VGND VGND VPWR VPWR _12851_/X sky130_fd_sc_hd__or2_4
XANTENNA__17641__B _17263_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11802_ _16231_/A VGND VGND VPWR VPWR _16677_/A sky130_fd_sc_hd__buf_2
XFILLER_27_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15442__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15570_ _14463_/A _15570_/B VGND VGND VPWR VPWR _15571_/C sky130_fd_sc_hd__or2_4
X_12782_ _13065_/A VGND VGND VPWR VPWR _15725_/A sky130_fd_sc_hd__buf_2
XANTENNA__24177__D _19750_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21703__A2 _21698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16257__B _23993_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14521_ _13699_/A _14518_/X _14520_/X VGND VGND VPWR VPWR _14521_/X sky130_fd_sc_hd__and3_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _16072_/A VGND VGND VPWR VPWR _11734_/A sky130_fd_sc_hd__buf_2
X_23719_ _23336_/CLK _21622_/X VGND VGND VPWR VPWR _23719_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14058__A _14046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _18249_/A VGND VGND VPWR VPWR _17240_/X sky130_fd_sc_hd__buf_2
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _12533_/A _14448_/X _14452_/C VGND VGND VPWR VPWR _14452_/X sky130_fd_sc_hd__or3_4
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A VGND VGND VPWR VPWR _12957_/A sky130_fd_sc_hd__buf_2
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _13351_/X _13403_/B _13402_/X VGND VGND VPWR VPWR _13403_/X sky130_fd_sc_hd__and3_4
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17171_ _14073_/X VGND VGND VPWR VPWR _17171_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13897__A _13890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383_ _15632_/A _14287_/B VGND VGND VPWR VPWR _14386_/B sky130_fd_sc_hd__or2_4
X_11595_ _11595_/A VGND VGND VPWR VPWR _11596_/A sky130_fd_sc_hd__buf_2
XFILLER_35_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16122_ _11982_/A _16122_/B VGND VGND VPWR VPWR _16122_/X sky130_fd_sc_hd__and2_4
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _13303_/X _13332_/X _13333_/X VGND VGND VPWR VPWR _13334_/X sky130_fd_sc_hd__and3_4
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16053_ _16019_/A _15981_/B VGND VGND VPWR VPWR _16053_/X sky130_fd_sc_hd__or2_4
X_13265_ _13243_/A _13263_/X _13264_/X VGND VGND VPWR VPWR _13265_/X sky130_fd_sc_hd__and3_4
XFILLER_100_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12306__A _15448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15004_ _15023_/A _15079_/B VGND VGND VPWR VPWR _15004_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12216_ _12216_/A VGND VGND VPWR VPWR _12217_/A sky130_fd_sc_hd__buf_2
XANTENNA__21619__A _21590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13196_ _15706_/A _13196_/B VGND VGND VPWR VPWR _13196_/X sky130_fd_sc_hd__or2_4
XFILLER_29_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20978__B1 _20977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19812_ _19603_/A _19643_/B _19812_/C VGND VGND VPWR VPWR _19812_/X sky130_fd_sc_hd__or3_4
XANTENNA_clkbuf_0_HCLK_A HCLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12147_ _11829_/A _23549_/Q VGND VGND VPWR VPWR _12147_/X sky130_fd_sc_hd__or2_4
XANTENNA__14521__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20242__B _20248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19743_ _19603_/A _19742_/X VGND VGND VPWR VPWR _19743_/X sky130_fd_sc_hd__or2_4
XANTENNA__15336__B _15277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12078_ _11997_/A _12140_/B VGND VGND VPWR VPWR _12079_/C sky130_fd_sc_hd__or2_4
X_16955_ _24121_/Q VGND VGND VPWR VPWR _16973_/A sky130_fd_sc_hd__inv_2
XANTENNA__22195__A2 _22193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19596__B1 HRDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13137__A _12221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15906_ _12672_/A _15890_/X _15906_/C VGND VGND VPWR VPWR _15907_/C sky130_fd_sc_hd__or3_4
XFILLER_110_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16886_ _16682_/X _16885_/X _16682_/X _16885_/X VGND VGND VPWR VPWR _16886_/X sky130_fd_sc_hd__a2bb2o_4
X_19674_ _19425_/Y VGND VGND VPWR VPWR _19674_/X sky130_fd_sc_hd__buf_2
XANTENNA__12041__A _11903_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15837_ _12890_/A _15835_/X _15836_/X VGND VGND VPWR VPWR _15837_/X sky130_fd_sc_hd__and3_4
X_18625_ _16935_/A _18613_/X _17006_/A _18624_/X VGND VGND VPWR VPWR _18625_/X sky130_fd_sc_hd__o22a_4
XFILLER_111_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16448__A _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15352__A _14810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15768_ _11680_/X _15768_/B _15767_/X VGND VGND VPWR VPWR _15768_/X sky130_fd_sc_hd__or3_4
X_18556_ _24190_/Q _16996_/A VGND VGND VPWR VPWR _18556_/X sky130_fd_sc_hd__or2_4
XFILLER_79_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14719_ _13918_/A _14719_/B _14718_/X VGND VGND VPWR VPWR _14719_/X sky130_fd_sc_hd__and3_4
X_17507_ _17504_/Y _17014_/X _17022_/A _17506_/X VGND VGND VPWR VPWR _17510_/B sky130_fd_sc_hd__o22a_4
X_18487_ _18486_/X VGND VGND VPWR VPWR _18487_/X sky130_fd_sc_hd__buf_2
X_15699_ _12738_/A _15699_/B VGND VGND VPWR VPWR _15699_/X sky130_fd_sc_hd__or2_4
XANTENNA__18571__B2 _18570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17438_ _17338_/X _17423_/Y _17430_/Y _17437_/Y VGND VGND VPWR VPWR _18153_/A sky130_fd_sc_hd__a211o_4
XANTENNA__15385__A1 _15185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23804__CLK _23840_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17369_ _17371_/B VGND VGND VPWR VPWR _18387_/B sky130_fd_sc_hd__inv_2
XANTENNA__17279__A _17277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21458__B2 _21453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22655__B1 _14308_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16183__A _16203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19520__B1 HRDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19108_ _19108_/A _19108_/B VGND VGND VPWR VPWR _19108_/X sky130_fd_sc_hd__and2_4
XANTENNA__13600__A _13600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20380_ _20380_/A _20258_/X VGND VGND VPWR VPWR _20380_/X sky130_fd_sc_hd__or2_4
XFILLER_118_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22913__A _23051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19039_ _19024_/X _19037_/Y _19038_/Y _19027_/X VGND VGND VPWR VPWR _19039_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16885__A1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22407__B1 _16158_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22050_ _21835_/X _22045_/X _23467_/Q _22049_/X VGND VGND VPWR VPWR _22050_/X sky130_fd_sc_hd__o22a_4
XFILLER_114_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18626__A2 _18606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21001_ _21001_/A VGND VGND VPWR VPWR _21293_/A sky130_fd_sc_hd__buf_2
XANTENNA__20433__A2 _20432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15527__A _12307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21630__B2 _21595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19334__A2_N _18378_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13047__A _13014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22952_ _22952_/A _22952_/B _22952_/C VGND VGND VPWR VPWR _22952_/X sky130_fd_sc_hd__and3_4
XANTENNA__24353__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21394__B1 _15180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21903_ _21843_/X _21901_/X _23560_/Q _21898_/X VGND VGND VPWR VPWR _21903_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19349__A2_N _18606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22883_ _22882_/X VGND VGND VPWR VPWR HADDR[0] sky130_fd_sc_hd__inv_2
XFILLER_3_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12886__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11790__A _11821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15262__A _14113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21834_ _21833_/X _21829_/X _23596_/Q _21824_/X VGND VGND VPWR VPWR _21834_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21697__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21765_ _21548_/X _21762_/X _15512_/B _21759_/X VGND VGND VPWR VPWR _23628_/D sky130_fd_sc_hd__o22a_4
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23504_ _24047_/CLK _21993_/X VGND VGND VPWR VPWR _23504_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22807__B _17109_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20716_ _18475_/X _20653_/X _20516_/X _20715_/Y VGND VGND VPWR VPWR _20717_/A sky130_fd_sc_hd__a211o_4
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21696_ _21514_/X _21691_/X _16472_/B _21695_/X VGND VGND VPWR VPWR _21696_/X sky130_fd_sc_hd__o22a_4
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20608__A _20534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22095__A _20486_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23435_ _23688_/CLK _22121_/X VGND VGND VPWR VPWR _23435_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20647_ HRDATA[14] _20699_/B VGND VGND VPWR VPWR _20647_/X sky130_fd_sc_hd__or2_4
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17117__A2 _17105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13510__A _12413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20578_ _20578_/A VGND VGND VPWR VPWR _20630_/A sky130_fd_sc_hd__buf_2
X_23366_ _23781_/CLK _22241_/X VGND VGND VPWR VPWR _14311_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_10_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22317_ _23309_/Q VGND VGND VPWR VPWR _22317_/X sky130_fd_sc_hd__buf_2
X_23297_ _23145_/CLK _22329_/X VGND VGND VPWR VPWR _15212_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13050_ _12512_/A _13120_/B VGND VGND VPWR VPWR _13051_/C sky130_fd_sc_hd__or2_4
X_22248_ _22145_/X _22243_/X _14898_/B _22212_/A VGND VGND VPWR VPWR _23360_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12001_ _11997_/A _23838_/Q VGND VGND VPWR VPWR _12002_/C sky130_fd_sc_hd__or2_4
XANTENNA__15437__A _13636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22179_ _22172_/A VGND VGND VPWR VPWR _22179_/X sky130_fd_sc_hd__buf_2
XANTENNA__21621__B2 _21616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12114__A1 _11992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22177__A2 _22172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16740_ _12112_/A _16740_/B _16740_/C VGND VGND VPWR VPWR _16741_/B sky130_fd_sc_hd__or3_4
X_13952_ _12216_/A _13952_/B _13951_/X VGND VGND VPWR VPWR _13956_/B sky130_fd_sc_hd__and3_4
XFILLER_4_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12903_ _12870_/A _12901_/X _12903_/C VGND VGND VPWR VPWR _12903_/X sky130_fd_sc_hd__and3_4
X_16671_ _16640_/X _16671_/B _16671_/C VGND VGND VPWR VPWR _16675_/B sky130_fd_sc_hd__and3_4
XFILLER_35_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13883_ _13700_/A _13883_/B _13883_/C VGND VGND VPWR VPWR _13884_/C sky130_fd_sc_hd__and3_4
XFILLER_62_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12796__A _12803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16268__A _11872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15622_ _15615_/A _15560_/B VGND VGND VPWR VPWR _15623_/C sky130_fd_sc_hd__or2_4
X_18410_ _17698_/X _18409_/X _17698_/X _18409_/X VGND VGND VPWR VPWR _18410_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15172__A _14725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12834_ _12769_/A _12832_/X _12833_/X VGND VGND VPWR VPWR _12838_/B sky130_fd_sc_hd__and3_4
X_19390_ _19389_/X _18316_/X _19389_/X _24208_/Q VGND VGND VPWR VPWR _19390_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18341_ _16977_/B VGND VGND VPWR VPWR _18341_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15553_ _15553_/A _23947_/Q VGND VGND VPWR VPWR _15553_/X sky130_fd_sc_hd__or2_4
X_12765_ _13097_/A VGND VGND VPWR VPWR _12765_/X sky130_fd_sc_hd__buf_2
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _13908_/A _14498_/X _14503_/X VGND VGND VPWR VPWR _14504_/X sky130_fd_sc_hd__or3_4
XFILLER_76_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19750__B1 _16677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _16025_/A VGND VGND VPWR VPWR _16072_/A sky130_fd_sc_hd__buf_2
X_18272_ _18392_/A _18271_/X VGND VGND VPWR VPWR _18272_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15900__A _13522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15484_/A _15476_/X _15484_/C VGND VGND VPWR VPWR _15484_/X sky130_fd_sc_hd__and3_4
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _15688_/A _12696_/B _12696_/C VGND VGND VPWR VPWR _12696_/X sky130_fd_sc_hd__or3_4
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17223_ _17130_/A VGND VGND VPWR VPWR _17826_/A sky130_fd_sc_hd__buf_2
XFILLER_50_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ _12441_/A _14501_/B VGND VGND VPWR VPWR _14435_/X sky130_fd_sc_hd__or2_4
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _11647_/A VGND VGND VPWR VPWR _12578_/A sky130_fd_sc_hd__buf_2
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17154_ _17135_/A VGND VGND VPWR VPWR _17154_/X sky130_fd_sc_hd__buf_2
X_14366_ _11766_/A VGND VGND VPWR VPWR _15628_/A sky130_fd_sc_hd__buf_2
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11578_ _16893_/A VGND VGND VPWR VPWR _16909_/B sky130_fd_sc_hd__buf_2
XANTENNA__22733__A SYSTICKCLKDIV[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16105_ _16130_/A _16098_/X _16105_/C VGND VGND VPWR VPWR _16105_/X sky130_fd_sc_hd__or3_4
X_13317_ _13317_/A VGND VGND VPWR VPWR _13483_/A sky130_fd_sc_hd__buf_2
X_17085_ _17084_/X VGND VGND VPWR VPWR _18048_/A sky130_fd_sc_hd__buf_2
X_14297_ _14322_/A _14295_/X _14297_/C VGND VGND VPWR VPWR _14298_/C sky130_fd_sc_hd__and3_4
XANTENNA__12036__A _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21860__B2 _21787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16036_ _11745_/X _16036_/B _16035_/X VGND VGND VPWR VPWR _16044_/B sky130_fd_sc_hd__or3_4
X_13248_ _13260_/A _13181_/B VGND VGND VPWR VPWR _13248_/X sky130_fd_sc_hd__or2_4
XFILLER_87_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16450__B _16383_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11875__A _16143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15347__A _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13179_ _12730_/A _13179_/B VGND VGND VPWR VPWR _13179_/X sky130_fd_sc_hd__or2_4
XFILLER_69_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17987_ _17961_/X _17965_/Y _17856_/X _17986_/Y VGND VGND VPWR VPWR _17987_/X sky130_fd_sc_hd__a211o_4
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22168__A2 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19569__B1 HRDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19726_ _19661_/A _19726_/B _19726_/C VGND VGND VPWR VPWR _19726_/X sky130_fd_sc_hd__or3_4
X_16938_ _17002_/A VGND VGND VPWR VPWR _17769_/A sky130_fd_sc_hd__inv_2
XANTENNA__20179__A1 _19884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19657_ _19524_/B _19872_/C _19722_/A _19656_/X VGND VGND VPWR VPWR _19657_/X sky130_fd_sc_hd__a211o_4
X_16869_ _14267_/B _16841_/X _14267_/B _16841_/X VGND VGND VPWR VPWR _16870_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18792__A1 _15911_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15082__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18608_ _17734_/A VGND VGND VPWR VPWR _18610_/A sky130_fd_sc_hd__buf_2
XFILLER_4_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19588_ _19553_/A HRDATA[11] VGND VGND VPWR VPWR _19588_/X sky130_fd_sc_hd__and2_4
XFILLER_20_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21812__A _21812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18539_ _18142_/A _17387_/X _18537_/Y _18398_/X _18538_/Y VGND VGND VPWR VPWR _18539_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22876__B1 _15910_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21679__B2 _21673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18544__A1 _18499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17347__A2 _17340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15810__A _12890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20887__C1 _20886_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21550_ _21265_/A VGND VGND VPWR VPWR _21550_/X sky130_fd_sc_hd__buf_2
XFILLER_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20501_ _20493_/X _20499_/X _19129_/A _20500_/X VGND VGND VPWR VPWR _20502_/B sky130_fd_sc_hd__o22a_4
X_21481_ _21467_/A VGND VGND VPWR VPWR _21481_/X sky130_fd_sc_hd__buf_2
XANTENNA__22628__B1 _16279_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14426__A _14336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20432_ _20293_/X _20431_/X _11528_/A _20303_/X VGND VGND VPWR VPWR _20432_/X sky130_fd_sc_hd__o22a_4
X_23220_ _24047_/CLK _23220_/D VGND VGND VPWR VPWR _23220_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22643__A _22636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20363_ _20251_/X _20362_/X _19231_/A _20327_/X VGND VGND VPWR VPWR _20363_/X sky130_fd_sc_hd__o22a_4
X_23151_ _24082_/CLK _23151_/D VGND VGND VPWR VPWR _13456_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17737__A _17737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21851__B2 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16641__A _16630_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_0_0_HCLK clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22102_ _22100_/X _22101_/X _23443_/Q _22096_/X VGND VGND VPWR VPWR _22102_/X sky130_fd_sc_hd__o22a_4
X_23082_ _23819_/CLK _23082_/D VGND VGND VPWR VPWR _23082_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21259__A _21247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20294_ _20257_/B VGND VGND VPWR VPWR _20556_/A sky130_fd_sc_hd__buf_2
X_22033_ _21807_/X _22031_/X _23479_/Q _22028_/X VGND VGND VPWR VPWR _22033_/X sky130_fd_sc_hd__o22a_4
XFILLER_103_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20406__A2 _20405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15257__A _11909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14161__A _14161_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21603__B2 _21602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23984_ _23157_/CLK _23984_/D VGND VGND VPWR VPWR _23984_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21906__A2 _21901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22935_ _22924_/X _18533_/A _22887_/X _22934_/X VGND VGND VPWR VPWR _22936_/A sky130_fd_sc_hd__a211o_4
XFILLER_84_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18783__A1 _17181_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13505__A _13500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22866_ _22872_/A _22866_/B VGND VGND VPWR VPWR HWDATA[26] sky130_fd_sc_hd__nor2_4
XANTENNA__24174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21817_ _21817_/A VGND VGND VPWR VPWR _21817_/X sky130_fd_sc_hd__buf_2
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22867__B1 _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22797_ _22821_/A VGND VGND VPWR VPWR _22807_/A sky130_fd_sc_hd__buf_2
XANTENNA__24103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12550_ _13031_/A _12657_/B VGND VGND VPWR VPWR _12550_/X sky130_fd_sc_hd__or2_4
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21748_ _21755_/A VGND VGND VPWR VPWR _21748_/X sky130_fd_sc_hd__buf_2
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20338__A _20338_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11501_ _24141_/Q VGND VGND VPWR VPWR _11625_/A sky130_fd_sc_hd__inv_2
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _12556_/A VGND VGND VPWR VPWR _12503_/A sky130_fd_sc_hd__buf_2
X_24467_ _24066_/CLK _24467_/D HRESETn VGND VGND VPWR VPWR _20010_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21679_ _21572_/X _21676_/X _15306_/B _21673_/X VGND VGND VPWR VPWR _21679_/X sky130_fd_sc_hd__o22a_4
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ _14345_/A _14217_/X _14220_/C VGND VGND VPWR VPWR _14220_/X sky130_fd_sc_hd__and3_4
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_16_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR _24230_/CLK sky130_fd_sc_hd__clkbuf_1
X_23418_ _23383_/CLK _22163_/X VGND VGND VPWR VPWR _16424_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24398_ _24334_/CLK _18844_/X HRESETn VGND VGND VPWR VPWR _24398_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17069__D _18866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_79_0_HCLK clkbuf_7_78_0_HCLK/A VGND VGND VPWR VPWR _23707_/CLK sky130_fd_sc_hd__clkbuf_1
X_14151_ _14151_/A VGND VGND VPWR VPWR _14152_/A sky130_fd_sc_hd__buf_2
X_23349_ _23987_/CLK _22270_/X VGND VGND VPWR VPWR _12580_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21842__B2 _21836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16551__A _11903_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13102_ _13102_/A _13093_/X _13102_/C VGND VGND VPWR VPWR _13103_/C sky130_fd_sc_hd__and3_4
XFILLER_101_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21169__A _21183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14082_ _15146_/A VGND VGND VPWR VPWR _14083_/A sky130_fd_sc_hd__buf_2
XANTENNA__23044__B1 _17766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20073__A _12100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13033_ _12917_/A _13031_/X _13033_/C VGND VGND VPWR VPWR _13034_/C sky130_fd_sc_hd__and3_4
X_17910_ _17244_/X VGND VGND VPWR VPWR _17910_/X sky130_fd_sc_hd__buf_2
XANTENNA__11695__A _13839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18890_ _12674_/X _18884_/X _24373_/Q _18885_/X VGND VGND VPWR VPWR _18890_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14071__A _14071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17841_ _17826_/X _17210_/X _17804_/A _17231_/X VGND VGND VPWR VPWR _17841_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14984_ _14202_/A _14984_/B _14984_/C VGND VGND VPWR VPWR _14985_/C sky130_fd_sc_hd__and3_4
X_17772_ _16927_/X _17637_/X _17639_/X _17771_/X VGND VGND VPWR VPWR _17772_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21358__B1 _23867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19511_ _19877_/B _19511_/B VGND VGND VPWR VPWR _19528_/C sky130_fd_sc_hd__or2_4
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13935_ _13951_/A VGND VGND VPWR VPWR _15037_/A sky130_fd_sc_hd__buf_2
X_16723_ _12083_/A _16791_/B VGND VGND VPWR VPWR _16725_/B sky130_fd_sc_hd__or2_4
XANTENNA__15614__B _23883_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13415__A _13415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16654_ _16617_/A _16654_/B VGND VGND VPWR VPWR _16654_/X sky130_fd_sc_hd__or2_4
X_19442_ _19485_/A _19442_/B VGND VGND VPWR VPWR _19450_/A sky130_fd_sc_hd__or2_4
XFILLER_90_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13866_ _11670_/A _13854_/X _13865_/X VGND VGND VPWR VPWR _13886_/B sky130_fd_sc_hd__and3_4
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20581__B2 _20497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22728__A SYSTICKCLKDIV[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15605_ _15617_/A _23659_/Q VGND VGND VPWR VPWR _15607_/B sky130_fd_sc_hd__or2_4
X_12817_ _12754_/X _12815_/X _12817_/C VGND VGND VPWR VPWR _12821_/B sky130_fd_sc_hd__and3_4
X_16585_ _16542_/A _16581_/X _16584_/X VGND VGND VPWR VPWR _16585_/X sky130_fd_sc_hd__or3_4
X_19373_ _19370_/X _18061_/Y _19370_/X _24216_/Q VGND VGND VPWR VPWR _24216_/D sky130_fd_sc_hd__a2bb2o_4
X_13797_ _15435_/A _13793_/X _13796_/X VGND VGND VPWR VPWR _13797_/X sky130_fd_sc_hd__or3_4
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15536_ _15536_/A _23659_/Q VGND VGND VPWR VPWR _15536_/X sky130_fd_sc_hd__or2_4
X_18324_ _17861_/A _18323_/X _17836_/A _17255_/X VGND VGND VPWR VPWR _18324_/X sky130_fd_sc_hd__o22a_4
XFILLER_91_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12748_ _13004_/A _12748_/B _12747_/X VGND VGND VPWR VPWR _12748_/X sky130_fd_sc_hd__or3_4
XFILLER_37_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20333__A1 _17880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21530__B1 _12774_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20248__A _20248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16445__B _16380_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18255_ _18254_/A _18254_/B _18048_/X VGND VGND VPWR VPWR _18255_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_72_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15467_ _12646_/A _15465_/X _15466_/X VGND VGND VPWR VPWR _15468_/C sky130_fd_sc_hd__and3_4
X_12679_ _12559_/X _12676_/X _12678_/Y VGND VGND VPWR VPWR _12680_/B sky130_fd_sc_hd__a21o_4
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14246__A _14246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18941__A _18994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17206_ _13278_/X _17161_/X _17192_/Y _17157_/X VGND VGND VPWR VPWR _17206_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14418_ _13845_/A _14324_/B VGND VGND VPWR VPWR _14419_/C sky130_fd_sc_hd__or2_4
X_18186_ _18040_/X _18073_/X _17868_/X VGND VGND VPWR VPWR _18186_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_15_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15398_ _15398_/A _15394_/X _15398_/C VGND VGND VPWR VPWR _15398_/X sky130_fd_sc_hd__or3_4
XFILLER_15_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24155__CLK _24162_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17137_ _17161_/A VGND VGND VPWR VPWR _17137_/X sky130_fd_sc_hd__buf_2
X_14349_ _15615_/A _14272_/B VGND VGND VPWR VPWR _14350_/C sky130_fd_sc_hd__or2_4
XFILLER_116_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17068_ _17068_/A VGND VGND VPWR VPWR _17068_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21079__A _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16019_ _16019_/A _16019_/B VGND VGND VPWR VPWR _16021_/B sky130_fd_sc_hd__or2_4
XANTENNA__15077__A _15115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21807__A _20442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18388__A _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12213__B _12213_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15805__A _12850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19709_ _19419_/X _19708_/X _12096_/A _19678_/X VGND VGND VPWR VPWR _19709_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22010__A1 _21852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22010__B2 _22006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20981_ _22460_/A VGND VGND VPWR VPWR _21291_/A sky130_fd_sc_hd__buf_2
XANTENNA__22561__A2 _22557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22720_ _22719_/X VGND VGND VPWR VPWR _22898_/A sky130_fd_sc_hd__buf_2
X_22651_ _22439_/X _22650_/X _23113_/Q _22647_/X VGND VGND VPWR VPWR _23113_/D sky130_fd_sc_hd__o22a_4
XFILLER_0_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19714__B1 _19784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21602_ _21602_/A VGND VGND VPWR VPWR _21602_/X sky130_fd_sc_hd__buf_2
X_22582_ _22408_/X _22579_/X _12274_/B _22576_/X VGND VGND VPWR VPWR _22582_/X sky130_fd_sc_hd__o22a_4
X_24321_ _24321_/CLK _24321_/D HRESETn VGND VGND VPWR VPWR _11503_/A sky130_fd_sc_hd__dfstp_4
X_21533_ _21531_/X _21532_/X _12858_/B _21527_/X VGND VGND VPWR VPWR _23763_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17740__A2 _17122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24252_ _24250_/CLK _24252_/D HRESETn VGND VGND VPWR VPWR _24252_/Q sky130_fd_sc_hd__dfrtp_4
X_21464_ _21234_/X _21463_/X _23800_/Q _21460_/X VGND VGND VPWR VPWR _23800_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23203_ _23433_/CLK _22509_/X VGND VGND VPWR VPWR _14772_/B sky130_fd_sc_hd__dfxtp_4
X_20415_ _20209_/X _20401_/Y _20413_/X _20414_/Y _20233_/X VGND VGND VPWR VPWR _20415_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13995__A _14841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17467__A _11924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21395_ _21291_/X _21390_/X _23840_/Q _21359_/A VGND VGND VPWR VPWR _23840_/D sky130_fd_sc_hd__o22a_4
X_24183_ _24187_/CLK _19652_/Y HRESETn VGND VGND VPWR VPWR _17552_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23134_ _23326_/CLK _22620_/X VGND VGND VPWR VPWR _11810_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20346_ _20251_/X _20345_/X _19232_/A _20327_/X VGND VGND VPWR VPWR _20346_/X sky130_fd_sc_hd__o22a_4
XFILLER_49_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20277_ _21789_/A VGND VGND VPWR VPWR _20277_/X sky130_fd_sc_hd__buf_2
X_23065_ _18605_/X _19955_/X _19956_/A _18605_/X VGND VGND VPWR VPWR _24478_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22016_ _23486_/Q VGND VGND VPWR VPWR _22016_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21052__A2 _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18298__A _18244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12123__B _12123_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15715__A _13130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22001__B2 _21999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11981_ _11980_/X VGND VGND VPWR VPWR _11982_/A sky130_fd_sc_hd__buf_2
X_23967_ _23130_/CLK _21160_/X VGND VGND VPWR VPWR _15079_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13720_ _15495_/A _13720_/B _13719_/X VGND VGND VPWR VPWR _13721_/C sky130_fd_sc_hd__and3_4
XANTENNA__13235__A _13211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22552__A2 _22550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22918_ _22886_/X _17724_/X _22887_/X _22917_/X VGND VGND VPWR VPWR _22919_/A sky130_fd_sc_hd__a211o_4
XFILLER_95_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20563__A1 _20468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23898_ _23706_/CLK _21310_/X VGND VGND VPWR VPWR _16413_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20563__B2 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21452__A _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13651_ _13651_/A _13651_/B VGND VGND VPWR VPWR _13651_/X sky130_fd_sc_hd__or2_4
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22849_ _22849_/A VGND VGND VPWR VPWR HWDATA[22] sky130_fd_sc_hd__inv_2
XFILLER_71_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12602_ _13726_/A VGND VGND VPWR VPWR _12650_/A sky130_fd_sc_hd__buf_2
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15450__A _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16370_ _16363_/X _16366_/X _16370_/C VGND VGND VPWR VPWR _16371_/C sky130_fd_sc_hd__or3_4
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13582_ _13136_/X _13273_/Y _13277_/A _13581_/Y VGND VGND VPWR VPWR _13582_/X sky130_fd_sc_hd__a211o_4
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12793__B _23156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15321_ _11638_/A _15321_/B _15320_/X VGND VGND VPWR VPWR _15331_/B sky130_fd_sc_hd__or3_4
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12533_ _12533_/A VGND VGND VPWR VPWR _13041_/A sky130_fd_sc_hd__buf_2
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14066__A _11647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18761__A _11844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18040_ _17861_/A VGND VGND VPWR VPWR _18040_/X sky130_fd_sc_hd__buf_2
X_15252_ _11879_/A _15252_/B VGND VGND VPWR VPWR _15254_/B sky130_fd_sc_hd__or2_4
X_12464_ _12464_/A _12462_/X _12463_/X VGND VGND VPWR VPWR _12464_/X sky130_fd_sc_hd__and3_4
XFILLER_12_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22283__A _22269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ _11738_/A VGND VGND VPWR VPWR _14367_/A sky130_fd_sc_hd__buf_2
XANTENNA__17377__A _15909_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15183_ _14172_/A _15183_/B VGND VGND VPWR VPWR _15183_/X sky130_fd_sc_hd__and2_4
XANTENNA__21815__B2 _21812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12395_ _15743_/A _12393_/X _12395_/C VGND VGND VPWR VPWR _12399_/B sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_4_11_0_HCLK_A clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14134_ _14318_/A _24041_/Q VGND VGND VPWR VPWR _14134_/X sky130_fd_sc_hd__or2_4
XFILLER_67_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19991_ _18127_/X _19985_/X _19990_/Y _19972_/X VGND VGND VPWR VPWR _19991_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15609__B _23531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14065_ _14065_/A _14063_/X _14065_/C VGND VGND VPWR VPWR _14070_/B sky130_fd_sc_hd__and3_4
X_18942_ _11532_/X VGND VGND VPWR VPWR _18942_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19592__A _19592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_9_0_HCLK clkbuf_6_4_0_HCLK/X VGND VGND VPWR VPWR _23522_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21579__B1 _23743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13016_ _13016_/A _23538_/Q VGND VGND VPWR VPWR _13017_/C sky130_fd_sc_hd__or2_4
XANTENNA__21043__A2 _21037_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18873_ _18873_/A VGND VGND VPWR VPWR _18898_/A sky130_fd_sc_hd__buf_2
XFILLER_80_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17824_ _17824_/A VGND VGND VPWR VPWR _17824_/X sky130_fd_sc_hd__buf_2
XFILLER_94_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14967_ _14925_/A _14965_/X _14966_/X VGND VGND VPWR VPWR _14967_/X sky130_fd_sc_hd__and3_4
X_17755_ _17755_/A _17755_/B VGND VGND VPWR VPWR _17755_/X sky130_fd_sc_hd__or2_4
XANTENNA__13145__A _12240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16706_ _12025_/A _16706_/B _16706_/C VGND VGND VPWR VPWR _16710_/B sky130_fd_sc_hd__and3_4
X_13918_ _13918_/A _13886_/X _13918_/C VGND VGND VPWR VPWR _13918_/X sky130_fd_sc_hd__and3_4
XANTENNA__20554__A1 _20511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14898_ _14895_/A _14898_/B VGND VGND VPWR VPWR _14898_/X sky130_fd_sc_hd__or2_4
X_17686_ _17685_/Y _17667_/X _17665_/A VGND VGND VPWR VPWR _17686_/X sky130_fd_sc_hd__a21o_4
XANTENNA__22458__A _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20554__B2 _20488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19425_ _19416_/B VGND VGND VPWR VPWR _19425_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21362__A _21369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13849_ _11707_/A VGND VGND VPWR VPWR _15314_/A sky130_fd_sc_hd__buf_2
X_16637_ _16662_/A _23676_/Q VGND VGND VPWR VPWR _16637_/X sky130_fd_sc_hd__or2_4
XFILLER_62_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12984__A _12622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16456__A _11715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17970__A2 _17828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15360__A _14009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19356_ _19356_/A VGND VGND VPWR VPWR _19356_/Y sky130_fd_sc_hd__inv_2
X_16568_ _16565_/A _24060_/Q VGND VGND VPWR VPWR _16569_/C sky130_fd_sc_hd__or2_4
XFILLER_50_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18307_ _18307_/A _18307_/B VGND VGND VPWR VPWR _18307_/X sky130_fd_sc_hd__or2_4
XFILLER_17_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15519_ _15453_/Y _15517_/X VGND VGND VPWR VPWR _15519_/X sky130_fd_sc_hd__or2_4
X_16499_ _16499_/A _16497_/X _16499_/C VGND VGND VPWR VPWR _16499_/X sky130_fd_sc_hd__and3_4
X_19287_ _19209_/X VGND VGND VPWR VPWR _19287_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17183__B1 _17182_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18238_ _22998_/B _18237_/Y _17667_/A _18237_/A VGND VGND VPWR VPWR _18238_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22193__A _22153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18169_ _18009_/X _18163_/X _18053_/X _18168_/X VGND VGND VPWR VPWR _18169_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16191__A _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21806__B2 _21800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_62_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR _23922_/CLK sky130_fd_sc_hd__clkbuf_1
X_20200_ _20199_/X VGND VGND VPWR VPWR _20279_/A sky130_fd_sc_hd__buf_2
XANTENNA__17486__A1 _11834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21180_ _21180_/A VGND VGND VPWR VPWR _21180_/X sky130_fd_sc_hd__buf_2
XANTENNA__15519__B _15517_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22921__A _23027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20131_ _19884_/X _18610_/A _20130_/X VGND VGND VPWR VPWR _20131_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_28_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12224__A _12691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20062_ _24456_/Q VGND VGND VPWR VPWR _20062_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17734__B _17111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22231__B2 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20441__A _20441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23821_ _23922_/CLK _21428_/X VGND VGND VPWR VPWR _23821_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_113_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18738__A1 _18735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22534__A2 _22529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13055__A _13055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23752_ _23304_/CLK _23752_/D VGND VGND VPWR VPWR _13713_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_66_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20964_ _20214_/Y _20962_/X _20963_/X VGND VGND VPWR VPWR _20964_/X sky130_fd_sc_hd__a21o_4
XFILLER_81_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22368__A _22368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21742__B1 _23645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22703_ _20819_/A _22700_/X _23079_/Q _22697_/X VGND VGND VPWR VPWR _22703_/X sky130_fd_sc_hd__o22a_4
X_23683_ _23270_/CLK _21678_/X VGND VGND VPWR VPWR _14779_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12894__A _12462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20895_ _20846_/B _20895_/B VGND VGND VPWR VPWR _20895_/X sky130_fd_sc_hd__or2_4
XANTENNA__16366__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15270__A _14161_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22634_ _22410_/X _22629_/X _12647_/B _22633_/X VGND VGND VPWR VPWR _22634_/X sky130_fd_sc_hd__o22a_4
XFILLER_74_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22298__B2 _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22565_ _21581_/A _21917_/B _21297_/A _21060_/A VGND VGND VPWR VPWR _22566_/A sky130_fd_sc_hd__or4_4
XANTENNA__17174__B1 _12992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18910__A1 _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24304_ _23260_/CLK _19168_/X HRESETn VGND VGND VPWR VPWR _24304_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22815__B _17298_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21516_ _21514_/X _21508_/X _16388_/B _21515_/X VGND VGND VPWR VPWR _23770_/D sky130_fd_sc_hd__o22a_4
X_22496_ _22432_/X _22493_/X _15511_/B _22490_/X VGND VGND VPWR VPWR _23212_/D sky130_fd_sc_hd__o22a_4
X_24235_ _24208_/CLK _24235_/D HRESETn VGND VGND VPWR VPWR _24235_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21447_ _23806_/Q VGND VGND VPWR VPWR _21447_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14614__A _14725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12180_ _11747_/X _12176_/X _12179_/X VGND VGND VPWR VPWR _12180_/X sky130_fd_sc_hd__or3_4
X_24166_ _23584_/CLK _19850_/Y HRESETn VGND VGND VPWR VPWR _22017_/A sky130_fd_sc_hd__dfrtp_4
X_21378_ _21261_/X _21376_/X _15839_/B _21373_/X VGND VGND VPWR VPWR _21378_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22470__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23117_ _23564_/CLK _22645_/X VGND VGND VPWR VPWR _15821_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_46_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20329_ _20322_/X _20328_/X _24348_/Q _20247_/X VGND VGND VPWR VPWR _20329_/X sky130_fd_sc_hd__o22a_4
X_24097_ _24290_/CLK _24097_/D HRESETn VGND VGND VPWR VPWR _24097_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12134__A _11746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17229__A1 _16814_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23048_ _23048_/A _23046_/X _23048_/C VGND VGND VPWR VPWR _23048_/X sky130_fd_sc_hd__and3_4
XFILLER_62_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17644__B _17535_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11973__A _12112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15870_ _13551_/X _23309_/Q VGND VGND VPWR VPWR _15870_/X sky130_fd_sc_hd__or2_4
XFILLER_114_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12788__B _23924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14821_ _13710_/A _14821_/B _14821_/C VGND VGND VPWR VPWR _14821_/X sky130_fd_sc_hd__and3_4
XFILLER_92_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22525__A2 _22522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14752_ _14752_/A _14748_/X _14752_/C VGND VGND VPWR VPWR _14752_/X sky130_fd_sc_hd__or3_4
X_17540_ _17540_/A _17957_/B VGND VGND VPWR VPWR _17627_/A sky130_fd_sc_hd__or2_4
X_11964_ _11997_/A _21110_/A VGND VGND VPWR VPWR _11965_/C sky130_fd_sc_hd__or2_4
XFILLER_91_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13703_ _15487_/A _13703_/B VGND VGND VPWR VPWR _13704_/C sky130_fd_sc_hd__or2_4
X_17471_ _12676_/X _17527_/B VGND VGND VPWR VPWR _17471_/X sky130_fd_sc_hd__or2_4
XFILLER_75_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14683_ _14714_/A _14683_/B VGND VGND VPWR VPWR _14683_/X sky130_fd_sc_hd__or2_4
X_11895_ _15393_/A VGND VGND VPWR VPWR _14463_/A sky130_fd_sc_hd__buf_2
X_19210_ _24261_/Q _19209_/X VGND VGND VPWR VPWR _19211_/B sky130_fd_sc_hd__and2_4
XFILLER_72_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23568__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15180__A _14151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13634_ _15436_/A _23304_/Q VGND VGND VPWR VPWR _13634_/X sky130_fd_sc_hd__or2_4
X_16422_ _16083_/A _16420_/X _16421_/X VGND VGND VPWR VPWR _16422_/X sky130_fd_sc_hd__and3_4
XFILLER_73_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22289__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22289__B2 _22283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16353_ _13415_/A _16349_/X _16353_/C VGND VGND VPWR VPWR _16353_/X sky130_fd_sc_hd__or3_4
X_19141_ _19139_/A _19138_/X _20244_/A _19140_/Y VGND VGND VPWR VPWR _24318_/D sky130_fd_sc_hd__o22a_4
X_13565_ _13551_/X _23471_/Q VGND VGND VPWR VPWR _13565_/X sky130_fd_sc_hd__or2_4
XANTENNA__19587__A HRDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18901__A1 _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15304_ _15030_/A _15304_/B VGND VGND VPWR VPWR _15305_/C sky130_fd_sc_hd__or2_4
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12516_ _12892_/A _12516_/B VGND VGND VPWR VPWR _12516_/X sky130_fd_sc_hd__and2_4
X_19072_ _19072_/A VGND VGND VPWR VPWR _19072_/Y sky130_fd_sc_hd__inv_2
X_16284_ _16151_/A _16282_/X _16284_/C VGND VGND VPWR VPWR _16285_/C sky130_fd_sc_hd__and3_4
X_13496_ _15876_/A _13427_/B VGND VGND VPWR VPWR _13496_/X sky130_fd_sc_hd__or2_4
XANTENNA__16912__B1 _16907_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16723__B _16791_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15235_ _14215_/A _15235_/B _15234_/X VGND VGND VPWR VPWR _15235_/X sky130_fd_sc_hd__and3_4
X_18023_ _18498_/A VGND VGND VPWR VPWR _18239_/A sky130_fd_sc_hd__buf_2
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12447_ _15045_/A VGND VGND VPWR VPWR _14748_/A sky130_fd_sc_hd__buf_2
Xclkbuf_6_49_0_HCLK clkbuf_6_49_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_49_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15166_ _14575_/X _15166_/B VGND VGND VPWR VPWR _15166_/X sky130_fd_sc_hd__or2_4
XANTENNA__21264__A2 _21259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12378_ _13908_/A VGND VGND VPWR VPWR _13211_/A sky130_fd_sc_hd__buf_2
XANTENNA__22461__B2 _22386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14117_ _14117_/A _14113_/X _14117_/C VGND VGND VPWR VPWR _14117_/X sky130_fd_sc_hd__and3_4
XFILLER_113_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15097_ _15109_/A _15097_/B VGND VGND VPWR VPWR _15099_/B sky130_fd_sc_hd__or2_4
X_19974_ _19970_/X _17766_/A _19934_/X _19973_/X VGND VGND VPWR VPWR _19974_/X sky130_fd_sc_hd__o22a_4
XFILLER_99_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14048_ _14813_/A _13966_/B VGND VGND VPWR VPWR _14048_/X sky130_fd_sc_hd__or2_4
X_18925_ _24348_/Q VGND VGND VPWR VPWR _18926_/C sky130_fd_sc_hd__inv_2
XANTENNA__12979__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11883__A _15784_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18856_ _18842_/A VGND VGND VPWR VPWR _18856_/X sky130_fd_sc_hd__buf_2
XANTENNA__20775__A1 _24233_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17807_ _17806_/X VGND VGND VPWR VPWR _17807_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16443__A2 _11618_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17640__B2 _17044_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0_HCLK clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18787_ _17194_/X _18781_/X _24432_/Q _18782_/X VGND VGND VPWR VPWR _24432_/D sky130_fd_sc_hd__o22a_4
X_15999_ _13448_/X VGND VGND VPWR VPWR _15999_/X sky130_fd_sc_hd__buf_2
XFILLER_36_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17738_ _17738_/A VGND VGND VPWR VPWR _17738_/X sky130_fd_sc_hd__buf_2
XFILLER_35_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21724__B1 _14283_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19393__B2 _24206_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15802__B _15802_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17669_ _17665_/X _17668_/Y VGND VGND VPWR VPWR _17669_/X sky130_fd_sc_hd__or2_4
XANTENNA__16186__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19408_ _19406_/X _18665_/X _19406_/X _24195_/Q VGND VGND VPWR VPWR _24195_/D sky130_fd_sc_hd__a2bb2o_4
X_20680_ _20447_/A VGND VGND VPWR VPWR _20680_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22916__A _18624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19339_ _19336_/X _18455_/X _19336_/X _24236_/Q VGND VGND VPWR VPWR _19339_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16914__A _16907_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22350_ _22093_/X _22347_/X _12241_/B _22344_/X VGND VGND VPWR VPWR _23286_/D sky130_fd_sc_hd__o22a_4
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17729__B _17106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21301_ _21316_/A VGND VGND VPWR VPWR _21301_/X sky130_fd_sc_hd__buf_2
X_22281_ _22115_/X _22279_/X _15848_/B _22276_/X VGND VGND VPWR VPWR _22281_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24020_ _24021_/CLK _21081_/X VGND VGND VPWR VPWR _24020_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21232_ _21802_/A VGND VGND VPWR VPWR _21232_/X sky130_fd_sc_hd__buf_2
XANTENNA__21255__A2 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21163_ _21162_/X VGND VGND VPWR VPWR _21168_/A sky130_fd_sc_hd__buf_2
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20114_ _11558_/A _20112_/Y _20113_/Y VGND VGND VPWR VPWR _20114_/X sky130_fd_sc_hd__o21a_4
X_21094_ _20723_/X _21089_/X _24011_/Q _21093_/X VGND VGND VPWR VPWR _21094_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12889__A _13029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20045_ _18456_/X _20033_/X _20043_/Y _20044_/X VGND VGND VPWR VPWR _20045_/X sky130_fd_sc_hd__o22a_4
XFILLER_86_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15265__A _14136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20766__B2 _20562_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21963__B1 _15213_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23804_ _23840_/CLK _23804_/D VGND VGND VPWR VPWR _23804_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21996_ _21828_/X _21995_/X _15715_/B _21992_/X VGND VGND VPWR VPWR _23502_/D sky130_fd_sc_hd__o22a_4
XFILLER_54_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22098__A _22413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _24088_/CLK _23735_/D VGND VGND VPWR VPWR _23735_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _20255_/A _20946_/X _19098_/A _18870_/X VGND VGND VPWR VPWR _20947_/X sky130_fd_sc_hd__o22a_4
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21191__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _12626_/A VGND VGND VPWR VPWR _11680_/X sky130_fd_sc_hd__buf_2
X_23666_ _23314_/CLK _21707_/X VGND VGND VPWR VPWR _23666_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ HRDATA[5] VGND VGND VPWR VPWR _20878_/Y sky130_fd_sc_hd__inv_2
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22617_ _22621_/A VGND VGND VPWR VPWR _22633_/A sky130_fd_sc_hd__inv_2
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23597_ _23826_/CLK _21832_/X VGND VGND VPWR VPWR _15879_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13350_ _13349_/X VGND VGND VPWR VPWR _13350_/Y sky130_fd_sc_hd__inv_2
X_22548_ _22434_/X _22543_/X _23179_/Q _22547_/X VGND VGND VPWR VPWR _23179_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21494__A2 _21491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22691__B2 _22690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12301_ _12301_/A VGND VGND VPWR VPWR _12302_/A sky130_fd_sc_hd__buf_2
XANTENNA__11968__A _12022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13281_ _15654_/A VGND VGND VPWR VPWR _13281_/X sky130_fd_sc_hd__buf_2
X_22479_ _22486_/A VGND VGND VPWR VPWR _22479_/X sky130_fd_sc_hd__buf_2
XANTENNA__14344__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15020_ _14165_/A _15088_/B VGND VGND VPWR VPWR _15021_/C sky130_fd_sc_hd__or2_4
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12232_ _12202_/A VGND VGND VPWR VPWR _13678_/A sky130_fd_sc_hd__buf_2
X_24218_ _24216_/CLK _24218_/D HRESETn VGND VGND VPWR VPWR _24218_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22443__B2 _22435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_3_0_HCLK_A clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12163_ _11734_/A _23421_/Q VGND VGND VPWR VPWR _12163_/X sky130_fd_sc_hd__or2_4
X_24149_ _24223_/CLK _24149_/D HRESETn VGND VGND VPWR VPWR _24149_/Q sky130_fd_sc_hd__dfrtp_4
X_12094_ _12065_/X _23421_/Q VGND VGND VPWR VPWR _12095_/C sky130_fd_sc_hd__or2_4
X_16971_ _17708_/A _16971_/B VGND VGND VPWR VPWR _16972_/B sky130_fd_sc_hd__or2_4
XFILLER_42_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18710_ _18011_/X _16997_/X _18556_/X VGND VGND VPWR VPWR _18710_/X sky130_fd_sc_hd__o21a_4
XFILLER_104_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15175__A _14146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15922_ _15909_/X VGND VGND VPWR VPWR _15922_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19690_ _19817_/C _19689_/Y _19877_/B VGND VGND VPWR VPWR _19690_/X sky130_fd_sc_hd__and3_4
XFILLER_81_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18641_ _18640_/X VGND VGND VPWR VPWR _18641_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21905__A _21884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15853_ _12386_/X _15792_/B VGND VGND VPWR VPWR _15853_/X sky130_fd_sc_hd__or2_4
XFILLER_40_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18486__A _17634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14804_ _12575_/A _14802_/X _14803_/X VGND VGND VPWR VPWR _14804_/X sky130_fd_sc_hd__and3_4
XFILLER_76_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15903__A _13511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18572_ _17746_/X _17747_/B _17746_/X _17747_/B VGND VGND VPWR VPWR _18572_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12996_ _12845_/X _12996_/B VGND VGND VPWR VPWR _12996_/X sky130_fd_sc_hd__or2_4
X_15784_ _15784_/A _15845_/B VGND VGND VPWR VPWR _15784_/X sky130_fd_sc_hd__or2_4
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17523_ _17461_/B VGND VGND VPWR VPWR _17523_/Y sky130_fd_sc_hd__inv_2
X_11947_ _11999_/A _11947_/B _11947_/C VGND VGND VPWR VPWR _11947_/X sky130_fd_sc_hd__or3_4
X_14735_ _14758_/A _14797_/B VGND VGND VPWR VPWR _14737_/B sky130_fd_sc_hd__or2_4
XANTENNA__15622__B _15560_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14519__A _13879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21182__B2 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13423__A _12787_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14666_ _14252_/A VGND VGND VPWR VPWR _14666_/X sky130_fd_sc_hd__buf_2
X_17454_ _17454_/A VGND VGND VPWR VPWR _17455_/B sky130_fd_sc_hd__inv_2
XFILLER_18_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11878_ _15146_/A VGND VGND VPWR VPWR _11879_/A sky130_fd_sc_hd__buf_2
XANTENNA__22736__A SYSTICKCLKDIV[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13617_ _15435_/A _13609_/X _13616_/X VGND VGND VPWR VPWR _13617_/X sky130_fd_sc_hd__or3_4
X_16405_ _13477_/X _16405_/B VGND VGND VPWR VPWR _16406_/C sky130_fd_sc_hd__or2_4
XANTENNA__21640__A _21636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_24_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14597_ _13600_/A _14592_/X _14597_/C VGND VGND VPWR VPWR _14597_/X sky130_fd_sc_hd__or3_4
X_17385_ _17384_/Y _17413_/B VGND VGND VPWR VPWR _17385_/X sky130_fd_sc_hd__or2_4
XANTENNA__16734__A _11993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12039__A _11888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19124_ _24303_/Q _19124_/B VGND VGND VPWR VPWR _19169_/A sky130_fd_sc_hd__and2_4
XFILLER_13_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13548_ _12959_/A VGND VGND VPWR VPWR _13548_/X sky130_fd_sc_hd__buf_2
X_16336_ _11727_/X _16336_/B _16336_/C VGND VGND VPWR VPWR _16337_/C sky130_fd_sc_hd__and3_4
XANTENNA__21485__A2 _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22682__A1 _20464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22682__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11878__A _15146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16267_ _11959_/X _16267_/B VGND VGND VPWR VPWR _16267_/X sky130_fd_sc_hd__or2_4
X_19055_ _19053_/Y _19054_/Y _11515_/B VGND VGND VPWR VPWR _19055_/X sky130_fd_sc_hd__o21a_4
XFILLER_16_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13479_ _13447_/X _13479_/B _13478_/X VGND VGND VPWR VPWR _13483_/B sky130_fd_sc_hd__and3_4
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14254__A _13839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15218_ _14644_/A _23873_/Q VGND VGND VPWR VPWR _15220_/B sky130_fd_sc_hd__or2_4
X_18006_ _16927_/X _18001_/X _17639_/X _18005_/X VGND VGND VPWR VPWR _18006_/X sky130_fd_sc_hd__o22a_4
XFILLER_86_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16198_ _16198_/A _16198_/B _16197_/X VGND VGND VPWR VPWR _16199_/C sky130_fd_sc_hd__or3_4
XANTENNA__15069__B _23903_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22471__A _22471_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15149_ _14121_/A _15149_/B VGND VGND VPWR VPWR _15149_/X sky130_fd_sc_hd__or2_4
XFILLER_86_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20996__A1 _18752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19957_ _19929_/X VGND VGND VPWR VPWR _19957_/X sky130_fd_sc_hd__buf_2
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22198__B1 _14899_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18908_ _14261_/X _18905_/X _24361_/Q _18906_/X VGND VGND VPWR VPWR _18908_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15085__A _14055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19888_ _19933_/A _19887_/X VGND VGND VPWR VPWR _19888_/X sky130_fd_sc_hd__or2_4
XFILLER_25_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12502__A _12540_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18839_ _13270_/X _18834_/X _24401_/Q _18835_/X VGND VGND VPWR VPWR _24401_/D sky130_fd_sc_hd__o22a_4
XFILLER_3_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21850_ _20870_/A VGND VGND VPWR VPWR _21850_/X sky130_fd_sc_hd__buf_2
XFILLER_97_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20801_ _20641_/X _20799_/X _20800_/X VGND VGND VPWR VPWR _20801_/X sky130_fd_sc_hd__and3_4
XFILLER_70_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15532__B _24011_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21781_ _21576_/X _21776_/X _23616_/Q _21737_/X VGND VGND VPWR VPWR _21781_/X sky130_fd_sc_hd__o22a_4
XFILLER_58_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14429__A _14336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23520_ _23391_/CLK _23520_/D VGND VGND VPWR VPWR _23520_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13333__A _13428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20732_ _20292_/X VGND VGND VPWR VPWR _20732_/X sky130_fd_sc_hd__buf_2
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23451_ _23293_/CLK _23451_/D VGND VGND VPWR VPWR _16708_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20663_ _20603_/A _20663_/B VGND VGND VPWR VPWR _20663_/Y sky130_fd_sc_hd__nor2_4
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16644__A _16599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23113__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22402_ _22401_/X _22392_/X _16240_/B _22399_/X VGND VGND VPWR VPWR _23257_/D sky130_fd_sc_hd__o22a_4
XFILLER_91_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23382_ _23473_/CLK _22218_/X VGND VGND VPWR VPWR _12297_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21476__A2 _21470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22673__A1 _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20594_ _20422_/X _19770_/X _20286_/A VGND VGND VPWR VPWR _20594_/X sky130_fd_sc_hd__a21o_4
XANTENNA__22673__B2 _22669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22333_ _22068_/A _21634_/B _21297_/A _21008_/A VGND VGND VPWR VPWR _22333_/X sky130_fd_sc_hd__or4_4
XANTENNA__11788__A _12169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14164__A _14992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24376__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24199__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22264_ _22086_/X _22258_/X _16244_/B _22262_/X VGND VGND VPWR VPWR _23353_/D sky130_fd_sc_hd__o22a_4
XFILLER_118_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24128__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24003_ _23363_/CLK _24003_/D VGND VGND VPWR VPWR _14797_/B sky130_fd_sc_hd__dfxtp_4
X_21215_ _21214_/X VGND VGND VPWR VPWR _21271_/A sky130_fd_sc_hd__buf_2
XANTENNA__22976__A2 _17893_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_32_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_65_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22195_ _22139_/X _22193_/X _14766_/B _22190_/X VGND VGND VPWR VPWR _22195_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21146_ _20748_/X _21140_/X _23978_/Q _21144_/X VGND VGND VPWR VPWR _23978_/D sky130_fd_sc_hd__o22a_4
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13508__A _15876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21077_ _20442_/X _21075_/X _16175_/B _21072_/X VGND VGND VPWR VPWR _21077_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12412__A _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20028_ _20027_/X VGND VGND VPWR VPWR _20028_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12850_ _12850_/A VGND VGND VPWR VPWR _12851_/A sky130_fd_sc_hd__buf_2
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11801_ _11800_/X VGND VGND VPWR VPWR _16231_/A sky130_fd_sc_hd__buf_2
X_12781_ _12799_/A _24020_/Q VGND VGND VPWR VPWR _12781_/X sky130_fd_sc_hd__or2_4
XFILLER_15_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21979_ _21799_/X _21974_/X _16381_/B _21978_/X VGND VGND VPWR VPWR _23514_/D sky130_fd_sc_hd__o22a_4
XFILLER_27_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17368__B1 _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14519_/X _14520_/B VGND VGND VPWR VPWR _14520_/X sky130_fd_sc_hd__or2_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13243__A _13243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11774_/A _11732_/B VGND VGND VPWR VPWR _11732_/X sky130_fd_sc_hd__or2_4
X_23718_ _23270_/CLK _21624_/X VGND VGND VPWR VPWR _14272_/B sky130_fd_sc_hd__dfxtp_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _12494_/A _14451_/B _14450_/X VGND VGND VPWR VPWR _14452_/C sky130_fd_sc_hd__and3_4
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21460__A _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _13886_/A VGND VGND VPWR VPWR _11664_/A sky130_fd_sc_hd__buf_2
X_23649_ _23073_/CLK _23649_/D VGND VGND VPWR VPWR _23649_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13354_/X _13326_/B VGND VGND VPWR VPWR _13402_/X sky130_fd_sc_hd__or2_4
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ _17322_/B VGND VGND VPWR VPWR _17845_/A sky130_fd_sc_hd__buf_2
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ _13847_/A VGND VGND VPWR VPWR _15632_/A sky130_fd_sc_hd__buf_2
XFILLER_70_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _11594_/A VGND VGND VPWR VPWR _11595_/A sky130_fd_sc_hd__buf_2
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16121_ _16121_/A _16121_/B _16121_/C VGND VGND VPWR VPWR _16122_/B sky130_fd_sc_hd__or3_4
Xclkbuf_7_114_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR _23699_/CLK sky130_fd_sc_hd__clkbuf_1
X_13333_ _13428_/A _24080_/Q VGND VGND VPWR VPWR _13333_/X sky130_fd_sc_hd__or2_4
XFILLER_70_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11698__A _12383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14074__A _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16052_ _11745_/X _16052_/B _16052_/C VGND VGND VPWR VPWR _16060_/B sky130_fd_sc_hd__or3_4
X_13264_ _13257_/A _13190_/B VGND VGND VPWR VPWR _13264_/X sky130_fd_sc_hd__or2_4
XFILLER_109_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15003_ _14588_/X _23647_/Q VGND VGND VPWR VPWR _15005_/B sky130_fd_sc_hd__or2_4
XFILLER_100_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12215_ _12250_/A VGND VGND VPWR VPWR _12216_/A sky130_fd_sc_hd__buf_2
X_13195_ _12435_/A _13193_/X _13194_/X VGND VGND VPWR VPWR _13195_/X sky130_fd_sc_hd__and3_4
XANTENNA__19832__A2 _19828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19811_ _19800_/B _19810_/X _19793_/B VGND VGND VPWR VPWR _19812_/C sky130_fd_sc_hd__o21a_4
X_12146_ _11827_/A _12146_/B VGND VGND VPWR VPWR _12146_/X sky130_fd_sc_hd__or2_4
XANTENNA__15617__B _23595_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19742_ _19742_/A _19742_/B VGND VGND VPWR VPWR _19742_/X sky130_fd_sc_hd__or2_4
X_12077_ _11996_/A _12139_/B VGND VGND VPWR VPWR _12077_/X sky130_fd_sc_hd__or2_4
X_16954_ _24122_/Q VGND VGND VPWR VPWR _16974_/A sky130_fd_sc_hd__inv_2
XANTENNA__12322__A _15706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15905_ _13572_/A _15905_/B _15905_/C VGND VGND VPWR VPWR _15906_/C sky130_fd_sc_hd__and3_4
X_19673_ _19607_/X _19669_/Y _19580_/X _19672_/X VGND VGND VPWR VPWR _19673_/X sky130_fd_sc_hd__a211o_4
X_16885_ _16525_/X _16816_/X _16815_/A VGND VGND VPWR VPWR _16885_/X sky130_fd_sc_hd__o21a_4
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16729__A _12068_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18624_ _17779_/X _18616_/X _18617_/Y _18619_/X _18623_/Y VGND VGND VPWR VPWR _18624_/X
+ sky130_fd_sc_hd__a32o_4
X_15836_ _12886_/A _15836_/B VGND VGND VPWR VPWR _15836_/X sky130_fd_sc_hd__or2_4
XFILLER_20_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19348__B2 _20833_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18555_ _16998_/A _16969_/B _16970_/B VGND VGND VPWR VPWR _22927_/B sky130_fd_sc_hd__a21bo_4
XFILLER_111_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12979_ _12955_/A _12979_/B _12979_/C VGND VGND VPWR VPWR _12987_/B sky130_fd_sc_hd__or3_4
X_15767_ _15743_/A _15765_/X _15766_/X VGND VGND VPWR VPWR _15767_/X sky130_fd_sc_hd__and3_4
XANTENNA__14249__A _14345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21155__B2 _21151_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22352__B1 _12607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17506_ _17506_/A _17506_/B VGND VGND VPWR VPWR _17506_/X sky130_fd_sc_hd__or2_4
XANTENNA__13153__A _12728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14718_ _14040_/X _14702_/X _14717_/X VGND VGND VPWR VPWR _14718_/X sky130_fd_sc_hd__or3_4
X_18486_ _17634_/X VGND VGND VPWR VPWR _18486_/X sky130_fd_sc_hd__buf_2
X_15698_ _12737_/A _15696_/X _15697_/X VGND VGND VPWR VPWR _15698_/X sky130_fd_sc_hd__and3_4
XFILLER_107_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17437_ _17436_/X VGND VGND VPWR VPWR _17437_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14649_ _15203_/A VGND VGND VPWR VPWR _14673_/A sky130_fd_sc_hd__buf_2
XANTENNA__15385__A2 _15251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17368_ _15713_/Y _17340_/X _17021_/A _17367_/X VGND VGND VPWR VPWR _17371_/B sky130_fd_sc_hd__o22a_4
XANTENNA__22655__B2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19107_ _19106_/X VGND VGND VPWR VPWR _24319_/D sky130_fd_sc_hd__inv_2
X_16319_ _16303_/X _16317_/X _16318_/X VGND VGND VPWR VPWR _16320_/C sky130_fd_sc_hd__and3_4
X_17299_ _17552_/A VGND VGND VPWR VPWR _17299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24292__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19038_ _24364_/Q VGND VGND VPWR VPWR _19038_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16885__A2 _16816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17295__A _14564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15808__A _12879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_19_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14712__A _14673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21000_ _24191_/Q _20370_/A _20999_/Y VGND VGND VPWR VPWR _21001_/A sky130_fd_sc_hd__o21a_4
XFILLER_114_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21091__B1 _15855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21630__A2 _21626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12232__A _12202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22951_ _18475_/X _22950_/X VGND VGND VPWR VPWR _22952_/C sky130_fd_sc_hd__or2_4
XFILLER_112_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16639__A _16621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21394__B2 _21359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21902_ _21840_/X _21901_/X _23561_/Q _21898_/X VGND VGND VPWR VPWR _23561_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22882_ _22719_/X _19925_/X _22932_/A _19894_/X VGND VGND VPWR VPWR _22882_/X sky130_fd_sc_hd__or4_4
XFILLER_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19339__B2 _24236_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21833_ _21263_/A VGND VGND VPWR VPWR _21833_/X sky130_fd_sc_hd__buf_2
XANTENNA__15262__B _15262_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21146__B2 _21144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22343__B1 _16759_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24061__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21764_ _21546_/X _21762_/X _15902_/B _21759_/X VGND VGND VPWR VPWR _21764_/X sky130_fd_sc_hd__o22a_4
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22894__A1 _22886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21697__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23503_ _24047_/CLK _21994_/X VGND VGND VPWR VPWR _23503_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23629__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20715_ _20715_/A _20715_/B VGND VGND VPWR VPWR _20715_/Y sky130_fd_sc_hd__nor2_4
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13998__A _13998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21695_ _21687_/X VGND VGND VPWR VPWR _21695_/X sky130_fd_sc_hd__buf_2
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23434_ _23978_/CLK _23434_/D VGND VGND VPWR VPWR _14027_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20646_ _20753_/B VGND VGND VPWR VPWR _20699_/B sky130_fd_sc_hd__buf_2
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22646__B2 _22640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23365_ _23365_/CLK _23365_/D VGND VGND VPWR VPWR _14472_/B sky130_fd_sc_hd__dfxtp_4
X_20577_ _20229_/A _20576_/X _20284_/X VGND VGND VPWR VPWR _20577_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__12407__A _13102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23779__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22316_ _15669_/B VGND VGND VPWR VPWR _23310_/D sky130_fd_sc_hd__buf_2
X_23296_ _24180_/CLK _22330_/X VGND VGND VPWR VPWR _14875_/B sky130_fd_sc_hd__dfxtp_4
X_22247_ _22143_/X _22243_/X _15228_/B _22212_/A VGND VGND VPWR VPWR _23361_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15718__A _15725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14622__A _13600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12000_ _11943_/A _11810_/B VGND VGND VPWR VPWR _12000_/X sky130_fd_sc_hd__or2_4
XFILLER_69_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21621__A2 _21619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22178_ _22110_/X _22172_/X _13554_/B _22176_/X VGND VGND VPWR VPWR _22178_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14639__A1 _12267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14341__B _14268_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21129_ _20464_/X _21126_/X _12248_/B _21123_/X VGND VGND VPWR VPWR _23990_/D sky130_fd_sc_hd__o22a_4
XFILLER_8_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19578__A1 _19722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13951_ _13951_/A _23562_/Q VGND VGND VPWR VPWR _13951_/X sky130_fd_sc_hd__or2_4
XANTENNA__17652__B _17652_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20963__A1_N _19437_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21385__A1 _21273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16549__A _12025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21385__B2 _21380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11981__A _11980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12902_ _12520_/X _23827_/Q VGND VGND VPWR VPWR _12903_/C sky130_fd_sc_hd__or2_4
XFILLER_86_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_39_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR _24008_/CLK sky130_fd_sc_hd__clkbuf_1
X_13882_ _13910_/A _23527_/Q VGND VGND VPWR VPWR _13883_/C sky130_fd_sc_hd__or2_4
X_16670_ _16670_/A _24092_/Q VGND VGND VPWR VPWR _16671_/C sky130_fd_sc_hd__or2_4
XFILLER_46_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12796__B _12711_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12833_ _12803_/A _24084_/Q VGND VGND VPWR VPWR _12833_/X sky130_fd_sc_hd__or2_4
X_15621_ _15586_/A _23115_/Q VGND VGND VPWR VPWR _15621_/X sky130_fd_sc_hd__or2_4
XFILLER_62_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14069__A _14046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18340_ _18198_/A VGND VGND VPWR VPWR _18340_/X sky130_fd_sc_hd__buf_2
XFILLER_76_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12764_ _12412_/A VGND VGND VPWR VPWR _13097_/A sky130_fd_sc_hd__buf_2
X_15552_ _15552_/A _23883_/Q VGND VGND VPWR VPWR _15554_/B sky130_fd_sc_hd__or2_4
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22286__A _22286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21190__A _21183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _11715_/A VGND VGND VPWR VPWR _16025_/A sky130_fd_sc_hd__buf_2
X_14503_ _14556_/A _14501_/X _14503_/C VGND VGND VPWR VPWR _14503_/X sky130_fd_sc_hd__and3_4
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _12626_/A _15479_/X _15483_/C VGND VGND VPWR VPWR _15484_/C sky130_fd_sc_hd__or3_4
X_18271_ _17796_/X _18270_/X _17836_/X _17936_/X VGND VGND VPWR VPWR _18271_/X sky130_fd_sc_hd__o22a_4
X_12695_ _12695_/A _12695_/B _12694_/X VGND VGND VPWR VPWR _12696_/C sky130_fd_sc_hd__and3_4
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _18728_/A _17173_/A _17221_/Y _17157_/A VGND VGND VPWR VPWR _17222_/X sky130_fd_sc_hd__o22a_4
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ _11646_/A VGND VGND VPWR VPWR _11647_/A sky130_fd_sc_hd__buf_2
X_14434_ _15578_/A VGND VGND VPWR VPWR _14464_/A sky130_fd_sc_hd__buf_2
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22637__B2 _22633_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ _15643_/A _14351_/X _14364_/X VGND VGND VPWR VPWR _14365_/X sky130_fd_sc_hd__and3_4
X_17153_ _14429_/B _17131_/X _16235_/X _17133_/X VGND VGND VPWR VPWR _17153_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11577_ _17069_/A VGND VGND VPWR VPWR _17083_/A sky130_fd_sc_hd__buf_2
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12317__A _12705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13316_ _13491_/A _13290_/X _13298_/X _13307_/X _13315_/X VGND VGND VPWR VPWR _13316_/X
+ sky130_fd_sc_hd__a32o_4
X_16104_ _16109_/A _16104_/B _16103_/X VGND VGND VPWR VPWR _16105_/C sky130_fd_sc_hd__and3_4
X_17084_ _17084_/A _17083_/X _17900_/A VGND VGND VPWR VPWR _17084_/X sky130_fd_sc_hd__or3_4
X_14296_ _11955_/A _14296_/B VGND VGND VPWR VPWR _14297_/C sky130_fd_sc_hd__or2_4
XANTENNA__21860__A2 _21853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20534__A _20534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13247_ _13231_/A _13247_/B _13246_/X VGND VGND VPWR VPWR _13251_/B sky130_fd_sc_hd__and3_4
X_16035_ _16063_/A _16035_/B _16034_/X VGND VGND VPWR VPWR _16035_/X sky130_fd_sc_hd__and3_4
XFILLER_115_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21073__B1 _16390_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13178_ _12728_/A _13178_/B VGND VGND VPWR VPWR _13178_/X sky130_fd_sc_hd__or2_4
XFILLER_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18939__A _19027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12129_ _12153_/A _23773_/Q VGND VGND VPWR VPWR _12129_/X sky130_fd_sc_hd__or2_4
XANTENNA__13148__A _15685_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17986_ _17968_/X _17985_/X VGND VGND VPWR VPWR _17986_/Y sky130_fd_sc_hd__nor2_4
XFILLER_46_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19725_ _19826_/B VGND VGND VPWR VPWR _19726_/C sky130_fd_sc_hd__inv_2
XFILLER_111_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16937_ _16991_/A VGND VGND VPWR VPWR _16937_/X sky130_fd_sc_hd__buf_2
XFILLER_65_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12987__A _13083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19656_ _19659_/A _19573_/Y VGND VGND VPWR VPWR _19656_/X sky130_fd_sc_hd__and2_4
X_16868_ _14430_/X _16867_/X _14430_/X _16867_/X VGND VGND VPWR VPWR _16868_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18607_ _16965_/C VGND VGND VPWR VPWR _18607_/X sky130_fd_sc_hd__buf_2
X_15819_ _15823_/A _15819_/B _15818_/X VGND VGND VPWR VPWR _15820_/C sky130_fd_sc_hd__and3_4
X_19587_ HRDATA[27] VGND VGND VPWR VPWR _20358_/B sky130_fd_sc_hd__buf_2
X_16799_ _16799_/A _23707_/Q VGND VGND VPWR VPWR _16799_/X sky130_fd_sc_hd__or2_4
XANTENNA__21128__B2 _21123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18538_ _18538_/A VGND VGND VPWR VPWR _18538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21679__A2 _21676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18469_ _18469_/A VGND VGND VPWR VPWR _18469_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16194__A _16194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20500_ _20500_/A VGND VGND VPWR VPWR _20500_/X sky130_fd_sc_hd__buf_2
XFILLER_33_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13611__A _13611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21480_ _21263_/X _21477_/X _23788_/Q _21474_/X VGND VGND VPWR VPWR _21480_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22924__A _22924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24402__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20431_ _20622_/A _20430_/Y _24279_/Q _20301_/X VGND VGND VPWR VPWR _20431_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12227__A _13054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23150_ _23692_/CLK _23150_/D VGND VGND VPWR VPWR _15732_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20362_ _20255_/X _20361_/X _18954_/A _18872_/B VGND VGND VPWR VPWR _20362_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21851__A2 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17737__B _17127_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20444__A _20444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22101_ _22101_/A VGND VGND VPWR VPWR _22101_/X sky130_fd_sc_hd__buf_2
X_23081_ _23561_/CLK _22701_/X VGND VGND VPWR VPWR _23081_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15538__A _15571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20293_ _20518_/A VGND VGND VPWR VPWR _20293_/X sky130_fd_sc_hd__buf_2
X_22032_ _21804_/X _22031_/X _23480_/Q _22028_/X VGND VGND VPWR VPWR _22032_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21603__A2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23983_ _23983_/CLK _23983_/D VGND VGND VPWR VPWR _13531_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12897__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16369__A _16447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21367__B2 _21366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15273__A _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22934_ _22952_/A _22932_/Y _22934_/C VGND VGND VPWR VPWR _22934_/X sky130_fd_sc_hd__and3_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22865_ _17542_/Y _22863_/X _22853_/X _22864_/X VGND VGND VPWR VPWR _22866_/B sky130_fd_sc_hd__o22a_4
XFILLER_77_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22818__B _14493_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21816_ _21246_/A VGND VGND VPWR VPWR _21816_/X sky130_fd_sc_hd__buf_2
XFILLER_19_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22796_ _22795_/X VGND VGND VPWR VPWR _22796_/X sky130_fd_sc_hd__buf_2
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21747_ _21517_/X _21741_/X _16368_/B _21745_/X VGND VGND VPWR VPWR _23641_/D sky130_fd_sc_hd__o22a_4
XFILLER_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12280__A1 _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14617__A _14617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11500_ _18652_/A VGND VGND VPWR VPWR _22888_/A sky130_fd_sc_hd__inv_2
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12480_ _12528_/A _12464_/X _12480_/C VGND VGND VPWR VPWR _12480_/X sky130_fd_sc_hd__or3_4
X_24466_ _24066_/CLK _18290_/X HRESETn VGND VGND VPWR VPWR _24466_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21678_ _21570_/X _21676_/X _14779_/B _21673_/X VGND VGND VPWR VPWR _21678_/X sky130_fd_sc_hd__o22a_4
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24143__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23417_ _23354_/CLK _23417_/D VGND VGND VPWR VPWR _16283_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20629_ _20493_/X _20628_/X _24302_/Q _20500_/X VGND VGND VPWR VPWR _20630_/B sky130_fd_sc_hd__o22a_4
X_24397_ _24334_/CLK _18845_/X HRESETn VGND VGND VPWR VPWR _24397_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14150_ _15041_/A VGND VGND VPWR VPWR _14151_/A sky130_fd_sc_hd__buf_2
XANTENNA__18750__C _18327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23348_ _23987_/CLK _22271_/X VGND VGND VPWR VPWR _12767_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21842__A2 _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13101_ _13101_/A _13101_/B _13101_/C VGND VGND VPWR VPWR _13102_/C sky130_fd_sc_hd__or3_4
XANTENNA__11976__A _11976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14081_ _12196_/A _14081_/B _14080_/X VGND VGND VPWR VPWR _14086_/B sky130_fd_sc_hd__and3_4
XFILLER_10_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15448__A _15448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23044__A1 _22886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23279_ _24047_/CLK _22360_/X VGND VGND VPWR VPWR _23279_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14352__A _14367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20073__B _12098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13032_ _13032_/A _24050_/Q VGND VGND VPWR VPWR _13033_/C sky130_fd_sc_hd__or2_4
XFILLER_117_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18759__A _18759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17840_ _17825_/X _17838_/X _17806_/X _17839_/X VGND VGND VPWR VPWR _17840_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__18471__A1 _18424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17771_ _17640_/X _17770_/X _17640_/X _17770_/X VGND VGND VPWR VPWR _17771_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14983_ _14658_/A _14983_/B _14983_/C VGND VGND VPWR VPWR _14984_/C sky130_fd_sc_hd__or3_4
XFILLER_43_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21358__A1 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21358__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22555__B1 _14275_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19510_ _19729_/B VGND VGND VPWR VPWR _19511_/B sky130_fd_sc_hd__inv_2
X_16722_ _16718_/A _16720_/X _16722_/C VGND VGND VPWR VPWR _16726_/B sky130_fd_sc_hd__and3_4
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15183__A _14172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13934_ _15036_/A _14011_/B VGND VGND VPWR VPWR _13934_/X sky130_fd_sc_hd__or2_4
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18223__B2 _18222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19441_ _19441_/A VGND VGND VPWR VPWR _19442_/B sky130_fd_sc_hd__buf_2
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16653_ _16622_/A _16653_/B _16652_/X VGND VGND VPWR VPWR _16661_/B sky130_fd_sc_hd__or3_4
X_13865_ _13893_/A _13858_/X _13865_/C VGND VGND VPWR VPWR _13865_/X sky130_fd_sc_hd__or3_4
XFILLER_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18494__A _17422_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15604_ _15604_/A _15600_/X _15604_/C VGND VGND VPWR VPWR _15612_/B sky130_fd_sc_hd__or3_4
XANTENNA__15911__A _15907_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12816_ _12816_/A _23828_/Q VGND VGND VPWR VPWR _12817_/C sky130_fd_sc_hd__or2_4
X_19372_ _19370_/X _18020_/Y _19370_/X _24217_/Q VGND VGND VPWR VPWR _24217_/D sky130_fd_sc_hd__a2bb2o_4
X_16584_ _16569_/A _16582_/X _16584_/C VGND VGND VPWR VPWR _16584_/X sky130_fd_sc_hd__and3_4
XFILLER_90_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13796_ _13796_/A _13796_/B _13796_/C VGND VGND VPWR VPWR _13796_/X sky130_fd_sc_hd__and3_4
XFILLER_62_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18323_ _17864_/A _18070_/X _17845_/X _18072_/X VGND VGND VPWR VPWR _18323_/X sky130_fd_sc_hd__o22a_4
XFILLER_91_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15535_ _15558_/A _15531_/X _15534_/X VGND VGND VPWR VPWR _15535_/X sky130_fd_sc_hd__or3_4
XFILLER_17_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15630__B _23787_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12747_ _12747_/A _12745_/X _12746_/X VGND VGND VPWR VPWR _12747_/X sky130_fd_sc_hd__and3_4
XFILLER_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21530__B2 _21527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20248__B _19926_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19333__A2_N _18337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13431__A _13463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18254_ _18254_/A _18254_/B VGND VGND VPWR VPWR _18254_/X sky130_fd_sc_hd__or2_4
XFILLER_15_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12678_ _12677_/X VGND VGND VPWR VPWR _12678_/Y sky130_fd_sc_hd__inv_2
X_15466_ _12585_/A _15403_/B VGND VGND VPWR VPWR _15466_/X sky130_fd_sc_hd__or2_4
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17205_ _17195_/Y _17131_/X _15909_/B _17133_/X VGND VGND VPWR VPWR _17205_/X sky130_fd_sc_hd__o22a_4
XFILLER_106_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11629_ _11628_/X VGND VGND VPWR VPWR _11629_/X sky130_fd_sc_hd__buf_2
X_14417_ _15632_/A _14417_/B VGND VGND VPWR VPWR _14417_/X sky130_fd_sc_hd__or2_4
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18185_ _18185_/A VGND VGND VPWR VPWR _18185_/Y sky130_fd_sc_hd__inv_2
X_15397_ _15424_/A _15397_/B _15396_/X VGND VGND VPWR VPWR _15398_/C sky130_fd_sc_hd__and3_4
XANTENNA__12047__A _11921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19756__C _19689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17136_ _17163_/A VGND VGND VPWR VPWR _17815_/A sky130_fd_sc_hd__buf_2
XFILLER_102_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21294__B1 _23903_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14348_ _14218_/X VGND VGND VPWR VPWR _15615_/A sky130_fd_sc_hd__buf_2
XANTENNA__19348__A2_N _18576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15358__A _14010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14279_ _15553_/A _14279_/B VGND VGND VPWR VPWR _14279_/X sky130_fd_sc_hd__or2_4
X_17067_ _17054_/A _16909_/B _16910_/X VGND VGND VPWR VPWR _18750_/A sky130_fd_sc_hd__o21a_4
XANTENNA__14262__A _14261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21046__B1 _13745_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16018_ _11684_/X _16011_/X _16018_/C VGND VGND VPWR VPWR _16029_/B sky130_fd_sc_hd__or3_4
XFILLER_69_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21597__B2 _21595_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17969_ _17864_/A VGND VGND VPWR VPWR _17969_/X sky130_fd_sc_hd__buf_2
XANTENNA__16189__A _16227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22546__B1 _15462_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19708_ _19534_/X _19701_/X _19704_/Y _19707_/X VGND VGND VPWR VPWR _19708_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15093__A _15115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22010__A2 _22009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20980_ _24192_/Q _20873_/X _20979_/X VGND VGND VPWR VPWR _22460_/A sky130_fd_sc_hd__o21a_4
XANTENNA__12510__A _13641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19639_ _19639_/A _19643_/B VGND VGND VPWR VPWR _19640_/B sky130_fd_sc_hd__or2_4
XANTENNA__13325__B _13325_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_22_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR _24187_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_85_0_HCLK clkbuf_6_42_0_HCLK/X VGND VGND VPWR VPWR _24277_/CLK sky130_fd_sc_hd__clkbuf_1
X_22650_ _22621_/A VGND VGND VPWR VPWR _22650_/X sky130_fd_sc_hd__buf_2
XFILLER_53_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20439__A _20484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21601_ _21524_/X _21598_/X _12224_/B _21595_/X VGND VGND VPWR VPWR _21601_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15540__B _23531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22581_ _22406_/X _22579_/X _16186_/B _22576_/X VGND VGND VPWR VPWR _23159_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21521__B2 _21515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24320_ _24320_/CLK _24320_/D HRESETn VGND VGND VPWR VPWR _24320_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__13341__A _15697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21532_ _21532_/A VGND VGND VPWR VPWR _21532_/X sky130_fd_sc_hd__buf_2
XANTENNA__22654__A _22633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24251_ _24216_/CLK _19316_/X HRESETn VGND VGND VPWR VPWR _24251_/Q sky130_fd_sc_hd__dfrtp_4
X_21463_ _21470_/A VGND VGND VPWR VPWR _21463_/X sky130_fd_sc_hd__buf_2
XANTENNA__16652__A _16652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23202_ _23812_/CLK _23202_/D VGND VGND VPWR VPWR _15299_/B sky130_fd_sc_hd__dfxtp_4
X_20414_ _20414_/A VGND VGND VPWR VPWR _20414_/Y sky130_fd_sc_hd__inv_2
X_24182_ _24180_/CLK _19679_/X HRESETn VGND VGND VPWR VPWR _11592_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21394_ _21289_/X _21390_/X _15180_/B _21359_/A VGND VGND VPWR VPWR _23841_/D sky130_fd_sc_hd__o22a_4
XFILLER_68_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23133_ _24092_/CLK _23133_/D VGND VGND VPWR VPWR _12159_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__11796__A _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20345_ _20255_/X _20344_/X _24379_/Q _18872_/B VGND VGND VPWR VPWR _20345_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14172__A _14172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23064_ _22898_/A _23064_/B _23064_/C _23062_/Y VGND VGND VPWR VPWR HTRANS[1] sky130_fd_sc_hd__or4_4
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20276_ _20276_/A VGND VGND VPWR VPWR _21789_/A sky130_fd_sc_hd__buf_2
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22015_ _21863_/X _21988_/A _23487_/Q _21970_/X VGND VGND VPWR VPWR _23487_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17483__A _13591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19650__B1 _20400_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15715__B _15715_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13516__A _13511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22001__A2 _21995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11980_ _11980_/A VGND VGND VPWR VPWR _11980_/X sky130_fd_sc_hd__buf_2
X_23966_ _23774_/CLK _21167_/X VGND VGND VPWR VPWR _21161_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__20012__A1 _19994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22917_ _22899_/X _22917_/B _22917_/C VGND VGND VPWR VPWR _22917_/X sky130_fd_sc_hd__and3_4
X_23897_ _23770_/CLK _23897_/D VGND VGND VPWR VPWR _16272_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21760__B2 _21759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24395__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15731__A _12765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13650_ _13647_/A VGND VGND VPWR VPWR _15442_/A sky130_fd_sc_hd__buf_2
X_22848_ _17466_/Y _22824_/X _22777_/X _22847_/X VGND VGND VPWR VPWR _22849_/A sky130_fd_sc_hd__a211o_4
XFILLER_32_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12601_ _12646_/A VGND VGND VPWR VPWR _12963_/A sky130_fd_sc_hd__buf_2
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13581_ _13280_/X _13580_/Y VGND VGND VPWR VPWR _13581_/Y sky130_fd_sc_hd__nor2_4
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ _18720_/X _22778_/Y _16910_/X VGND VGND VPWR VPWR _22779_/X sky130_fd_sc_hd__o21a_4
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13251__A _13211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12532_ _15398_/A VGND VGND VPWR VPWR _12533_/A sky130_fd_sc_hd__buf_2
X_15320_ _15334_/A _15317_/X _15320_/C VGND VGND VPWR VPWR _15320_/X sky130_fd_sc_hd__and3_4
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18761__B _18866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12463_ _12865_/A _12463_/B VGND VGND VPWR VPWR _12463_/X sky130_fd_sc_hd__or2_4
X_15251_ _15251_/A VGND VGND VPWR VPWR _15251_/X sky130_fd_sc_hd__buf_2
XFILLER_71_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19469__B1 HRDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24449_ _24203_/CLK _24449_/D HRESETn VGND VGND VPWR VPWR _24449_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23347__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16562__A _11982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14202_ _14202_/A _14190_/X _14202_/C VGND VGND VPWR VPWR _14202_/X sky130_fd_sc_hd__and3_4
X_15182_ _15032_/A _15178_/X _15182_/C VGND VGND VPWR VPWR _15183_/B sky130_fd_sc_hd__or3_4
X_12394_ _12828_/A _12287_/B VGND VGND VPWR VPWR _12395_/C sky130_fd_sc_hd__or2_4
XANTENNA__21815__A2 _21805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14133_ _14315_/A _23593_/Q VGND VGND VPWR VPWR _14135_/B sky130_fd_sc_hd__or2_4
X_19990_ _19990_/A VGND VGND VPWR VPWR _19990_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14082__A _15146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14064_ _14035_/A _24074_/Q VGND VGND VPWR VPWR _14065_/C sky130_fd_sc_hd__or2_4
X_18941_ _18994_/A VGND VGND VPWR VPWR _18941_/X sky130_fd_sc_hd__buf_2
XFILLER_113_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21908__A _21901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21579__B2 _21515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13015_ _13015_/A _23314_/Q VGND VGND VPWR VPWR _13017_/B sky130_fd_sc_hd__or2_4
X_18872_ _18762_/A _18872_/B VGND VGND VPWR VPWR _18873_/A sky130_fd_sc_hd__or2_4
XANTENNA__15906__A _12672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14810__A _14810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17823_ _17975_/A VGND VGND VPWR VPWR _17823_/X sky130_fd_sc_hd__buf_2
XFILLER_79_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15625__B _23403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22528__B1 _16248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13426__A _13350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17754_ _17697_/A _17754_/B _17753_/X VGND VGND VPWR VPWR _18164_/A sky130_fd_sc_hd__and3_4
XFILLER_110_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14966_ _15074_/A _14899_/B VGND VGND VPWR VPWR _14966_/X sky130_fd_sc_hd__or2_4
XANTENNA__12330__A _12744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20003__A1 _19994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16705_ _11903_/A _23579_/Q VGND VGND VPWR VPWR _16706_/C sky130_fd_sc_hd__or2_4
X_13917_ _11799_/A _13901_/X _13917_/C VGND VGND VPWR VPWR _13918_/C sky130_fd_sc_hd__or3_4
X_17685_ _17685_/A VGND VGND VPWR VPWR _17685_/Y sky130_fd_sc_hd__inv_2
X_14897_ _13982_/A _14895_/X _14897_/C VGND VGND VPWR VPWR _14901_/B sky130_fd_sc_hd__and3_4
XFILLER_35_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16737__A _11943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21751__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19424_ _19424_/A VGND VGND VPWR VPWR _19545_/A sky130_fd_sc_hd__buf_2
XFILLER_39_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16636_ _16629_/X VGND VGND VPWR VPWR _16662_/A sky130_fd_sc_hd__buf_2
XFILLER_78_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13848_ _13878_/A _23335_/Q VGND VGND VPWR VPWR _13848_/X sky130_fd_sc_hd__or2_4
XFILLER_35_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19355_ _19370_/A VGND VGND VPWR VPWR _19355_/X sky130_fd_sc_hd__buf_2
X_16567_ _16567_/A _23612_/Q VGND VGND VPWR VPWR _16569_/B sky130_fd_sc_hd__or2_4
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13779_ _12861_/A _13777_/X _13778_/X VGND VGND VPWR VPWR _13783_/B sky130_fd_sc_hd__and3_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20306__A2 _20304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18306_ _18189_/X _18278_/X _18189_/X _18275_/X VGND VGND VPWR VPWR _18307_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13161__A _15695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15518_ _15453_/Y _15517_/X VGND VGND VPWR VPWR _15518_/X sky130_fd_sc_hd__and2_4
X_19286_ _24261_/Q _19209_/X _19285_/Y VGND VGND VPWR VPWR _24261_/D sky130_fd_sc_hd__o21a_4
X_16498_ _16473_/X _16435_/B VGND VGND VPWR VPWR _16499_/C sky130_fd_sc_hd__or2_4
XANTENNA__17183__A1 _14263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18237_ _18237_/A VGND VGND VPWR VPWR _18237_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15449_ _15449_/A _15449_/B _15448_/X VGND VGND VPWR VPWR _15449_/X sky130_fd_sc_hd__or3_4
XANTENNA__21267__B1 _23915_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18168_ _17755_/X _18167_/X _17755_/X _18167_/X VGND VGND VPWR VPWR _18168_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21806__A2 _21805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17119_ _17150_/A VGND VGND VPWR VPWR _17120_/A sky130_fd_sc_hd__inv_2
X_18099_ _18239_/A _17567_/X VGND VGND VPWR VPWR _18099_/X sky130_fd_sc_hd__or2_4
XANTENNA__12505__A _13029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20130_ _19313_/A _20129_/X VGND VGND VPWR VPWR _20130_/X sky130_fd_sc_hd__or2_4
XFILLER_67_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18399__A _17338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20722__A _20722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12224__B _12224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20061_ _20060_/X VGND VGND VPWR VPWR _20061_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15816__A _12859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22231__A2 _22229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19632__B1 _19866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14720__A _14719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20793__A2 _20784_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21990__B2 _21985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23820_ _23698_/CLK _23820_/D VGND VGND VPWR VPWR _23820_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_113_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12240__A _12240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23751_ _23847_/CLK _21561_/X VGND VGND VPWR VPWR _23751_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20963_ _19437_/Y _20850_/Y _20576_/B _20699_/B VGND VGND VPWR VPWR _20963_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20545__A2 _20544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22702_ _21843_/A _22700_/X _13756_/B _22697_/X VGND VGND VPWR VPWR _22702_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21742__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23682_ _23363_/CLK _21679_/X VGND VGND VPWR VPWR _15306_/B sky130_fd_sc_hd__dfxtp_4
X_20894_ _20872_/X _20893_/X _24068_/Q _20839_/X VGND VGND VPWR VPWR _24068_/D sky130_fd_sc_hd__o22a_4
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15421__A1 _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22633_ _22633_/A VGND VGND VPWR VPWR _22633_/X sky130_fd_sc_hd__buf_2
XANTENNA__22298__A2 _22293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22564_ _11779_/B VGND VGND VPWR VPWR _22564_/Y sky130_fd_sc_hd__inv_2
X_21515_ _21515_/A VGND VGND VPWR VPWR _21515_/X sky130_fd_sc_hd__buf_2
X_24303_ _23324_/CLK _24303_/D HRESETn VGND VGND VPWR VPWR _24303_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22495_ _22430_/X _22493_/X _15831_/B _22490_/X VGND VGND VPWR VPWR _23213_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16382__A _15948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24234_ _24202_/CLK _24234_/D HRESETn VGND VGND VPWR VPWR _20743_/A sky130_fd_sc_hd__dfrtp_4
X_21446_ _21293_/X _21419_/A _23807_/Q _21401_/X VGND VGND VPWR VPWR _23807_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18123__B1 _17634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24165_ _24165_/CLK _19860_/X HRESETn VGND VGND VPWR VPWR _24165_/Q sky130_fd_sc_hd__dfrtp_4
X_21377_ _21258_/X _21376_/X _15766_/B _21373_/X VGND VGND VPWR VPWR _21377_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12415__A _12386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23116_ _23304_/CLK _23116_/D VGND VGND VPWR VPWR _15493_/B sky130_fd_sc_hd__dfxtp_4
X_20328_ _20251_/X _20324_/X _24284_/Q _20327_/X VGND VGND VPWR VPWR _20328_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24096_ _24290_/CLK _22750_/X HRESETn VGND VGND VPWR VPWR _22727_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_116_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23047_ _17880_/X _23038_/B VGND VGND VPWR VPWR _23048_/C sky130_fd_sc_hd__or2_4
XANTENNA__18426__A1 _18424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15726__A _12777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20259_ _20258_/X VGND VGND VPWR VPWR _20449_/A sky130_fd_sc_hd__buf_2
XFILLER_1_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18102__A _18242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14820_ _13851_/A _14820_/B VGND VGND VPWR VPWR _14821_/C sky130_fd_sc_hd__or2_4
XFILLER_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12150__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21463__A _21470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14751_ _14778_/A _14751_/B _14751_/C VGND VGND VPWR VPWR _14752_/C sky130_fd_sc_hd__and3_4
X_11963_ _11962_/X VGND VGND VPWR VPWR _11997_/A sky130_fd_sc_hd__buf_2
X_23949_ _23698_/CLK _21192_/X VGND VGND VPWR VPWR _15815_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_56_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16557__A _12025_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13702_ _15486_/A _13702_/B VGND VGND VPWR VPWR _13702_/X sky130_fd_sc_hd__or2_4
X_17470_ _17466_/Y _17014_/X _17022_/A _17469_/Y VGND VGND VPWR VPWR _17527_/B sky130_fd_sc_hd__o22a_4
X_11894_ _11894_/A VGND VGND VPWR VPWR _15393_/A sky130_fd_sc_hd__buf_2
X_14682_ _14341_/A _14682_/B VGND VGND VPWR VPWR _14682_/X sky130_fd_sc_hd__or2_4
XFILLER_72_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16421_ _16002_/A _16421_/B VGND VGND VPWR VPWR _16421_/X sky130_fd_sc_hd__or2_4
X_13633_ _12203_/A VGND VGND VPWR VPWR _15436_/A sky130_fd_sc_hd__buf_2
XANTENNA__15180__B _15180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22289__A2 _22286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19140_ _19138_/X VGND VGND VPWR VPWR _19140_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24295__CLK _24299_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21497__B1 _23775_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16352_ _11727_/X _16350_/X _16352_/C VGND VGND VPWR VPWR _16353_/C sky130_fd_sc_hd__and3_4
X_13564_ _12753_/X _13560_/X _13563_/X VGND VGND VPWR VPWR _13572_/B sky130_fd_sc_hd__or3_4
XFILLER_73_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15303_ _14588_/X _15303_/B VGND VGND VPWR VPWR _15303_/X sky130_fd_sc_hd__or2_4
XFILLER_34_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12515_ _13048_/A _12515_/B _12514_/X VGND VGND VPWR VPWR _12516_/B sky130_fd_sc_hd__or3_4
X_19071_ _11511_/A _11511_/B _19066_/Y VGND VGND VPWR VPWR _19071_/Y sky130_fd_sc_hd__a21oi_4
X_13495_ _12958_/A VGND VGND VPWR VPWR _15876_/A sky130_fd_sc_hd__buf_2
X_16283_ _15934_/X _16283_/B VGND VGND VPWR VPWR _16284_/C sky130_fd_sc_hd__or2_4
XFILLER_9_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16292__A _15980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14805__A _14813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18022_ _18202_/A VGND VGND VPWR VPWR _18022_/X sky130_fd_sc_hd__buf_2
X_12446_ _11905_/Y VGND VGND VPWR VPWR _15045_/A sky130_fd_sc_hd__buf_2
X_15234_ _15234_/A _15177_/B VGND VGND VPWR VPWR _15234_/X sky130_fd_sc_hd__or2_4
X_12377_ _15882_/A _12370_/X _12376_/X VGND VGND VPWR VPWR _12390_/B sky130_fd_sc_hd__or3_4
X_15165_ _15142_/A _15228_/B VGND VGND VPWR VPWR _15165_/X sky130_fd_sc_hd__or2_4
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12325__A _12740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22461__A2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14116_ _14143_/A _23529_/Q VGND VGND VPWR VPWR _14117_/C sky130_fd_sc_hd__or2_4
X_15096_ _15104_/A _15096_/B _15096_/C VGND VGND VPWR VPWR _15100_/B sky130_fd_sc_hd__and3_4
X_19973_ _17948_/X _19961_/X _19971_/Y _19972_/X VGND VGND VPWR VPWR _19973_/X sky130_fd_sc_hd__o22a_4
XFILLER_113_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21638__A _21637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18924_ _11531_/X VGND VGND VPWR VPWR _18924_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14047_ _14847_/A _14043_/X _14047_/C VGND VGND VPWR VPWR _14055_/B sky130_fd_sc_hd__or3_4
XANTENNA__19108__A _19108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18855_ _18841_/A VGND VGND VPWR VPWR _18855_/X sky130_fd_sc_hd__buf_2
XANTENNA__19090__A1 _18965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17806_ _17817_/A VGND VGND VPWR VPWR _17806_/X sky130_fd_sc_hd__buf_2
XANTENNA__13156__A _15706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21972__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18786_ _13270_/X _18781_/X _20558_/A _18782_/X VGND VGND VPWR VPWR _18786_/X sky130_fd_sc_hd__o22a_4
X_15998_ _15948_/A _15998_/B _15998_/C VGND VGND VPWR VPWR _16004_/B sky130_fd_sc_hd__and3_4
XFILLER_67_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15651__A1 _15582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22469__A _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21373__A _21373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17737_ _17737_/A _17127_/Y VGND VGND VPWR VPWR _17738_/A sky130_fd_sc_hd__or2_4
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14949_ _15072_/A _14875_/B VGND VGND VPWR VPWR _14949_/X sky130_fd_sc_hd__or2_4
XFILLER_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_20_0_HCLK_A clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21724__B2 _21723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15371__A _14810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23512__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17668_ _24129_/Q _17442_/A _17667_/X VGND VGND VPWR VPWR _17668_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16186__B _16186_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19407_ _19403_/X _18645_/X _19406_/X _24196_/Q VGND VGND VPWR VPWR _24196_/D sky130_fd_sc_hd__a2bb2o_4
X_16619_ _16618_/X VGND VGND VPWR VPWR _16651_/A sky130_fd_sc_hd__buf_2
XFILLER_63_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17599_ _18567_/B _17598_/Y _17397_/X VGND VGND VPWR VPWR _17599_/Y sky130_fd_sc_hd__o21ai_4
X_19338_ _19336_/X _18432_/X _19336_/X _24237_/Q VGND VGND VPWR VPWR _24237_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19269_ _19219_/B VGND VGND VPWR VPWR _19269_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14715__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21300_ _21300_/A VGND VGND VPWR VPWR _21316_/A sky130_fd_sc_hd__inv_2
X_22280_ _22112_/X _22279_/X _15655_/B _22276_/X VGND VGND VPWR VPWR _23342_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22932__A _22932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21231_ _21229_/X _21223_/X _16404_/B _21230_/X VGND VGND VPWR VPWR _21231_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24018__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12235__A _12235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21162_ _21348_/A _21112_/B _21162_/C _20199_/B VGND VGND VPWR VPWR _21162_/X sky130_fd_sc_hd__or4_4
X_20113_ _11558_/B VGND VGND VPWR VPWR _20113_/Y sky130_fd_sc_hd__inv_2
X_21093_ _21079_/A VGND VGND VPWR VPWR _21093_/X sky130_fd_sc_hd__buf_2
XANTENNA__18408__B2 _18407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14450__A _13020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12889__B _23443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20044_ _19996_/A VGND VGND VPWR VPWR _20044_/X sky130_fd_sc_hd__buf_2
XFILLER_98_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21963__B2 _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24336__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23803_ _23867_/CLK _21459_/X VGND VGND VPWR VPWR _23803_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19908__B2 _20358_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21995_ _21988_/A VGND VGND VPWR VPWR _21995_/X sky130_fd_sc_hd__buf_2
XFILLER_27_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16377__A _16302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21715__B2 _21709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20946_ _24385_/Q _20405_/A _11541_/A _20449_/A VGND VGND VPWR VPWR _20946_/X sky130_fd_sc_hd__o22a_4
X_23734_ _23920_/CLK _21601_/X VGND VGND VPWR VPWR _12224_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21191__A2 _21190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16096__B _16096_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _20841_/X _20876_/X VGND VGND VPWR VPWR _20877_/X sky130_fd_sc_hd__and2_4
X_23665_ _23122_/CLK _23665_/D VGND VGND VPWR VPWR _13153_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_55_0_HCLK clkbuf_6_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21479__B1 _15836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22616_ _22616_/A VGND VGND VPWR VPWR _22621_/A sky130_fd_sc_hd__buf_2
XFILLER_39_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23596_ _23794_/CLK _21834_/X VGND VGND VPWR VPWR _23596_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22140__B2 _22132_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12129__B _23773_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22547_ _22533_/A VGND VGND VPWR VPWR _22547_/X sky130_fd_sc_hd__buf_2
XANTENNA__22620__A2_N _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18895__A1 _13274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22691__A2 _22686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12300_ _12706_/A _12295_/X _12299_/X VGND VGND VPWR VPWR _12300_/X sky130_fd_sc_hd__or3_4
XFILLER_33_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13280_ _13277_/X _13280_/B VGND VGND VPWR VPWR _13280_/X sky130_fd_sc_hd__or2_4
X_22478_ _22401_/X _22472_/X _16289_/B _22476_/X VGND VGND VPWR VPWR _23225_/D sky130_fd_sc_hd__o22a_4
XFILLER_10_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12231_ _12198_/X VGND VGND VPWR VPWR _12695_/A sky130_fd_sc_hd__buf_2
X_21429_ _21263_/X _21426_/X _23820_/Q _21423_/X VGND VGND VPWR VPWR _23820_/D sky130_fd_sc_hd__o22a_4
X_24217_ _24216_/CLK _24217_/D HRESETn VGND VGND VPWR VPWR _24217_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18647__A1 _17742_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22443__A2 _22440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12145__A _12169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12162_ _11774_/A _12162_/B VGND VGND VPWR VPWR _12162_/X sky130_fd_sc_hd__or2_4
X_24148_ _24223_/CLK _24148_/D HRESETn VGND VGND VPWR VPWR _24148_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17655__B _17652_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15456__A _15495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12093_ _12093_/A _12162_/B VGND VGND VPWR VPWR _12095_/B sky130_fd_sc_hd__or2_4
X_16970_ _16970_/A _16970_/B VGND VGND VPWR VPWR _16971_/B sky130_fd_sc_hd__or2_4
X_24079_ _23311_/CLK _20612_/X VGND VGND VPWR VPWR _13566_/B sky130_fd_sc_hd__dfxtp_4
X_15921_ _15915_/X _15919_/Y _15920_/Y VGND VGND VPWR VPWR _15921_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_42_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21954__A1 _21843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21954__B2 _21949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18640_ _18487_/X _18632_/Y _18633_/X _17998_/X _18639_/X VGND VGND VPWR VPWR _18640_/X
+ sky130_fd_sc_hd__a32o_4
X_15852_ _12384_/X _15852_/B VGND VGND VPWR VPWR _15852_/X sky130_fd_sc_hd__or2_4
XFILLER_76_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14803_ _13862_/A _14803_/B VGND VGND VPWR VPWR _14803_/X sky130_fd_sc_hd__or2_4
X_18571_ _18458_/X _18560_/X _18485_/X _18570_/X VGND VGND VPWR VPWR _18571_/X sky130_fd_sc_hd__o22a_4
X_15783_ _15783_/A _15782_/X VGND VGND VPWR VPWR _15914_/C sky130_fd_sc_hd__or2_4
X_12995_ _12924_/X _12992_/X _12994_/Y VGND VGND VPWR VPWR _12996_/B sky130_fd_sc_hd__a21o_4
XANTENNA__21706__A1 _21531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21706__B2 _21702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17522_ _17476_/X _17521_/X VGND VGND VPWR VPWR _17522_/Y sky130_fd_sc_hd__nor2_4
XFILLER_45_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15191__A _15203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14734_ _14734_/A _14734_/B _14734_/C VGND VGND VPWR VPWR _14734_/X sky130_fd_sc_hd__and3_4
XFILLER_91_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11946_ _11998_/A _11946_/B _11945_/X VGND VGND VPWR VPWR _11947_/C sky130_fd_sc_hd__and3_4
XFILLER_55_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17386__A1 _17383_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17386__B2 _17385_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17453_ _12841_/X _17525_/B VGND VGND VPWR VPWR _17454_/A sky130_fd_sc_hd__or2_4
XANTENNA__21921__A _21920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19598__A _19598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14665_ _14679_/A _24004_/Q VGND VGND VPWR VPWR _14665_/X sky130_fd_sc_hd__or2_4
XANTENNA__20390__B1 _20389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11877_ _14912_/A VGND VGND VPWR VPWR _15146_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16404_ _16394_/X _16404_/B VGND VGND VPWR VPWR _16404_/X sky130_fd_sc_hd__or2_4
X_13616_ _15424_/A _13614_/X _13616_/C VGND VGND VPWR VPWR _13616_/X sky130_fd_sc_hd__and3_4
XFILLER_32_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17384_ _17273_/A VGND VGND VPWR VPWR _17384_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14596_ _12449_/A _14596_/B _14596_/C VGND VGND VPWR VPWR _14597_/C sky130_fd_sc_hd__and3_4
X_19123_ _24302_/Q _19123_/B VGND VGND VPWR VPWR _19124_/B sky130_fd_sc_hd__and2_4
XFILLER_9_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16335_ _16365_/A _16260_/B VGND VGND VPWR VPWR _16336_/C sky130_fd_sc_hd__or2_4
X_13547_ _13546_/X _13547_/B VGND VGND VPWR VPWR _13547_/X sky130_fd_sc_hd__or2_4
XANTENNA__18886__A1 _16374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22682__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19054_ _11514_/B VGND VGND VPWR VPWR _19054_/Y sky130_fd_sc_hd__inv_2
X_16266_ _16090_/A _16266_/B VGND VGND VPWR VPWR _16266_/X sky130_fd_sc_hd__or2_4
XANTENNA__21890__B1 _23569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13478_ _13477_/X _13566_/B VGND VGND VPWR VPWR _13478_/X sky130_fd_sc_hd__or2_4
X_18005_ _17651_/A _18004_/X _17651_/A _18004_/X VGND VGND VPWR VPWR _18005_/X sky130_fd_sc_hd__a2bb2o_4
X_15217_ _11661_/A _15217_/B _15217_/C VGND VGND VPWR VPWR _15249_/B sky130_fd_sc_hd__or3_4
XFILLER_12_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12429_ _11657_/X _12429_/B _12429_/C VGND VGND VPWR VPWR _12429_/X sky130_fd_sc_hd__and3_4
X_16197_ _16162_/X _16195_/X _16196_/X VGND VGND VPWR VPWR _16197_/X sky130_fd_sc_hd__and3_4
XANTENNA__12055__A _11875_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16750__A _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21642__B1 _23709_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15148_ _14998_/A _15146_/X _15147_/X VGND VGND VPWR VPWR _15148_/X sky130_fd_sc_hd__and3_4
XFILLER_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15366__A _14000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11894__A _11894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15079_ _12583_/A _15079_/B VGND VGND VPWR VPWR _15079_/X sky130_fd_sc_hd__or2_4
X_19956_ _19956_/A VGND VGND VPWR VPWR _19956_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14270__A _12320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22198__B2 _22162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18907_ _17171_/X _18905_/X _24362_/Q _18906_/X VGND VGND VPWR VPWR _18907_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19887_ _22824_/B VGND VGND VPWR VPWR _19887_/X sky130_fd_sc_hd__buf_2
XANTENNA__18810__A1 _15119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18838_ _13274_/X _18834_/X _24402_/Q _18835_/X VGND VGND VPWR VPWR _18838_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18810__B2 _18782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16821__B1 _16897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18769_ _11837_/X _18765_/X _24446_/Q _18768_/X VGND VGND VPWR VPWR _18769_/X sky130_fd_sc_hd__o22a_4
X_20800_ _20800_/A _20754_/B VGND VGND VPWR VPWR _20800_/X sky130_fd_sc_hd__or2_4
XANTENNA__13614__A _13614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21780_ _21574_/X _21776_/X _23617_/Q _21737_/X VGND VGND VPWR VPWR _21780_/X sky130_fd_sc_hd__o22a_4
XFILLER_97_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14429__B _14429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22370__B2 _22365_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20731_ _20492_/A VGND VGND VPWR VPWR _20731_/X sky130_fd_sc_hd__buf_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23450_ _23383_/CLK _22085_/X VGND VGND VPWR VPWR _16408_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20662_ _20517_/X _20661_/X _19122_/A _20527_/X VGND VGND VPWR VPWR _20663_/B sky130_fd_sc_hd__o22a_4
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20447__A _20447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22401_ _20393_/A VGND VGND VPWR VPWR _22401_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23381_ _23635_/CLK _23381_/D VGND VGND VPWR VPWR _12651_/B sky130_fd_sc_hd__dfxtp_4
X_20593_ _20511_/X _20591_/X _24080_/Q _20592_/X VGND VGND VPWR VPWR _24080_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22673__A2 _22672_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14445__A _12460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22332_ _11760_/B VGND VGND VPWR VPWR _22332_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20684__A1 _20681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20684__B2 _20625_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22263_ _22083_/X _22258_/X _16383_/B _22262_/X VGND VGND VPWR VPWR _23354_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16660__A _16599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24002_ _24066_/CLK _24002_/D VGND VGND VPWR VPWR _15262_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_105_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21214_ _21112_/A _21112_/B _21162_/C _21634_/D VGND VGND VPWR VPWR _21214_/X sky130_fd_sc_hd__or4_4
XFILLER_117_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21278__A _21242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22194_ _22136_/X _22193_/X _14620_/B _22190_/X VGND VGND VPWR VPWR _23396_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17301__A1 _17298_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17301__B2 _17300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21145_ _20723_/X _21140_/X _23979_/Q _21144_/X VGND VGND VPWR VPWR _23979_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15276__A _14588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15312__B1 _11594_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22189__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22189__B2 _22183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21076_ _20419_/X _21075_/X _24024_/Q _21072_/X VGND VGND VPWR VPWR _21076_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18587__A _18499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21936__B2 _21935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20027_ _20018_/X _17681_/A _20024_/X _20026_/X VGND VGND VPWR VPWR _20027_/X sky130_fd_sc_hd__o22a_4
XFILLER_98_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18801__A1 _14425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11800_ _12392_/A VGND VGND VPWR VPWR _11800_/X sky130_fd_sc_hd__buf_2
XFILLER_92_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12780_ _15724_/A VGND VGND VPWR VPWR _12799_/A sky130_fd_sc_hd__buf_2
XANTENNA__17368__A1 _15713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _21970_/X VGND VGND VPWR VPWR _21978_/X sky130_fd_sc_hd__buf_2
XFILLER_42_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17368__B2 _17367_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21741__A _21755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11731_ _16071_/A VGND VGND VPWR VPWR _11774_/A sky130_fd_sc_hd__buf_2
X_23717_ _23973_/CLK _21625_/X VGND VGND VPWR VPWR _14502_/B sky130_fd_sc_hd__dfxtp_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _20732_/X _20928_/X _19111_/A _20739_/X VGND VGND VPWR VPWR _20930_/B sky130_fd_sc_hd__o22a_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _13020_/A _14450_/B VGND VGND VPWR VPWR _14450_/X sky130_fd_sc_hd__or2_4
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _14039_/A VGND VGND VPWR VPWR _13886_/A sky130_fd_sc_hd__buf_2
X_23648_ _24180_/CLK _23648_/D VGND VGND VPWR VPWR _14872_/B sky130_fd_sc_hd__dfxtp_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13352_/X _13325_/B VGND VGND VPWR VPWR _13403_/B sky130_fd_sc_hd__or2_4
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11979__A _15812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ _11592_/X VGND VGND VPWR VPWR _11594_/A sky130_fd_sc_hd__buf_2
X_14381_ _13710_/A VGND VGND VPWR VPWR _15626_/A sky130_fd_sc_hd__buf_2
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23579_ _24026_/CLK _23579_/D VGND VGND VPWR VPWR _23579_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16120_ _16147_/A _16118_/X _16120_/C VGND VGND VPWR VPWR _16121_/C sky130_fd_sc_hd__and3_4
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ _13300_/A _23472_/Q VGND VGND VPWR VPWR _13332_/X sky130_fd_sc_hd__or2_4
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22572__A _22586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14074__B _14073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16051_ _16063_/A _16051_/B _16051_/C VGND VGND VPWR VPWR _16052_/C sky130_fd_sc_hd__and3_4
X_13263_ _13256_/A _13188_/B VGND VGND VPWR VPWR _13263_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15002_ _14119_/X _15002_/B _15002_/C VGND VGND VPWR VPWR _15002_/X sky130_fd_sc_hd__or3_4
X_12214_ _15654_/A _12206_/X _12213_/X VGND VGND VPWR VPWR _12214_/X sky130_fd_sc_hd__and3_4
XFILLER_48_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21624__B1 _14272_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13194_ _12315_/A _13254_/B VGND VGND VPWR VPWR _13194_/X sky130_fd_sc_hd__or2_4
XANTENNA__20978__A2 _20444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12145_ _12169_/A _12145_/B _12145_/C VGND VGND VPWR VPWR _12145_/X sky130_fd_sc_hd__and3_4
X_19810_ _19625_/Y _19801_/X _19809_/Y VGND VGND VPWR VPWR _19810_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12603__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12076_ _11995_/A _12074_/X _12076_/C VGND VGND VPWR VPWR _12080_/B sky130_fd_sc_hd__and3_4
X_16953_ _24123_/Q VGND VGND VPWR VPWR _17699_/A sky130_fd_sc_hd__inv_2
X_19741_ _19818_/A VGND VGND VPWR VPWR _19742_/B sky130_fd_sc_hd__inv_2
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17056__B1 _20206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21927__B2 _21921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15904_ _13507_/X _15904_/B _15904_/C VGND VGND VPWR VPWR _15905_/C sky130_fd_sc_hd__or3_4
X_19672_ _19670_/X _19442_/B _19672_/C _19672_/D VGND VGND VPWR VPWR _19672_/X sky130_fd_sc_hd__and4_4
XFILLER_77_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16884_ _12845_/X _16883_/X _12845_/X _16883_/X VGND VGND VPWR VPWR _16887_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18623_ _18623_/A VGND VGND VPWR VPWR _18623_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15835_ _12879_/A _15835_/B VGND VGND VPWR VPWR _15835_/X sky130_fd_sc_hd__or2_4
XANTENNA__15633__B _15577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18554_ _18381_/A VGND VGND VPWR VPWR _18554_/X sky130_fd_sc_hd__buf_2
XFILLER_20_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15766_ _12795_/A _15766_/B VGND VGND VPWR VPWR _15766_/X sky130_fd_sc_hd__or2_4
XFILLER_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12978_ _12954_/A _12978_/B _12978_/C VGND VGND VPWR VPWR _12979_/C sky130_fd_sc_hd__and3_4
XFILLER_111_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21155__A2 _21154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24382__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17505_ _16624_/X _17364_/X _17365_/X VGND VGND VPWR VPWR _17506_/B sky130_fd_sc_hd__o21a_4
XFILLER_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22352__B2 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14717_ _15643_/A _14709_/X _14716_/X VGND VGND VPWR VPWR _14717_/X sky130_fd_sc_hd__and3_4
X_11929_ _11929_/A VGND VGND VPWR VPWR _13813_/A sky130_fd_sc_hd__buf_2
X_18485_ _18202_/A VGND VGND VPWR VPWR _18485_/X sky130_fd_sc_hd__buf_2
X_15697_ _15697_/A _15697_/B VGND VGND VPWR VPWR _15697_/X sky130_fd_sc_hd__or2_4
X_17436_ _15782_/B _18387_/B _18405_/A _17435_/X VGND VGND VPWR VPWR _17436_/X sky130_fd_sc_hd__o22a_4
X_14648_ _13709_/A VGND VGND VPWR VPWR _15203_/A sky130_fd_sc_hd__buf_2
XANTENNA__18308__B1 _18048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22104__A1 _22103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22104__B2 _22096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _17506_/A _17367_/B VGND VGND VPWR VPWR _17367_/X sky130_fd_sc_hd__or2_4
XANTENNA__18859__A1 _14851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14579_ _15142_/A _14661_/B VGND VGND VPWR VPWR _14579_/X sky130_fd_sc_hd__or2_4
XANTENNA__22655__A2 _22650_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19106_ _18934_/A _19104_/Y _19102_/X _19105_/Y VGND VGND VPWR VPWR _19106_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20666__A1 _20640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16318_ _16323_/A _16253_/B VGND VGND VPWR VPWR _16318_/X sky130_fd_sc_hd__or2_4
XFILLER_119_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17298_ _14640_/X VGND VGND VPWR VPWR _17298_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17531__A1 _18153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19037_ _24332_/Q _11517_/B _19032_/Y VGND VGND VPWR VPWR _19037_/Y sky130_fd_sc_hd__a21oi_4
X_16249_ _16150_/A _16249_/B VGND VGND VPWR VPWR _16249_/X sky130_fd_sc_hd__or2_4
XANTENNA__22407__A2 _22404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16480__A _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21615__B1 _15459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15808__B _15863_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13609__A _15404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21091__B2 _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12513__A _13032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19939_ _20057_/A VGND VGND VPWR VPWR _19985_/A sky130_fd_sc_hd__buf_2
XANTENNA__23850__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15824__A _12518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22040__B1 _23474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22950_ _22980_/A VGND VGND VPWR VPWR _22950_/X sky130_fd_sc_hd__buf_2
XFILLER_68_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18200__A _18174_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21394__A2 _21390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22591__B2 _22590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21901_ _21901_/A VGND VGND VPWR VPWR _21901_/X sky130_fd_sc_hd__buf_2
XANTENNA__15543__B _23915_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22881_ _22862_/A _22881_/B VGND VGND VPWR VPWR HWDATA[31] sky130_fd_sc_hd__nor2_4
XFILLER_83_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13344__A _15785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_120_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR _24047_/CLK sky130_fd_sc_hd__clkbuf_1
X_21832_ _21831_/X _21829_/X _15879_/B _21824_/X VGND VGND VPWR VPWR _21832_/X sky130_fd_sc_hd__o22a_4
XFILLER_43_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22657__A _22621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21146__A2 _21140_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22343__B2 _22337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21763_ _21543_/X _21762_/X _15700_/B _21759_/X VGND VGND VPWR VPWR _23630_/D sky130_fd_sc_hd__o22a_4
XFILLER_73_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20714_ _20517_/X _20713_/X _19120_/A _20527_/X VGND VGND VPWR VPWR _20715_/B sky130_fd_sc_hd__o22a_4
X_23502_ _23564_/CLK _23502_/D VGND VGND VPWR VPWR _15715_/B sky130_fd_sc_hd__dfxtp_4
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21694_ _21512_/X _21691_/X _23675_/Q _21688_/X VGND VGND VPWR VPWR _23675_/D sky130_fd_sc_hd__o22a_4
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24104__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11799__A _11799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20645_ _20644_/X VGND VGND VPWR VPWR _20753_/B sky130_fd_sc_hd__inv_2
X_23433_ _23433_/CLK _23433_/D VGND VGND VPWR VPWR _23433_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22646__A2 _22643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18870__A _20407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23364_ _24066_/CLK _22244_/X VGND VGND VPWR VPWR _14698_/B sky130_fd_sc_hd__dfxtp_4
X_20576_ _20285_/X _20576_/B VGND VGND VPWR VPWR _20576_/X sky130_fd_sc_hd__and2_4
XANTENNA__22392__A _22416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14336__A1 _13594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22315_ _23311_/Q VGND VGND VPWR VPWR _22315_/X sky130_fd_sc_hd__buf_2
X_23295_ _23391_/CLK _22331_/X VGND VGND VPWR VPWR _15081_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16390__A _15999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14903__A _14906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22246_ _22141_/X _22243_/X _15292_/B _22240_/X VGND VGND VPWR VPWR _23362_/D sky130_fd_sc_hd__o22a_4
XFILLER_65_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13519__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22177_ _22107_/X _22172_/X _13329_/B _22176_/X VGND VGND VPWR VPWR _22177_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21128_ _20442_/X _21126_/X _23991_/Q _21123_/X VGND VGND VPWR VPWR _23991_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21736__A _21740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21909__A1 _21852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21909__B2 _21905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15734__A _15774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19578__A2 _19536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13950_ _11611_/A _23914_/Q VGND VGND VPWR VPWR _13952_/B sky130_fd_sc_hd__or2_4
X_21059_ _21007_/A _22017_/B _21212_/B VGND VGND VPWR VPWR _21060_/A sky130_fd_sc_hd__or3_4
XFILLER_4_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21385__A2 _21383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18786__B1 _20558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12901_ _12518_/X _12965_/B VGND VGND VPWR VPWR _12901_/X sky130_fd_sc_hd__or2_4
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13881_ _13909_/A _13794_/B VGND VGND VPWR VPWR _13883_/B sky130_fd_sc_hd__or2_4
X_15620_ _15604_/A _15616_/X _15620_/C VGND VGND VPWR VPWR _15620_/X sky130_fd_sc_hd__or3_4
XANTENNA__13254__A _13242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12832_ _12802_/A _12735_/B VGND VGND VPWR VPWR _12832_/X sky130_fd_sc_hd__or2_4
XFILLER_41_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22567__A _22600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15551_ _13597_/X _15528_/X _15535_/X _15542_/X _15550_/X VGND VGND VPWR VPWR _15551_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_43_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12763_ _12754_/X _12758_/X _12763_/C VGND VGND VPWR VPWR _12770_/B sky130_fd_sc_hd__and3_4
XFILLER_15_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14502_ _14533_/A _14502_/B VGND VGND VPWR VPWR _14503_/C sky130_fd_sc_hd__or2_4
XANTENNA__17210__B1 _14429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11713_/X VGND VGND VPWR VPWR _11715_/A sky130_fd_sc_hd__buf_2
X_18270_ _17969_/X _17979_/X _17975_/X _17983_/X VGND VGND VPWR VPWR _18270_/X sky130_fd_sc_hd__o22a_4
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _13097_/A _15482_/B _15481_/X VGND VGND VPWR VPWR _15483_/C sky130_fd_sc_hd__and3_4
XFILLER_43_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12240_/X _12784_/B VGND VGND VPWR VPWR _12694_/X sky130_fd_sc_hd__or2_4
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_25_0_HCLK clkbuf_5_24_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_25_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _15118_/X VGND VGND VPWR VPWR _17221_/Y sky130_fd_sc_hd__inv_2
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _15571_/A _14433_/B _14433_/C VGND VGND VPWR VPWR _14433_/X sky130_fd_sc_hd__and3_4
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11645_/A VGND VGND VPWR VPWR _11646_/A sky130_fd_sc_hd__buf_2
XANTENNA__22637__A2 _22636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17152_ _17130_/A VGND VGND VPWR VPWR _17152_/X sky130_fd_sc_hd__buf_2
XFILLER_89_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14364_ _14397_/A _14357_/X _14364_/C VGND VGND VPWR VPWR _14364_/X sky130_fd_sc_hd__or3_4
X_11576_ _20965_/A _11533_/X _24385_/Q _20070_/A VGND VGND VPWR VPWR _11576_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16103_ _16108_/A _16103_/B VGND VGND VPWR VPWR _16103_/X sky130_fd_sc_hd__or2_4
X_13315_ _12716_/X _13314_/X VGND VGND VPWR VPWR _13315_/X sky130_fd_sc_hd__and2_4
X_17083_ _17083_/A _17083_/B _17068_/A VGND VGND VPWR VPWR _17083_/X sky130_fd_sc_hd__and3_4
XANTENNA__15909__A _15844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14295_ _15543_/A _14373_/B VGND VGND VPWR VPWR _14295_/X sky130_fd_sc_hd__or2_4
XANTENNA__14813__A _14813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16034_ _16069_/A _15969_/B VGND VGND VPWR VPWR _16034_/X sky130_fd_sc_hd__or2_4
X_13246_ _13239_/A _13179_/B VGND VGND VPWR VPWR _13246_/X sky130_fd_sc_hd__or2_4
XANTENNA__13429__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21073__B2 _21072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13177_ _13317_/A _13173_/X _13176_/X VGND VGND VPWR VPWR _13177_/X sky130_fd_sc_hd__or3_4
XANTENNA__12333__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11561__A1 _24432_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20820__A1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12128_ _12152_/A _12128_/B VGND VGND VPWR VPWR _12128_/X sky130_fd_sc_hd__or2_4
XFILLER_96_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20820__B2 _20724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13148__B _24017_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17985_ _17862_/A _17980_/X _17836_/X _17984_/X VGND VGND VPWR VPWR _17985_/X sky130_fd_sc_hd__o22a_4
XFILLER_111_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12059_ _12091_/A _12132_/B VGND VGND VPWR VPWR _12060_/C sky130_fd_sc_hd__or2_4
X_16936_ _24139_/Q VGND VGND VPWR VPWR _16991_/A sky130_fd_sc_hd__inv_2
X_19724_ _19721_/Y _19723_/X _19667_/A VGND VGND VPWR VPWR _19724_/X sky130_fd_sc_hd__o21a_4
XFILLER_81_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15644__A _11799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22573__B2 _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16459__B _16390_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16867_ _15388_/X _14568_/Y _14566_/X VGND VGND VPWR VPWR _16867_/X sky130_fd_sc_hd__o21a_4
X_19655_ _19726_/B VGND VGND VPWR VPWR _19872_/C sky130_fd_sc_hd__buf_2
XFILLER_96_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13164__A _12709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15818_ _12895_/A _15818_/B VGND VGND VPWR VPWR _15818_/X sky130_fd_sc_hd__or2_4
X_18606_ _17745_/C _17745_/B _17745_/C _17745_/B VGND VGND VPWR VPWR _18606_/X sky130_fd_sc_hd__a2bb2o_4
X_19586_ _19549_/X _19555_/X _19584_/X _17273_/A _19585_/X VGND VGND VPWR VPWR _19586_/X
+ sky130_fd_sc_hd__a32o_4
X_16798_ _16757_/X _16796_/X _16797_/X VGND VGND VPWR VPWR _16798_/X sky130_fd_sc_hd__and3_4
XFILLER_46_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18537_ _17390_/B _18537_/B VGND VGND VPWR VPWR _18537_/Y sky130_fd_sc_hd__nand2_4
X_15749_ _13100_/A _15749_/B _15748_/X VGND VGND VPWR VPWR _15753_/B sky130_fd_sc_hd__and3_4
XFILLER_80_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20887__A1 _18641_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18468_ _18244_/A _18468_/B _18468_/C _18468_/D VGND VGND VPWR VPWR _18469_/A sky130_fd_sc_hd__or4_4
XFILLER_61_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17419_ _17418_/X VGND VGND VPWR VPWR _17419_/Y sky130_fd_sc_hd__inv_2
X_18399_ _17338_/X VGND VGND VPWR VPWR _18399_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22628__A2 _22622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20430_ _20430_/A VGND VGND VPWR VPWR _20430_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20361_ _24410_/Q _18814_/X _24442_/Q _20260_/X VGND VGND VPWR VPWR _20361_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15819__A _15823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22100_ _22100_/A VGND VGND VPWR VPWR _22100_/X sky130_fd_sc_hd__buf_2
XANTENNA__24442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23080_ _23368_/CLK _22702_/X VGND VGND VPWR VPWR _13756_/B sky130_fd_sc_hd__dfxtp_4
X_20292_ _20517_/A VGND VGND VPWR VPWR _20292_/X sky130_fd_sc_hd__buf_2
XFILLER_115_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22940__A _18528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_45_0_HCLK clkbuf_6_22_0_HCLK/X VGND VGND VPWR VPWR _23561_/CLK sky130_fd_sc_hd__clkbuf_1
X_22031_ _22031_/A VGND VGND VPWR VPWR _22031_/X sky130_fd_sc_hd__buf_2
XANTENNA__13339__A _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22261__B1 _16749_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12243__A _13048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21556__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15554__A _12307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22013__B1 _15126_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23982_ _24044_/CLK _23982_/D VGND VGND VPWR VPWR _15667_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21367__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22933_ _18548_/X _22945_/B VGND VGND VPWR VPWR _22934_/C sky130_fd_sc_hd__or2_4
XFILLER_60_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15273__B _15273_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20575__B1 _24081_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18865__A _12036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13074__A _13104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13057__A1 _12892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22864_ _22854_/X _22804_/X _17411_/Y _22855_/X VGND VGND VPWR VPWR _22864_/X sky130_fd_sc_hd__o22a_4
XFILLER_84_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22387__A _22386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21291__A _21291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21815_ _21814_/X _21805_/X _23604_/Q _21812_/X VGND VGND VPWR VPWR _21815_/X sky130_fd_sc_hd__o22a_4
X_22795_ _18720_/X _18752_/X VGND VGND VPWR VPWR _22795_/X sky130_fd_sc_hd__or2_4
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16385__A _11915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13802__A _13641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21746_ _21514_/X _21741_/X _16508_/B _21745_/X VGND VGND VPWR VPWR _23642_/D sky130_fd_sc_hd__o22a_4
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24465_ _24066_/CLK _18313_/X HRESETn VGND VGND VPWR VPWR _24465_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21677_ _21567_/X _21676_/X _14706_/B _21673_/X VGND VGND VPWR VPWR _21677_/X sky130_fd_sc_hd__o22a_4
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23416_ _23383_/CLK _23416_/D VGND VGND VPWR VPWR _23416_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20628_ _20494_/X _20627_/X _11519_/A _20453_/X VGND VGND VPWR VPWR _20628_/X sky130_fd_sc_hd__o22a_4
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24396_ _24334_/CLK _18846_/X HRESETn VGND VGND VPWR VPWR _24396_/Q sky130_fd_sc_hd__dfrtp_4
X_20559_ _20558_/Y _20521_/B VGND VGND VPWR VPWR _20559_/X sky130_fd_sc_hd__or2_4
X_23347_ _24082_/CLK _23347_/D VGND VGND VPWR VPWR _12928_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15729__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13100_ _13100_/A _13100_/B _13100_/C VGND VGND VPWR VPWR _13101_/C sky130_fd_sc_hd__and3_4
XANTENNA__24183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14080_ _14089_/A _23497_/Q VGND VGND VPWR VPWR _14080_/X sky130_fd_sc_hd__or2_4
X_23278_ _23922_/CLK _22362_/X VGND VGND VPWR VPWR _15725_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13031_ _13031_/A _23602_/Q VGND VGND VPWR VPWR _13031_/X sky130_fd_sc_hd__or2_4
XANTENNA__13249__A _13242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21055__B2 _21012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22229_ _22222_/A VGND VGND VPWR VPWR _22229_/X sky130_fd_sc_hd__buf_2
XFILLER_65_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17663__B _17664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_2_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11992__A _11982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17770_ _17641_/X _17768_/Y _17769_/X VGND VGND VPWR VPWR _17770_/X sky130_fd_sc_hd__o21a_4
X_14982_ _11642_/A _14980_/X _14982_/C VGND VGND VPWR VPWR _14983_/C sky130_fd_sc_hd__and3_4
XANTENNA__16279__B _16279_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16721_ _16698_/A _23835_/Q VGND VGND VPWR VPWR _16722_/C sky130_fd_sc_hd__or2_4
XANTENNA__22555__B2 _22554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13933_ _14782_/A _13928_/X _13933_/C VGND VGND VPWR VPWR _13933_/X sky130_fd_sc_hd__or3_4
XANTENNA__18223__A2 _19382_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18775__A _18782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19440_ _19545_/A _19436_/Y _19437_/Y _19439_/X VGND VGND VPWR VPWR _19441_/A sky130_fd_sc_hd__o22a_4
X_16652_ _16652_/A _16650_/X _16652_/C VGND VGND VPWR VPWR _16652_/X sky130_fd_sc_hd__and3_4
XFILLER_21_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13864_ _13880_/A _13859_/X _13864_/C VGND VGND VPWR VPWR _13865_/C sky130_fd_sc_hd__and3_4
XFILLER_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15603_ _15631_/A _15603_/B _15603_/C VGND VGND VPWR VPWR _15604_/C sky130_fd_sc_hd__and3_4
X_12815_ _12808_/A _23124_/Q VGND VGND VPWR VPWR _12815_/X sky130_fd_sc_hd__or2_4
X_19371_ _19367_/X _17953_/X _19370_/X _24218_/Q VGND VGND VPWR VPWR _24218_/D sky130_fd_sc_hd__a2bb2o_4
X_16583_ _16583_/A _23644_/Q VGND VGND VPWR VPWR _16584_/C sky130_fd_sc_hd__or2_4
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13795_ _13630_/A _23527_/Q VGND VGND VPWR VPWR _13796_/C sky130_fd_sc_hd__or2_4
XANTENNA__16295__A _11872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14808__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18322_ _18322_/A VGND VGND VPWR VPWR _18322_/Y sky130_fd_sc_hd__inv_2
X_15534_ _15534_/A _15532_/X _15533_/X VGND VGND VPWR VPWR _15534_/X sky130_fd_sc_hd__and3_4
XFILLER_63_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13712__A _11648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12746_ _12315_/A _23860_/Q VGND VGND VPWR VPWR _12746_/X sky130_fd_sc_hd__or2_4
XFILLER_16_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21530__A2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18253_ _18189_/X _18154_/X _18189_/X _18217_/B VGND VGND VPWR VPWR _18254_/B sky130_fd_sc_hd__a2bb2o_4
X_15465_ _15477_/A _15465_/B VGND VGND VPWR VPWR _15465_/X sky130_fd_sc_hd__or2_4
X_12677_ _12559_/X _12675_/Y VGND VGND VPWR VPWR _12677_/X sky130_fd_sc_hd__or2_4
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12328__A _12710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _17141_/X _17202_/X _17163_/A _17203_/X VGND VGND VPWR VPWR _17204_/X sky130_fd_sc_hd__o22a_4
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__B1 _11596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ _15626_/A _14414_/X _14415_/X VGND VGND VPWR VPWR _14416_/X sky130_fd_sc_hd__and3_4
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11628_ _20077_/D VGND VGND VPWR VPWR _11628_/X sky130_fd_sc_hd__buf_2
X_18184_ _17862_/A _18182_/X _18183_/X _18077_/X VGND VGND VPWR VPWR _18185_/A sky130_fd_sc_hd__o22a_4
XFILLER_54_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15396_ _13620_/A _15459_/B VGND VGND VPWR VPWR _15396_/X sky130_fd_sc_hd__or2_4
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ _17135_/A VGND VGND VPWR VPWR _17163_/A sky130_fd_sc_hd__buf_2
X_14347_ _15586_/A _14271_/B VGND VGND VPWR VPWR _14350_/B sky130_fd_sc_hd__or2_4
XANTENNA__21294__B2 _21230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22491__B1 _13336_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11559_ _11553_/X _11559_/B VGND VGND VPWR VPWR _20089_/D sky130_fd_sc_hd__or2_4
XANTENNA__18015__A _24190_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17066_ _17065_/X VGND VGND VPWR VPWR _18728_/B sky130_fd_sc_hd__buf_2
XFILLER_13_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14278_ _15552_/A _14278_/B VGND VGND VPWR VPWR _14278_/X sky130_fd_sc_hd__or2_4
XANTENNA__21046__A1 _20797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16017_ _16058_/A _16014_/X _16016_/X VGND VGND VPWR VPWR _16018_/C sky130_fd_sc_hd__and3_4
XANTENNA__13159__A _15697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13229_ _12373_/A VGND VGND VPWR VPWR _13242_/A sky130_fd_sc_hd__buf_2
XANTENNA__17854__A _18249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21046__B2 _21041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12063__A _11943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21376__A _21369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20280__A _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12998__A _12850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15374__A _12567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17968_ _18142_/A VGND VGND VPWR VPWR _17968_/X sky130_fd_sc_hd__buf_2
XFILLER_66_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22546__B2 _22540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16189__B _16189_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19707_ _19637_/Y _19705_/X _19445_/A _19706_/X VGND VGND VPWR VPWR _19707_/X sky130_fd_sc_hd__a211o_4
X_16919_ _16919_/A VGND VGND VPWR VPWR _16919_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17899_ _18203_/A _17282_/A VGND VGND VPWR VPWR _17899_/X sky130_fd_sc_hd__or2_4
XFILLER_66_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19638_ _19638_/A VGND VGND VPWR VPWR _19643_/B sky130_fd_sc_hd__inv_2
XFILLER_80_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15821__B _15821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19569_ _19424_/A _19568_/X HRDATA[4] _19439_/X VGND VGND VPWR VPWR _19570_/A sky130_fd_sc_hd__o22a_4
XFILLER_94_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14718__A _14040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21600_ _21522_/X _21598_/X _23735_/Q _21595_/X VGND VGND VPWR VPWR _23735_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13622__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22580_ _22403_/X _22579_/X _15967_/B _22576_/X VGND VGND VPWR VPWR _23160_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21521__A2 _21520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21531_ _21246_/A VGND VGND VPWR VPWR _21531_/X sky130_fd_sc_hd__buf_2
X_21462_ _21232_/X _21456_/X _16294_/B _21460_/X VGND VGND VPWR VPWR _23801_/D sky130_fd_sc_hd__o22a_4
X_24250_ _24250_/CLK _24250_/D HRESETn VGND VGND VPWR VPWR _24250_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20413_ _18087_/X _20238_/X _20319_/X _20412_/Y VGND VGND VPWR VPWR _20413_/X sky130_fd_sc_hd__a211o_4
X_23201_ _23145_/CLK _23201_/D VGND VGND VPWR VPWR _15243_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15549__A _12459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22482__B1 _12323_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21393_ _21287_/X _21390_/X _15307_/B _21387_/X VGND VGND VPWR VPWR _21393_/X sky130_fd_sc_hd__o22a_4
X_24181_ _23584_/CLK _24181_/D HRESETn VGND VGND VPWR VPWR _11974_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20174__B _20173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20344_ _24411_/Q _18814_/X _24443_/Q _20260_/X VGND VGND VPWR VPWR _20344_/X sky130_fd_sc_hd__o22a_4
X_23132_ _23324_/CLK _22624_/X VGND VGND VPWR VPWR _16654_/B sky130_fd_sc_hd__dfxtp_4
X_23063_ _20206_/A _23062_/Y VGND VGND VPWR VPWR HWRITE sky130_fd_sc_hd__and2_4
XANTENNA__13069__A _13104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22234__B1 _23371_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20275_ _20370_/A _20210_/X _20273_/X _24222_/Q _20484_/A VGND VGND VPWR VPWR _20276_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22014_ _21861_/X _22009_/X _14857_/B _21970_/X VGND VGND VPWR VPWR _23488_/D sky130_fd_sc_hd__o22a_4
XFILLER_118_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23299__CLK _23494_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19650__A1 _19497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20190__A _20190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12701__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22537__B2 _22533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23965_ _24026_/CLK _21170_/X VGND VGND VPWR VPWR _23965_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19402__B2 _24199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20012__A2 _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22916_ _18624_/X _22945_/B VGND VGND VPWR VPWR _22917_/C sky130_fd_sc_hd__or2_4
XFILLER_112_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23896_ _24088_/CLK _21313_/X VGND VGND VPWR VPWR _23896_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21760__A2 _21755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22847_ _14493_/Y _22778_/Y _22794_/A VGND VGND VPWR VPWR _22847_/X sky130_fd_sc_hd__o21a_4
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14628__A _12883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12600_ _12617_/A VGND VGND VPWR VPWR _12646_/A sky130_fd_sc_hd__buf_2
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13532__A _13529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20349__B _20348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _13426_/X _13578_/Y _13579_/X VGND VGND VPWR VPWR _13580_/Y sky130_fd_sc_hd__o21ai_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22778_ _16913_/X _18752_/X VGND VGND VPWR VPWR _22778_/Y sky130_fd_sc_hd__nor2_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14347__B _14271_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12531_ _12531_/A VGND VGND VPWR VPWR _15398_/A sky130_fd_sc_hd__buf_2
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21729_ _21572_/X _21726_/X _15266_/B _21723_/X VGND VGND VPWR VPWR _23650_/D sky130_fd_sc_hd__o22a_4
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15250_ _15249_/X VGND VGND VPWR VPWR _15251_/A sky130_fd_sc_hd__inv_2
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18761__C _11620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12462_ _12462_/A _12462_/B VGND VGND VPWR VPWR _12462_/X sky130_fd_sc_hd__or2_4
X_24448_ _24203_/CLK _24448_/D HRESETn VGND VGND VPWR VPWR _20180_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19469__B2 _19433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14201_ _14201_/A _14201_/B _14200_/X VGND VGND VPWR VPWR _14202_/C sky130_fd_sc_hd__or3_4
XFILLER_32_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15181_ _14617_/A _15181_/B _15181_/C VGND VGND VPWR VPWR _15182_/C sky130_fd_sc_hd__and3_4
XANTENNA__15459__A _12585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21276__B2 _21266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12393_ _12826_/A _12285_/B VGND VGND VPWR VPWR _12393_/X sky130_fd_sc_hd__or2_4
X_24379_ _24344_/CLK _24379_/D HRESETn VGND VGND VPWR VPWR _24379_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__24074__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14132_ _11909_/A _14132_/B _14132_/C VGND VGND VPWR VPWR _14136_/B sky130_fd_sc_hd__and3_4
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19873__B _19873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21028__B2 _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14063_ _14031_/A _23466_/Q VGND VGND VPWR VPWR _14063_/X sky130_fd_sc_hd__or2_4
X_18940_ _18940_/A VGND VGND VPWR VPWR _18994_/A sky130_fd_sc_hd__buf_2
XANTENNA__17674__A _17674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21579__A2 _21532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13014_ _13014_/A _13012_/X _13014_/C VGND VGND VPWR VPWR _13014_/X sky130_fd_sc_hd__and3_4
XFILLER_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18871_ _18870_/X VGND VGND VPWR VPWR _18872_/B sky130_fd_sc_hd__buf_2
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_91_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR _24026_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_79_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17822_ _17845_/A VGND VGND VPWR VPWR _17975_/A sky130_fd_sc_hd__buf_2
XFILLER_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21924__A _21938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14965_ _14970_/A _14898_/B VGND VGND VPWR VPWR _14965_/X sky130_fd_sc_hd__or2_4
X_17753_ _17698_/X _17753_/B _17753_/C VGND VGND VPWR VPWR _17753_/X sky130_fd_sc_hd__or3_4
XANTENNA__13426__B _13425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20003__A2 _16945_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13916_ _11670_/A _13908_/X _13916_/C VGND VGND VPWR VPWR _13917_/C sky130_fd_sc_hd__and3_4
X_16704_ _11888_/A _23931_/Q VGND VGND VPWR VPWR _16706_/B sky130_fd_sc_hd__or2_4
XFILLER_48_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21200__B2 _21194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17684_ _17684_/A _17684_/B _17683_/X VGND VGND VPWR VPWR _17684_/X sky130_fd_sc_hd__and3_4
XFILLER_75_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14896_ _14867_/X _23808_/Q VGND VGND VPWR VPWR _14897_/C sky130_fd_sc_hd__or2_4
XFILLER_62_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21751__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21505__A2_N _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16737__B _23707_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16635_ _16622_/A _16635_/B _16634_/X VGND VGND VPWR VPWR _16635_/X sky130_fd_sc_hd__or3_4
X_19423_ _19422_/X VGND VGND VPWR VPWR _19424_/A sky130_fd_sc_hd__buf_2
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13847_ _13847_/A VGND VGND VPWR VPWR _13878_/A sky130_fd_sc_hd__buf_2
XANTENNA__14538__A _13747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13442__A _12466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16566_ _12011_/A _16566_/B _16566_/C VGND VGND VPWR VPWR _16570_/B sky130_fd_sc_hd__and3_4
X_19354_ _19317_/A VGND VGND VPWR VPWR _19370_/A sky130_fd_sc_hd__buf_2
X_13778_ _15393_/A _23495_/Q VGND VGND VPWR VPWR _13778_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15517_ _11656_/A _15485_/X _15516_/X VGND VGND VPWR VPWR _15517_/X sky130_fd_sc_hd__and3_4
X_18305_ _18107_/X _18446_/B _18249_/X _18304_/X VGND VGND VPWR VPWR _18305_/X sky130_fd_sc_hd__a211o_4
X_12729_ _12743_/A VGND VGND VPWR VPWR _12730_/A sky130_fd_sc_hd__buf_2
X_19285_ _19211_/B VGND VGND VPWR VPWR _19285_/Y sky130_fd_sc_hd__inv_2
X_16497_ _16471_/X _16434_/B VGND VGND VPWR VPWR _16497_/X sky130_fd_sc_hd__or2_4
XANTENNA__12058__A _11994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18236_ _17672_/A _18236_/B VGND VGND VPWR VPWR _18237_/A sky130_fd_sc_hd__or2_4
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15448_ _15448_/A _15448_/B _15448_/C VGND VGND VPWR VPWR _15448_/X sky130_fd_sc_hd__and3_4
XFILLER_31_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11897__A _12852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18167_ _17756_/Y _18166_/X _17690_/A VGND VGND VPWR VPWR _18167_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15369__A _13992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21267__B2 _21266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15379_ _11652_/X _15347_/X _15378_/X VGND VGND VPWR VPWR _15379_/X sky130_fd_sc_hd__and3_4
XFILLER_89_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14273__A _13670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17118_ _17115_/Y _17010_/X _17018_/A _17117_/X VGND VGND VPWR VPWR _17150_/A sky130_fd_sc_hd__o22a_4
X_18098_ _23021_/B _18097_/X _23021_/B _18097_/X VGND VGND VPWR VPWR _18098_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15088__B _15088_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22490__A _22483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17049_ _17047_/Y _17049_/B VGND VGND VPWR VPWR _17077_/A sky130_fd_sc_hd__or2_4
XANTENNA__21019__B2 _21013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22216__B1 _15984_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20060_ _20042_/X _18348_/A _20048_/X _20059_/X VGND VGND VPWR VPWR _20060_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13617__A _15435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12521__A _12520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21990__A2 _21988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13336__B _13336_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23750_ _23845_/CLK _21564_/X VGND VGND VPWR VPWR _14276_/B sky130_fd_sc_hd__dfxtp_4
X_20962_ _20223_/A _20960_/X _20961_/X HRDATA[9] _20846_/X VGND VGND VPWR VPWR _20962_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_81_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21742__A2 _21741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22701_ _21555_/A _22700_/X _23081_/Q _22697_/X VGND VGND VPWR VPWR _22701_/X sky130_fd_sc_hd__o22a_4
XFILLER_96_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23681_ _23819_/CLK _21680_/X VGND VGND VPWR VPWR _23681_/Q sky130_fd_sc_hd__dfxtp_4
X_20893_ _21282_/A VGND VGND VPWR VPWR _20893_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14448__A _12862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13352__A _12802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22632_ _22408_/X _22629_/X _12293_/B _22626_/X VGND VGND VPWR VPWR _23126_/D sky130_fd_sc_hd__o22a_4
XFILLER_74_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22563_ _22462_/X _22536_/A _23167_/Q _22518_/X VGND VGND VPWR VPWR _22563_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24302_ _23324_/CLK _19172_/X HRESETn VGND VGND VPWR VPWR _24302_/Q sky130_fd_sc_hd__dfrtp_4
X_21514_ _21799_/A VGND VGND VPWR VPWR _21514_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22494_ _22427_/X _22493_/X _15699_/B _22490_/X VGND VGND VPWR VPWR _23214_/D sky130_fd_sc_hd__o22a_4
XFILLER_10_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24233_ _24203_/CLK _24233_/D HRESETn VGND VGND VPWR VPWR _24233_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15279__A _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21445_ _21291_/X _21440_/X _23808_/Q _21401_/X VGND VGND VPWR VPWR _23808_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18123__A1 _17568_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24359__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21376_ _21369_/A VGND VGND VPWR VPWR _21376_/X sky130_fd_sc_hd__buf_2
X_24164_ _24165_/CLK _24164_/D HRESETn VGND VGND VPWR VPWR _17024_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19871__A1 _19730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20327_ _20497_/A VGND VGND VPWR VPWR _20327_/X sky130_fd_sc_hd__buf_2
X_23115_ _23336_/CLK _23115_/D VGND VGND VPWR VPWR _23115_/Q sky130_fd_sc_hd__dfxtp_4
X_24095_ _24320_/CLK _24095_/D HRESETn VGND VGND VPWR VPWR _18934_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14911__A _15015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_15_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_30_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20258_ _20471_/A VGND VGND VPWR VPWR _20258_/X sky130_fd_sc_hd__buf_2
X_23046_ _23051_/A _23046_/B VGND VGND VPWR VPWR _23046_/X sky130_fd_sc_hd__or2_4
XFILLER_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13527__A _12754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20189_ _21005_/A _19830_/A _19841_/A VGND VGND VPWR VPWR _20199_/A sky130_fd_sc_hd__or3_4
XANTENNA__12431__A _12338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14750_ _13960_/A _14806_/B VGND VGND VPWR VPWR _14751_/C sky130_fd_sc_hd__or2_4
XANTENNA__15742__A _12795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11962_ _16139_/A VGND VGND VPWR VPWR _11962_/X sky130_fd_sc_hd__buf_2
X_23948_ _24044_/CLK _23948_/D VGND VGND VPWR VPWR _15487_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_1_1_1_HCLK clkbuf_1_1_0_HCLK/X VGND VGND VPWR VPWR clkbuf_2_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13701_ _12578_/A VGND VGND VPWR VPWR _15486_/A sky130_fd_sc_hd__buf_2
XFILLER_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14681_ _14664_/X _14679_/X _14681_/C VGND VGND VPWR VPWR _14681_/X sky130_fd_sc_hd__and3_4
X_11893_ _15023_/A VGND VGND VPWR VPWR _11894_/A sky130_fd_sc_hd__buf_2
X_23879_ _23816_/CLK _21336_/X VGND VGND VPWR VPWR _13807_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20941__B1 HRDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16420_ _16400_/A _16489_/B VGND VGND VPWR VPWR _16420_/X sky130_fd_sc_hd__or2_4
XANTENNA__23314__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13262__A _12350_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13632_ _13632_/A VGND VGND VPWR VPWR _15411_/A sky130_fd_sc_hd__buf_2
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16351_ _16365_/A _16283_/B VGND VGND VPWR VPWR _16352_/C sky130_fd_sc_hd__or2_4
X_13563_ _13563_/A _13561_/X _13563_/C VGND VGND VPWR VPWR _13563_/X sky130_fd_sc_hd__and3_4
XANTENNA__21497__B2 _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16573__A _16569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15302_ _11929_/A _15298_/X _15302_/C VGND VGND VPWR VPWR _15302_/X sky130_fd_sc_hd__or3_4
XFILLER_73_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12514_ _13014_/A _12507_/X _12514_/C VGND VGND VPWR VPWR _12514_/X sky130_fd_sc_hd__and3_4
X_19070_ _19060_/X _19069_/X _19060_/X _19065_/A VGND VGND VPWR VPWR _24327_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16282_ _16286_/A _16282_/B VGND VGND VPWR VPWR _16282_/X sky130_fd_sc_hd__or2_4
XFILLER_51_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13494_ _12655_/A VGND VGND VPWR VPWR _13494_/X sky130_fd_sc_hd__buf_2
XFILLER_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18021_ _16931_/X VGND VGND VPWR VPWR _18202_/A sky130_fd_sc_hd__buf_2
XANTENNA__23464__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15233_ _14186_/A _15176_/B VGND VGND VPWR VPWR _15235_/B sky130_fd_sc_hd__or2_4
XANTENNA__15189__A _15201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12445_ _15823_/A _12443_/X _12444_/X VGND VGND VPWR VPWR _12445_/X sky130_fd_sc_hd__and3_4
XANTENNA__19884__A _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14093__A _11879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12606__A _12652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20457__C1 _20456_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15164_ _14098_/A _15162_/X _15163_/X VGND VGND VPWR VPWR _15164_/X sky130_fd_sc_hd__and3_4
XANTENNA__21919__A _21919_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12376_ _12398_/A _12372_/X _12376_/C VGND VGND VPWR VPWR _12376_/X sky130_fd_sc_hd__and3_4
XFILLER_5_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14115_ _14165_/A VGND VGND VPWR VPWR _14143_/A sky130_fd_sc_hd__buf_2
XFILLER_119_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15095_ _14068_/A _23807_/Q VGND VGND VPWR VPWR _15096_/C sky130_fd_sc_hd__or2_4
X_19972_ _19996_/A VGND VGND VPWR VPWR _19972_/X sky130_fd_sc_hd__buf_2
XANTENNA__14821__A _13710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22749__A1 SYSTICKCLKDIV[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14046_ _14046_/A _14044_/X _14046_/C VGND VGND VPWR VPWR _14047_/C sky130_fd_sc_hd__and3_4
X_18923_ _11532_/A VGND VGND VPWR VPWR _18923_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15636__B _23467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13437__A _12518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18854_ _14425_/A _18848_/X _24390_/Q _18849_/X VGND VGND VPWR VPWR _24390_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21421__B2 _21416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17805_ _17802_/X _17146_/X _17804_/X _17162_/X VGND VGND VPWR VPWR _17805_/X sky130_fd_sc_hd__o22a_4
XFILLER_62_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15997_ _15997_/A _23800_/Q VGND VGND VPWR VPWR _15998_/C sky130_fd_sc_hd__or2_4
X_18785_ _13274_/X _18781_/X _24434_/Q _18782_/X VGND VGND VPWR VPWR _18785_/X sky130_fd_sc_hd__o22a_4
XFILLER_62_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16748__A _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15652__A _12221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14948_ _15063_/A _14946_/X _14947_/X VGND VGND VPWR VPWR _14952_/B sky130_fd_sc_hd__and3_4
X_17736_ _17736_/A VGND VGND VPWR VPWR _17737_/A sky130_fd_sc_hd__inv_2
XANTENNA__21185__B1 _23954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21724__A2 _21719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16467__B _16407_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14879_ _11610_/A _14879_/B VGND VGND VPWR VPWR _14881_/B sky130_fd_sc_hd__or2_4
X_17667_ _17667_/A _17667_/B VGND VGND VPWR VPWR _17667_/X sky130_fd_sc_hd__or2_4
XANTENNA__14268__A _12233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13172__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19406_ _19302_/X VGND VGND VPWR VPWR _19406_/X sky130_fd_sc_hd__buf_2
X_16618_ _11758_/X VGND VGND VPWR VPWR _16618_/X sky130_fd_sc_hd__buf_2
XFILLER_91_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17598_ _17395_/X VGND VGND VPWR VPWR _17598_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16549_ _12025_/A VGND VGND VPWR VPWR _16715_/A sky130_fd_sc_hd__buf_2
X_19337_ _19332_/X _18410_/X _19336_/X _24238_/Q VGND VGND VPWR VPWR _24238_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22685__B1 _12823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19268_ _19219_/A _19219_/B _19267_/Y VGND VGND VPWR VPWR _24270_/D sky130_fd_sc_hd__o21a_4
X_18219_ _18216_/X _17444_/X _18217_/X _18082_/X _18218_/Y VGND VGND VPWR VPWR _18219_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15099__A _15107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19794__A _19730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19199_ _19110_/B VGND VGND VPWR VPWR _19199_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12516__A _12892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21230_ _21230_/A VGND VGND VPWR VPWR _21230_/X sky130_fd_sc_hd__buf_2
XANTENNA__21829__A _21817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19853__A1 _19872_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20733__A _20293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16930__B _16929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21161_ _21161_/A VGND VGND VPWR VPWR _21161_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15827__A _12458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21660__B2 _21659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14731__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18203__A _18203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20112_ _20111_/Y _11542_/X _11538_/B VGND VGND VPWR VPWR _20112_/Y sky130_fd_sc_hd__a21oi_4
X_21092_ _20697_/X _21089_/X _15465_/B _21086_/X VGND VGND VPWR VPWR _21092_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19605__A1 _19876_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15546__B _23147_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20043_ _20043_/A VGND VGND VPWR VPWR _20043_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13347__A _12682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21963__A2 _21959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23802_ _23706_/CLK _21461_/X VGND VGND VPWR VPWR _16435_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15562__A _15536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21994_ _21826_/X _21988_/X _23503_/Q _21992_/X VGND VGND VPWR VPWR _21994_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21715__A2 _21712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23733_ _24021_/CLK _21603_/X VGND VGND VPWR VPWR _12586_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_27_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20945_ _20942_/X _20944_/X _20240_/X VGND VGND VPWR VPWR _20945_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20923__B1 _20539_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18592__A1 _18697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ _23157_/CLK _23664_/D VGND VGND VPWR VPWR _23664_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_6_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _20842_/X _20874_/X _20875_/X HRDATA[13] _20847_/X VGND VGND VPWR VPWR _20876_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_39_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22615_ _21784_/A _21917_/B _22383_/C _21060_/A VGND VGND VPWR VPWR _22616_/A sky130_fd_sc_hd__or4_4
XFILLER_35_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21479__B2 _21474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23595_ _24044_/CLK _23595_/D VGND VGND VPWR VPWR _23595_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17703__A2_N _17346_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16393__A _16121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14906__A _14906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13810__A _15429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22140__A2 _22137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22546_ _22432_/X _22543_/X _15462_/B _22540_/X VGND VGND VPWR VPWR _22546_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22477_ _22398_/X _22472_/X _16430_/B _22476_/X VGND VGND VPWR VPWR _22477_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12426__A _15882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12230_ _13017_/A _12228_/X _12230_/C VGND VGND VPWR VPWR _12230_/X sky130_fd_sc_hd__and3_4
X_24216_ _24216_/CLK _24216_/D HRESETn VGND VGND VPWR VPWR _24216_/Q sky130_fd_sc_hd__dfrtp_4
X_21428_ _21261_/X _21426_/X _23821_/Q _21423_/X VGND VGND VPWR VPWR _21428_/X sky130_fd_sc_hd__o22a_4
X_12161_ _11692_/X _12159_/X _12160_/X VGND VGND VPWR VPWR _12161_/X sky130_fd_sc_hd__and3_4
X_24147_ _24250_/CLK _24147_/D HRESETn VGND VGND VPWR VPWR _24147_/Q sky130_fd_sc_hd__dfrtp_4
X_21359_ _21359_/A VGND VGND VPWR VPWR _21359_/X sky130_fd_sc_hd__buf_2
XANTENNA__14641__A _11638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21651__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12092_ _12088_/A _12092_/B _12092_/C VGND VGND VPWR VPWR _12096_/B sky130_fd_sc_hd__and3_4
X_24078_ _24044_/CLK _24078_/D VGND VGND VPWR VPWR _15697_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14360__B _14278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13257__A _13257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15920_ _15518_/X _15650_/Y _15519_/X VGND VGND VPWR VPWR _15920_/Y sky130_fd_sc_hd__o21ai_4
X_23029_ _23018_/A _23027_/Y _23029_/C VGND VGND VPWR VPWR _23029_/X sky130_fd_sc_hd__and3_4
XFILLER_81_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21403__B2 _21402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12161__A _11692_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21954__A2 _21952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15851_ _15889_/A _15851_/B _15851_/C VGND VGND VPWR VPWR _15851_/X sky130_fd_sc_hd__or3_4
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18280__B1 _18082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21474__A _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14802_ _13694_/A _14802_/B VGND VGND VPWR VPWR _14802_/X sky130_fd_sc_hd__or2_4
XANTENNA__15472__A _12638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15782_ _15712_/X _15782_/B VGND VGND VPWR VPWR _15782_/X sky130_fd_sc_hd__and2_4
X_18570_ _18486_/X _18562_/X _18563_/Y _18565_/X _18569_/Y VGND VGND VPWR VPWR _18570_/X
+ sky130_fd_sc_hd__a32o_4
X_12994_ _12993_/X VGND VGND VPWR VPWR _12994_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21706__A2 _21705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14733_ _14756_/A _14733_/B VGND VGND VPWR VPWR _14734_/C sky130_fd_sc_hd__or2_4
X_17521_ _17175_/Y _17515_/Y _18281_/A _17520_/X VGND VGND VPWR VPWR _17521_/X sky130_fd_sc_hd__o22a_4
X_11945_ _11994_/A _11760_/B VGND VGND VPWR VPWR _11945_/X sky130_fd_sc_hd__or2_4
XFILLER_45_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20914__B1 _20913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17386__A2 _17012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17452_ _17181_/X _17525_/B VGND VGND VPWR VPWR _17452_/X sky130_fd_sc_hd__and2_4
X_14664_ _14246_/A VGND VGND VPWR VPWR _14664_/X sky130_fd_sc_hd__buf_2
XFILLER_44_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11876_ _14101_/A VGND VGND VPWR VPWR _14912_/A sky130_fd_sc_hd__buf_2
XFILLER_17_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20818__A _22129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16403_ _16152_/A _16399_/X _16403_/C VGND VGND VPWR VPWR _16403_/X sky130_fd_sc_hd__or3_4
X_13615_ _12475_/A _13703_/B VGND VGND VPWR VPWR _13616_/C sky130_fd_sc_hd__or2_4
X_17383_ _13837_/X VGND VGND VPWR VPWR _17383_/Y sky130_fd_sc_hd__inv_2
X_14595_ _14763_/A _14683_/B VGND VGND VPWR VPWR _14596_/C sky130_fd_sc_hd__or2_4
XFILLER_60_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18335__B2 _18334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16334_ _16364_/A _16259_/B VGND VGND VPWR VPWR _16336_/B sky130_fd_sc_hd__or2_4
X_19122_ _19122_/A _19122_/B VGND VGND VPWR VPWR _19123_/B sky130_fd_sc_hd__and2_4
XANTENNA__13720__A _15495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13546_ _12965_/A VGND VGND VPWR VPWR _13546_/X sky130_fd_sc_hd__buf_2
XFILLER_9_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19053_ _24329_/Q VGND VGND VPWR VPWR _19053_/Y sky130_fd_sc_hd__inv_2
X_16265_ _15937_/X _16263_/X _16264_/X VGND VGND VPWR VPWR _16265_/X sky130_fd_sc_hd__and3_4
XANTENNA__20693__A2 _20679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13477_ _12874_/A VGND VGND VPWR VPWR _13477_/X sky130_fd_sc_hd__buf_2
XANTENNA__21890__B2 _21884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15216_ _14243_/A _15207_/X _15216_/C VGND VGND VPWR VPWR _15217_/C sky130_fd_sc_hd__and3_4
X_18004_ _17651_/B _18003_/X _17647_/X VGND VGND VPWR VPWR _18004_/X sky130_fd_sc_hd__o21a_4
XFILLER_103_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12428_ _12672_/A _12407_/X _12428_/C VGND VGND VPWR VPWR _12429_/C sky130_fd_sc_hd__or3_4
X_16196_ _16227_/A _23543_/Q VGND VGND VPWR VPWR _16196_/X sky130_fd_sc_hd__or2_4
XANTENNA__20553__A _21249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15147_ _14990_/A _23553_/Q VGND VGND VPWR VPWR _15147_/X sky130_fd_sc_hd__or2_4
XANTENNA__15647__A _15646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24342__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12359_ _13243_/A VGND VGND VPWR VPWR _12398_/A sky130_fd_sc_hd__buf_2
XANTENNA__21642__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18023__A _18498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15078_ _15069_/A _23647_/Q VGND VGND VPWR VPWR _15080_/B sky130_fd_sc_hd__or2_4
X_19955_ _16927_/X _19954_/X _17639_/X _19309_/X VGND VGND VPWR VPWR _19955_/X sky130_fd_sc_hd__o22a_4
XFILLER_64_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22198__A2 _22193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14029_ _14847_/A _14029_/B _14028_/X VGND VGND VPWR VPWR _14038_/B sky130_fd_sc_hd__or3_4
X_18906_ _18877_/A VGND VGND VPWR VPWR _18906_/X sky130_fd_sc_hd__buf_2
XANTENNA__13167__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12071__A _12098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19886_ _19885_/Y VGND VGND VPWR VPWR _20644_/A sky130_fd_sc_hd__buf_2
XFILLER_64_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_61_0_HCLK clkbuf_6_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18837_ _12990_/X _18834_/X _20519_/A _18835_/X VGND VGND VPWR VPWR _24403_/D sky130_fd_sc_hd__o22a_4
XANTENNA__18810__A2 _18781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16478__A _16203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24467__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18768_ _18782_/A VGND VGND VPWR VPWR _18768_/X sky130_fd_sc_hd__buf_2
XFILLER_23_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17719_ _18558_/A _17287_/X VGND VGND VPWR VPWR _17723_/B sky130_fd_sc_hd__and2_4
X_18699_ _18698_/X VGND VGND VPWR VPWR _18699_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22370__A2 _22368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19771__B1 _19770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20730_ _20619_/X _20729_/X _20617_/X VGND VGND VPWR VPWR _20730_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20381__A1 _20407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20381__B2 _20253_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20728__A _20358_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20661_ _20518_/X _20660_/X _24333_/Q _20525_/X VGND VGND VPWR VPWR _20661_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14726__A _11894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22400_ _22398_/X _22392_/X _16380_/B _22399_/X VGND VGND VPWR VPWR _22400_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13630__A _13630_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20592_ _20488_/A VGND VGND VPWR VPWR _20592_/X sky130_fd_sc_hd__buf_2
X_23380_ _23635_/CLK _22221_/X VGND VGND VPWR VPWR _23380_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22331_ _15081_/B VGND VGND VPWR VPWR _22331_/X sky130_fd_sc_hd__buf_2
XANTENNA__12246__A _12725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21881__B2 _21877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22262_ _22262_/A VGND VGND VPWR VPWR _22262_/X sky130_fd_sc_hd__buf_2
XANTENNA__20463__A _20463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24001_ _24065_/CLK _24001_/D VGND VGND VPWR VPWR _15196_/B sky130_fd_sc_hd__dfxtp_4
X_21213_ _21213_/A VGND VGND VPWR VPWR _21634_/D sky130_fd_sc_hd__buf_2
XANTENNA__15557__A _15571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22193_ _22153_/A VGND VGND VPWR VPWR _22193_/X sky130_fd_sc_hd__buf_2
XFILLER_82_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21144_ _21130_/A VGND VGND VPWR VPWR _21144_/X sky130_fd_sc_hd__buf_2
XANTENNA__15312__A1 _11841_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22189__A2 _22186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21075_ _21075_/A VGND VGND VPWR VPWR _21075_/X sky130_fd_sc_hd__buf_2
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19690__C _19877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20026_ _18338_/X _20009_/X _20025_/Y _20020_/X VGND VGND VPWR VPWR _20026_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16388__A _15997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15292__A _14158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13805__A _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21149__B1 _13630_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24137__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13524__B _13456_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19699__A HRDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21977_ _21797_/X _21974_/X _23515_/Q _21971_/X VGND VGND VPWR VPWR _23515_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17368__A2 _17340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11729_/X VGND VGND VPWR VPWR _11730_/X sky130_fd_sc_hd__buf_2
X_23716_ _23363_/CLK _23716_/D VGND VGND VPWR VPWR _14654_/B sky130_fd_sc_hd__dfxtp_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ _20733_/X _20927_/X _19092_/A _20453_/A VGND VGND VPWR VPWR _20928_/X sky130_fd_sc_hd__o22a_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23014__A _22985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11661_/A VGND VGND VPWR VPWR _14039_/A sky130_fd_sc_hd__buf_2
X_23647_ _23487_/CLK _21732_/X VGND VGND VPWR VPWR _23647_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20859_ _20704_/X _20858_/Y _24261_/Q _20325_/X VGND VGND VPWR VPWR _20859_/X sky130_fd_sc_hd__o22a_4
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14636__A _13611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _13370_/A _13400_/B _13400_/C VGND VGND VPWR VPWR _13408_/B sky130_fd_sc_hd__or3_4
XANTENNA__13540__A _15884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17012__A _17012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ _15607_/A _14378_/X _14380_/C VGND VGND VPWR VPWR _14380_/X sky130_fd_sc_hd__and3_4
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ _11592_/A VGND VGND VPWR VPWR _11592_/X sky130_fd_sc_hd__buf_2
X_23578_ _23699_/CLK _21878_/X VGND VGND VPWR VPWR _16405_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14355__B _14275_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ _12503_/A _13327_/X _13330_/X VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__or3_4
XANTENNA__20076__C _18940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22529_ _22536_/A VGND VGND VPWR VPWR _22529_/X sky130_fd_sc_hd__buf_2
Xclkbuf_2_1_0_HCLK clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ _16050_/A _24056_/Q VGND VGND VPWR VPWR _16051_/C sky130_fd_sc_hd__or2_4
X_13262_ _12350_/A _13262_/B _13262_/C VGND VGND VPWR VPWR _13266_/B sky130_fd_sc_hd__and3_4
XANTENNA__15551__A1 _13597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20373__A _21799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15001_ _15028_/A _15001_/B _15000_/X VGND VGND VPWR VPWR _15002_/C sky130_fd_sc_hd__and3_4
X_12213_ _13046_/A _12213_/B VGND VGND VPWR VPWR _12213_/X sky130_fd_sc_hd__or2_4
XFILLER_87_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15467__A _12646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13193_ _12745_/A _13193_/B VGND VGND VPWR VPWR _13193_/X sky130_fd_sc_hd__or2_4
XFILLER_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21624__B2 _21623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23502__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20832__C1 _20831_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12144_ _12168_/A _23997_/Q VGND VGND VPWR VPWR _12145_/C sky130_fd_sc_hd__or2_4
XFILLER_29_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19740_ _19740_/A _19740_/B VGND VGND VPWR VPWR _19740_/X sky130_fd_sc_hd__or2_4
XFILLER_110_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12075_ _11994_/A _23581_/Q VGND VGND VPWR VPWR _12076_/C sky130_fd_sc_hd__or2_4
X_16952_ _16952_/A VGND VGND VPWR VPWR _17694_/A sky130_fd_sc_hd__inv_2
XFILLER_96_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21927__A2 _21924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15903_ _13511_/X _15901_/X _15903_/C VGND VGND VPWR VPWR _15904_/C sky130_fd_sc_hd__and3_4
XFILLER_81_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18253__B1 _18189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19671_ _19722_/A VGND VGND VPWR VPWR _19672_/C sky130_fd_sc_hd__buf_2
X_16883_ _12996_/B _16899_/B _12993_/X VGND VGND VPWR VPWR _16883_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16298__A _15937_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18622_ _17295_/X _18620_/X _18063_/A _18621_/X VGND VGND VPWR VPWR _18623_/A sky130_fd_sc_hd__a211o_4
XFILLER_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15834_ _12914_/A _15834_/B _15834_/C VGND VGND VPWR VPWR _15834_/X sky130_fd_sc_hd__or3_4
XFILLER_49_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18553_ _18512_/X _18552_/X _24456_/Q _18512_/X VGND VGND VPWR VPWR _24456_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12977_ _12953_/A _23859_/Q VGND VGND VPWR VPWR _12978_/C sky130_fd_sc_hd__or2_4
X_15765_ _12792_/A _15765_/B VGND VGND VPWR VPWR _15765_/X sky130_fd_sc_hd__or2_4
XFILLER_20_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22352__A2 _22347_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17504_ _13202_/X VGND VGND VPWR VPWR _17504_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15930__A _15929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11928_ _14752_/A VGND VGND VPWR VPWR _11929_/A sky130_fd_sc_hd__buf_2
X_14716_ _14397_/A _14712_/X _14716_/C VGND VGND VPWR VPWR _14716_/X sky130_fd_sc_hd__or3_4
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15696_ _15696_/A _15769_/B VGND VGND VPWR VPWR _15696_/X sky130_fd_sc_hd__or2_4
X_18484_ _18484_/A VGND VGND VPWR VPWR _18484_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14647_ _15114_/A _14645_/X _14647_/C VGND VGND VPWR VPWR _14656_/B sky130_fd_sc_hd__and3_4
X_17435_ _18428_/A _17433_/X _17434_/Y VGND VGND VPWR VPWR _17435_/X sky130_fd_sc_hd__o21a_4
X_11859_ _11859_/A VGND VGND VPWR VPWR _13004_/A sky130_fd_sc_hd__buf_2
XFILLER_21_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22104__A2 _22101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ _14145_/A _14578_/B _14577_/X VGND VGND VPWR VPWR _14578_/X sky130_fd_sc_hd__or3_4
X_17366_ _16800_/A _17364_/X _17365_/X VGND VGND VPWR VPWR _17367_/B sky130_fd_sc_hd__o21a_4
XFILLER_20_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24158__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19105_ _24351_/Q _19084_/X VGND VGND VPWR VPWR _19105_/Y sky130_fd_sc_hd__nor2_4
XFILLER_14_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13529_ _12967_/A VGND VGND VPWR VPWR _13529_/X sky130_fd_sc_hd__buf_2
X_16317_ _16322_/A _24025_/Q VGND VGND VPWR VPWR _16317_/X sky130_fd_sc_hd__or2_4
X_17297_ _14719_/X VGND VGND VPWR VPWR _17297_/X sky130_fd_sc_hd__buf_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16761__A _11834_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16248_ _16145_/A _16248_/B VGND VGND VPWR VPWR _16248_/X sky130_fd_sc_hd__or2_4
X_19036_ _19030_/X _19035_/X _19030_/X _24333_/Q VGND VGND VPWR VPWR _24333_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20283__A _20421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15377__A _13991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16179_ _16229_/A _16172_/X _16179_/C VGND VGND VPWR VPWR _16180_/C sky130_fd_sc_hd__or3_4
XANTENNA__21615__B2 _21609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18087__A3 _18080_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21091__A2 _21089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19938_ _18603_/Y _20176_/A VGND VGND VPWR VPWR _20057_/A sky130_fd_sc_hd__or2_4
XFILLER_114_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21379__B1 _23852_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22040__B2 _22035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19869_ _19867_/X _19868_/X _19881_/A VGND VGND VPWR VPWR _19869_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_99_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18200__B _18174_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21900_ _21838_/X _21894_/X _23562_/Q _21898_/X VGND VGND VPWR VPWR _23562_/D sky130_fd_sc_hd__o22a_4
XFILLER_96_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13625__A _13813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22591__A2 _22586_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22880_ _12031_/B _22827_/X _19887_/X _22879_/X VGND VGND VPWR VPWR _22881_/B sky130_fd_sc_hd__o22a_4
XFILLER_7_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16001__A _13477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22938__A _22978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24230__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21831_ _21831_/A VGND VGND VPWR VPWR _21831_/X sky130_fd_sc_hd__buf_2
XANTENNA__22879__B1 _15713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15840__A _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19312__A _19933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21762_ _21755_/A VGND VGND VPWR VPWR _21762_/X sky130_fd_sc_hd__buf_2
XFILLER_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_68_0_HCLK clkbuf_6_34_0_HCLK/X VGND VGND VPWR VPWR _24321_/CLK sky130_fd_sc_hd__clkbuf_1
X_23501_ _23826_/CLK _21997_/X VGND VGND VPWR VPWR _23501_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20713_ _20518_/X _20712_/X _24331_/Q _20525_/X VGND VGND VPWR VPWR _20713_/X sky130_fd_sc_hd__o22a_4
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21693_ _21510_/X _21691_/X _23676_/Q _21688_/X VGND VGND VPWR VPWR _23676_/D sky130_fd_sc_hd__o22a_4
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23432_ _23304_/CLK _22128_/X VGND VGND VPWR VPWR _13729_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20644_ _20644_/A _22855_/A VGND VGND VPWR VPWR _20644_/X sky130_fd_sc_hd__or2_4
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21854__A1 _21852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23363_ _23363_/CLK _23363_/D VGND VGND VPWR VPWR _14765_/B sky130_fd_sc_hd__dfxtp_4
X_20575_ _20511_/X _20574_/X _24081_/Q _20488_/X VGND VGND VPWR VPWR _20575_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16671__A _16640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21854__B2 _21848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22314_ _13304_/B VGND VGND VPWR VPWR _22314_/X sky130_fd_sc_hd__buf_2
XANTENNA__21289__A _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23294_ _23326_/CLK _23294_/D VGND VGND VPWR VPWR _11760_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16390__B _16390_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14903__B _14903_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15287__A _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21606__A1 _21531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22245_ _22139_/X _22243_/X _14765_/B _22240_/X VGND VGND VPWR VPWR _23363_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21606__B2 _21602_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14191__A _11738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12704__A _15693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22176_ _22169_/A VGND VGND VPWR VPWR _22176_/X sky130_fd_sc_hd__buf_2
XANTENNA__12423__B _12323_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24389__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21127_ _20419_/X _21126_/X _23992_/Q _21123_/X VGND VGND VPWR VPWR _21127_/X sky130_fd_sc_hd__o22a_4
XFILLER_87_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21909__A2 _21908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21058_ _24030_/Q VGND VGND VPWR VPWR _21058_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18786__A1 _13270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12900_ _12528_/A _12896_/X _12900_/C VGND VGND VPWR VPWR _12900_/X sky130_fd_sc_hd__or3_4
XFILLER_101_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22582__A2 _22579_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20009_ _19985_/A VGND VGND VPWR VPWR _20009_/X sky130_fd_sc_hd__buf_2
XFILLER_47_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13880_ _13880_/A _13880_/B _13879_/X VGND VGND VPWR VPWR _13884_/B sky130_fd_sc_hd__and3_4
XANTENNA__20593__A1 _20511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20593__B2 _20592_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12831_ _12753_/X _12831_/B _12830_/X VGND VGND VPWR VPWR _12831_/X sky130_fd_sc_hd__or3_4
XFILLER_41_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21752__A _21752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15550_ _12269_/A _15549_/X VGND VGND VPWR VPWR _15550_/X sky130_fd_sc_hd__and2_4
X_12762_ _12816_/A _23508_/Q VGND VGND VPWR VPWR _12763_/C sky130_fd_sc_hd__or2_4
XFILLER_61_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20368__A _24250_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14500_/X _14501_/B VGND VGND VPWR VPWR _14501_/X sky130_fd_sc_hd__or2_4
XANTENNA__17210__A1 _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _12381_/A VGND VGND VPWR VPWR _11713_/X sky130_fd_sc_hd__buf_2
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15512_/A _15410_/B VGND VGND VPWR VPWR _15481_/X sky130_fd_sc_hd__or2_4
XFILLER_54_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _24020_/Q VGND VGND VPWR VPWR _12695_/B sky130_fd_sc_hd__or2_4
XFILLER_70_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14366__A _11766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14432_/A _14497_/B VGND VGND VPWR VPWR _14433_/C sky130_fd_sc_hd__or2_4
X_17220_ _17220_/A VGND VGND VPWR VPWR _17825_/A sky130_fd_sc_hd__buf_2
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11644_/A VGND VGND VPWR VPWR _11645_/A sky130_fd_sc_hd__buf_2
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19876__B _19876_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22583__A _22583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17151_ _17220_/A VGND VGND VPWR VPWR _17151_/X sky130_fd_sc_hd__buf_2
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _15607_/A _14360_/X _14362_/X VGND VGND VPWR VPWR _14364_/C sky130_fd_sc_hd__and3_4
XFILLER_50_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11575_ _11538_/X _11548_/X _20089_/D _20071_/A VGND VGND VPWR VPWR _20070_/A sky130_fd_sc_hd__or4_4
XFILLER_10_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16102_ _16146_/A VGND VGND VPWR VPWR _16108_/A sky130_fd_sc_hd__buf_2
XANTENNA__18710__A1 _18011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13314_ _13317_/A _13310_/X _13313_/X VGND VGND VPWR VPWR _13314_/X sky130_fd_sc_hd__or3_4
XANTENNA__24450__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17082_ _17083_/B _17082_/B VGND VGND VPWR VPWR _17084_/A sky130_fd_sc_hd__and2_4
X_14294_ _15448_/A _14292_/X _14294_/C VGND VGND VPWR VPWR _14298_/B sky130_fd_sc_hd__and3_4
XANTENNA__15909__B _15909_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16033_ _16064_/A _15967_/B VGND VGND VPWR VPWR _16035_/B sky130_fd_sc_hd__or2_4
X_13245_ _13228_/A _13178_/B VGND VGND VPWR VPWR _13247_/B sky130_fd_sc_hd__or2_4
XANTENNA__15197__A _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18474__B1 _18048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13176_ _15687_/A _13174_/X _13176_/C VGND VGND VPWR VPWR _13176_/X sky130_fd_sc_hd__and3_4
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22270__B2 _22269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11561__A2 IRQ[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12127_ _11685_/X _12121_/X _12127_/C VGND VGND VPWR VPWR _12127_/X sky130_fd_sc_hd__or3_4
X_17984_ _17975_/X _17935_/X _17798_/X _17983_/X VGND VGND VPWR VPWR _17984_/X sky130_fd_sc_hd__o22a_4
XFILLER_2_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19723_ _19857_/C _19723_/B VGND VGND VPWR VPWR _19723_/X sky130_fd_sc_hd__and2_4
X_12058_ _11994_/A VGND VGND VPWR VPWR _12091_/A sky130_fd_sc_hd__buf_2
X_16935_ _16935_/A VGND VGND VPWR VPWR _16935_/X sky130_fd_sc_hd__buf_2
XANTENNA__18777__A1 _17164_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22573__A2 _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19654_ _19516_/A VGND VGND VPWR VPWR _19726_/B sky130_fd_sc_hd__inv_2
X_16866_ _16865_/X VGND VGND VPWR VPWR _16870_/B sky130_fd_sc_hd__inv_2
XFILLER_65_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18605_ _11628_/X VGND VGND VPWR VPWR _18605_/X sky130_fd_sc_hd__buf_2
XANTENNA__21662__A _21662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15817_ _12851_/A _15879_/B VGND VGND VPWR VPWR _15819_/B sky130_fd_sc_hd__or2_4
XFILLER_0_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19585_ _19419_/A VGND VGND VPWR VPWR _19585_/X sky130_fd_sc_hd__buf_2
X_16797_ _16768_/X _23803_/Q VGND VGND VPWR VPWR _16797_/X sky130_fd_sc_hd__or2_4
XANTENNA__16756__A _11823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18529__B2 _18528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15660__A _12286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18536_ _18536_/A VGND VGND VPWR VPWR _18536_/Y sky130_fd_sc_hd__inv_2
X_15748_ _13130_/A _15748_/B VGND VGND VPWR VPWR _15748_/X sky130_fd_sc_hd__or2_4
XFILLER_61_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18467_ _18421_/A _17349_/Y VGND VGND VPWR VPWR _18468_/D sky130_fd_sc_hd__and2_4
XFILLER_72_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15679_ _12713_/A _15679_/B _15678_/X VGND VGND VPWR VPWR _15679_/X sky130_fd_sc_hd__or3_4
XANTENNA__14276__A _12260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18971__A _18971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17752__A2 _17354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17418_ _14261_/X _17427_/B VGND VGND VPWR VPWR _17418_/X sky130_fd_sc_hd__or2_4
X_18398_ _18713_/A VGND VGND VPWR VPWR _18398_/X sky130_fd_sc_hd__buf_2
XFILLER_53_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17349_ _17349_/A VGND VGND VPWR VPWR _17349_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20360_ _20578_/A VGND VGND VPWR VPWR _20502_/A sky130_fd_sc_hd__buf_2
XANTENNA__14723__B _14723_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19019_ _11520_/B VGND VGND VPWR VPWR _19019_/Y sky130_fd_sc_hd__inv_2
X_20291_ _20467_/A VGND VGND VPWR VPWR _20291_/X sky130_fd_sc_hd__buf_2
XANTENNA__12524__A _12915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22030_ _21802_/X _22024_/X _23481_/Q _22028_/X VGND VGND VPWR VPWR _23481_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22261__B2 _22255_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11552__A2 IRQ[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15835__A _12879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22013__B2 _21970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23981_ _23698_/CLK _23981_/D VGND VGND VPWR VPWR _15799_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_31_0_HCLK clkbuf_5_30_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22932_ _22932_/A _22932_/B VGND VGND VPWR VPWR _22932_/Y sky130_fd_sc_hd__nand2_4
XFILLER_99_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20575__A1 _20511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22668__A _22683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20575__B2 _20488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18865__B _12096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22863_ _22779_/X VGND VGND VPWR VPWR _22863_/X sky130_fd_sc_hd__buf_2
XANTENNA__19717__B1 _12100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15570__A _14463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21814_ _20509_/A VGND VGND VPWR VPWR _21814_/X sky130_fd_sc_hd__buf_2
XFILLER_37_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22794_ _22794_/A VGND VGND VPWR VPWR _22794_/X sky130_fd_sc_hd__buf_2
XFILLER_38_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21745_ _21737_/X VGND VGND VPWR VPWR _21745_/X sky130_fd_sc_hd__buf_2
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24464_ _24066_/CLK _18339_/X HRESETn VGND VGND VPWR VPWR _20025_/A sky130_fd_sc_hd__dfrtp_4
X_21676_ _21636_/A VGND VGND VPWR VPWR _21676_/X sky130_fd_sc_hd__buf_2
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12418__B _12312_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23415_ _23383_/CLK _23415_/D VGND VGND VPWR VPWR _16135_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21827__A1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20627_ _20622_/X _20626_/X _19219_/A _20497_/X VGND VGND VPWR VPWR _20627_/X sky130_fd_sc_hd__o22a_4
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24395_ _24365_/CLK _24395_/D HRESETn VGND VGND VPWR VPWR _24395_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21827__B2 _21824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23346_ _23826_/CLK _23346_/D VGND VGND VPWR VPWR _13069_/B sky130_fd_sc_hd__dfxtp_4
X_20558_ _20558_/A VGND VGND VPWR VPWR _20558_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23277_ _23122_/CLK _23277_/D VGND VGND VPWR VPWR _15795_/B sky130_fd_sc_hd__dfxtp_4
X_20489_ _20396_/X _20487_/X _24085_/Q _20488_/X VGND VGND VPWR VPWR _20489_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13030_ _12887_/A _13028_/X _13030_/C VGND VGND VPWR VPWR _13030_/X sky130_fd_sc_hd__and3_4
X_22228_ _22110_/X _22222_/X _13552_/B _22226_/X VGND VGND VPWR VPWR _23375_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21055__A2 _21051_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15745__A _13102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22159_ _22075_/X _22158_/X _23421_/Q _22155_/X VGND VGND VPWR VPWR _23421_/D sky130_fd_sc_hd__o22a_4
XFILLER_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22004__A1 _21843_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22004__B2 _21999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14981_ _11709_/A _23616_/Q VGND VGND VPWR VPWR _14982_/C sky130_fd_sc_hd__or2_4
XANTENNA__22555__A2 _22550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16720_ _16713_/A _16788_/B VGND VGND VPWR VPWR _16720_/X sky130_fd_sc_hd__or2_4
XFILLER_102_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13265__A _13243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13932_ _13611_/A _13932_/B _13932_/C VGND VGND VPWR VPWR _13933_/C sky130_fd_sc_hd__and3_4
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21763__B1 _15700_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13863_ _13879_/A _13863_/B VGND VGND VPWR VPWR _13864_/C sky130_fd_sc_hd__or2_4
X_16651_ _16651_/A _24060_/Q VGND VGND VPWR VPWR _16652_/C sky130_fd_sc_hd__or2_4
XFILLER_78_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16576__A _12011_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17982__A2 _17848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19708__B1 _19704_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12814_ _12771_/X _12814_/B _12814_/C VGND VGND VPWR VPWR _12822_/B sky130_fd_sc_hd__or3_4
X_15602_ _15633_/A _23435_/Q VGND VGND VPWR VPWR _15603_/C sky130_fd_sc_hd__or2_4
X_19370_ _19370_/A VGND VGND VPWR VPWR _19370_/X sky130_fd_sc_hd__buf_2
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21167__A2_N _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13794_ _13794_/A _13794_/B VGND VGND VPWR VPWR _13796_/B sky130_fd_sc_hd__or2_4
X_16582_ _16686_/A _16672_/B VGND VGND VPWR VPWR _16582_/X sky130_fd_sc_hd__or2_4
XFILLER_56_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18321_ _18267_/A _18321_/B _18319_/X _18321_/D VGND VGND VPWR VPWR _18322_/A sky130_fd_sc_hd__or4_4
X_12745_ _12745_/A _12827_/B VGND VGND VPWR VPWR _12745_/X sky130_fd_sc_hd__or2_4
X_15533_ _15533_/A _23275_/Q VGND VGND VPWR VPWR _15533_/X sky130_fd_sc_hd__or2_4
XANTENNA__19887__A _22824_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14096__A _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12609__A _12964_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16821__A1_N _16897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_51_0_HCLK clkbuf_7_50_0_HCLK/A VGND VGND VPWR VPWR _23304_/CLK sky130_fd_sc_hd__clkbuf_1
X_15464_ _13765_/A _15462_/X _15463_/X VGND VGND VPWR VPWR _15464_/X sky130_fd_sc_hd__and3_4
X_18252_ _18107_/X _18248_/Y _18249_/X _18251_/Y VGND VGND VPWR VPWR _18252_/X sky130_fd_sc_hd__a211o_4
X_12676_ _12675_/Y VGND VGND VPWR VPWR _12676_/X sky130_fd_sc_hd__buf_2
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__A1 _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _15637_/A _14320_/B VGND VGND VPWR VPWR _14415_/X sky130_fd_sc_hd__or2_4
X_17203_ _12992_/X _17173_/X _17172_/Y _17145_/X VGND VGND VPWR VPWR _17203_/X sky130_fd_sc_hd__o22a_4
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _22888_/A _11626_/Y VGND VGND VPWR VPWR _20077_/D sky130_fd_sc_hd__or2_4
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23840__CLK _23840_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21818__A1 _21816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15395_ _13614_/A _15458_/B VGND VGND VPWR VPWR _15397_/B sky130_fd_sc_hd__or2_4
X_18183_ _17256_/A VGND VGND VPWR VPWR _18183_/X sky130_fd_sc_hd__buf_2
XFILLER_15_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21818__B2 _21812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14824__A _14050_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19487__A2 _19481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17498__A1 _13059_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ _14359_/A VGND VGND VPWR VPWR _15586_/A sky130_fd_sc_hd__buf_2
X_17134_ _15251_/X _17131_/X _17132_/Y _17133_/X VGND VGND VPWR VPWR _17134_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ _11558_/A _11558_/B VGND VGND VPWR VPWR _11559_/B sky130_fd_sc_hd__or2_4
XANTENNA__17498__B2 _17497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21294__A2 _21247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22491__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15639__B _23211_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17065_ _17157_/A VGND VGND VPWR VPWR _17065_/X sky130_fd_sc_hd__buf_2
X_14277_ _13670_/A _14275_/X _14276_/X VGND VGND VPWR VPWR _14277_/X sky130_fd_sc_hd__and3_4
XFILLER_116_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12344__A _12826_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16016_ _16047_/A _23736_/Q VGND VGND VPWR VPWR _16016_/X sky130_fd_sc_hd__or2_4
X_13228_ _13228_/A _13153_/B VGND VGND VPWR VPWR _13231_/B sky130_fd_sc_hd__or2_4
XANTENNA__21046__A2 _21044_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_14_0_HCLK_A clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15655__A _12284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13159_ _15697_/A _23537_/Q VGND VGND VPWR VPWR _13159_/X sky130_fd_sc_hd__or2_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23220__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17967_ _17966_/X VGND VGND VPWR VPWR _18142_/A sky130_fd_sc_hd__buf_2
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22546__A2 _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19706_ _19706_/A _19669_/Y VGND VGND VPWR VPWR _19706_/X sky130_fd_sc_hd__and2_4
XANTENNA__13175__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16918_ _11632_/X _11634_/X _16918_/C VGND VGND VPWR VPWR _16923_/A sky130_fd_sc_hd__or3_4
XFILLER_61_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17898_ _17766_/A _17896_/X _16939_/A _17897_/Y VGND VGND VPWR VPWR _17898_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21754__B1 _12836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19637_ _19637_/A VGND VGND VPWR VPWR _19637_/Y sky130_fd_sc_hd__inv_2
X_16849_ _15914_/D _16838_/X _15909_/X VGND VGND VPWR VPWR _16850_/B sky130_fd_sc_hd__o21a_4
XANTENNA__19701__A1_N _19674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13903__A _13879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19568_ _24146_/Q _19435_/X HRDATA[20] _19432_/X VGND VGND VPWR VPWR _19568_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18519_ _17966_/X _18491_/X _17966_/X _18488_/X VGND VGND VPWR VPWR _18519_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13622__B _24008_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19499_ _19499_/A VGND VGND VPWR VPWR _19499_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17725__A2 _17290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12519__A _12518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21530_ _21529_/X _21520_/X _12774_/B _21527_/X VGND VGND VPWR VPWR _21530_/X sky130_fd_sc_hd__o22a_4
XFILLER_90_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20736__A _20497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21461_ _21229_/X _21456_/X _16435_/B _21460_/X VGND VGND VPWR VPWR _21461_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18206__A _18206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23200_ _23233_/CLK _22512_/X VGND VGND VPWR VPWR _14905_/B sky130_fd_sc_hd__dfxtp_4
X_20412_ _20502_/A _20411_/X VGND VGND VPWR VPWR _20412_/Y sky130_fd_sc_hd__nor2_4
X_24180_ _24180_/CLK _19709_/X HRESETn VGND VGND VPWR VPWR _12529_/A sky130_fd_sc_hd__dfrtp_4
X_21392_ _21285_/X _21390_/X _14780_/B _21387_/X VGND VGND VPWR VPWR _23843_/D sky130_fd_sc_hd__o22a_4
XFILLER_107_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22951__A _18475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23131_ _24059_/CLK _23131_/D VGND VGND VPWR VPWR _16788_/B sky130_fd_sc_hd__dfxtp_4
X_20343_ _20229_/X _20342_/X _20213_/X VGND VGND VPWR VPWR _20343_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_49_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12254__A _13670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23062_ _23062_/A VGND VGND VPWR VPWR _23062_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18438__B1 _18016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20274_ _18577_/Y VGND VGND VPWR VPWR _20484_/A sky130_fd_sc_hd__buf_2
XANTENNA__22234__B2 _22233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22013_ _21859_/X _22009_/X _15126_/B _21970_/X VGND VGND VPWR VPWR _22013_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18453__A3 _18447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19650__A2 HRDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18876__A _18898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22537__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23964_ _23515_/CLK _23964_/D VGND VGND VPWR VPWR _23964_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23713__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22398__A _20372_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22915_ _23038_/B VGND VGND VPWR VPWR _22945_/B sky130_fd_sc_hd__buf_2
XFILLER_29_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19953__A3 _19947_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23895_ _23632_/CLK _23895_/D VGND VGND VPWR VPWR _16124_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24319__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13813__A _13813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22846_ _22846_/A VGND VGND VPWR VPWR HWDATA[21] sky130_fd_sc_hd__inv_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22777_ _22777_/A VGND VGND VPWR VPWR _22777_/X sky130_fd_sc_hd__buf_2
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12429__A _11657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12530_ _15032_/A VGND VGND VPWR VPWR _12531_/A sky130_fd_sc_hd__buf_2
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_38_0_HCLK clkbuf_6_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_38_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21728_ _21570_/X _21726_/X _14739_/B _21723_/X VGND VGND VPWR VPWR _21728_/X sky130_fd_sc_hd__o22a_4
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23022__A _18124_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12461_ _12891_/A VGND VGND VPWR VPWR _12528_/A sky130_fd_sc_hd__buf_2
X_24447_ _24203_/CLK _24447_/D HRESETn VGND VGND VPWR VPWR _24447_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18761__D _18812_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21659_ _21659_/A VGND VGND VPWR VPWR _21659_/X sky130_fd_sc_hd__buf_2
X_14200_ _14215_/A _14200_/B _14200_/C VGND VGND VPWR VPWR _14200_/X sky130_fd_sc_hd__and3_4
XFILLER_21_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15180_ _14151_/A _15180_/B VGND VGND VPWR VPWR _15181_/C sky130_fd_sc_hd__or2_4
XANTENNA__18677__B1 _17779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21276__A2 _21271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12392_ _12392_/A VGND VGND VPWR VPWR _12672_/A sky130_fd_sc_hd__buf_2
X_24378_ _24344_/CLK _24378_/D HRESETn VGND VGND VPWR VPWR _18954_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__22473__B2 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15459__B _15459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14131_ _11954_/A _23945_/Q VGND VGND VPWR VPWR _14132_/C sky130_fd_sc_hd__or2_4
X_23329_ _23104_/CLK _23329_/D VGND VGND VPWR VPWR _15128_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17955__A _18205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14062_ _14037_/A _14062_/B _14062_/C VGND VGND VPWR VPWR _14062_/X sky130_fd_sc_hd__or3_4
XANTENNA__18429__B1 _18048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21477__A _21470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17674__B _17506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22225__B2 _22219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13013_ _13032_/A _23986_/Q VGND VGND VPWR VPWR _13014_/C sky130_fd_sc_hd__or2_4
XANTENNA__15475__A _13087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18870_ _20407_/A VGND VGND VPWR VPWR _18870_/X sky130_fd_sc_hd__buf_2
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20787__A1 _20622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21984__B1 _12213_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17821_ _17800_/X _17810_/Y _17812_/X _17820_/Y VGND VGND VPWR VPWR _17821_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22528__A2 _22522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17752_ _16974_/A _17354_/X _17701_/X _17751_/X VGND VGND VPWR VPWR _17753_/C sky130_fd_sc_hd__o22a_4
XANTENNA__23393__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14964_ _15063_/A _14962_/X _14964_/C VGND VGND VPWR VPWR _14968_/B sky130_fd_sc_hd__and3_4
XFILLER_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16703_ _12096_/A _16703_/B _16703_/C VGND VGND VPWR VPWR _16703_/X sky130_fd_sc_hd__or3_4
X_13915_ _11740_/A _13915_/B _13915_/C VGND VGND VPWR VPWR _13916_/C sky130_fd_sc_hd__or3_4
XANTENNA__21200__A2 _21197_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17683_ _17677_/X _17678_/X _18286_/A VGND VGND VPWR VPWR _17683_/X sky130_fd_sc_hd__or3_4
XFILLER_47_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14895_ _14895_/A _14962_/B VGND VGND VPWR VPWR _14895_/X sky130_fd_sc_hd__or2_4
XANTENNA__22101__A _22101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14819__A _13872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19422_ _19458_/A VGND VGND VPWR VPWR _19422_/X sky130_fd_sc_hd__buf_2
X_16634_ _16652_/A _16634_/B _16634_/C VGND VGND VPWR VPWR _16634_/X sky130_fd_sc_hd__and3_4
X_13846_ _13896_/A _13846_/B _13846_/C VGND VGND VPWR VPWR _13846_/X sky130_fd_sc_hd__and3_4
XFILLER_63_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19353_ _19350_/X _18687_/X _19350_/X _20932_/A VGND VGND VPWR VPWR _19353_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13777_ _15392_/A _13841_/B VGND VGND VPWR VPWR _13777_/X sky130_fd_sc_hd__or2_4
X_16565_ _16565_/A _23964_/Q VGND VGND VPWR VPWR _16566_/C sky130_fd_sc_hd__or2_4
XFILLER_108_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12339__A _11645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22161__B1 _16792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18904__A1 _15646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18304_ _18425_/A _18304_/B VGND VGND VPWR VPWR _18304_/X sky130_fd_sc_hd__and2_4
X_15516_ _12392_/A _15516_/B _15515_/X VGND VGND VPWR VPWR _15516_/X sky130_fd_sc_hd__or3_4
XFILLER_56_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12728_ _12728_/A _23380_/Q VGND VGND VPWR VPWR _12728_/X sky130_fd_sc_hd__or2_4
X_19284_ _19211_/A _19211_/B _19283_/Y VGND VGND VPWR VPWR _19284_/X sky130_fd_sc_hd__o21a_4
X_16496_ _11770_/X _16488_/X _16496_/C VGND VGND VPWR VPWR _16496_/X sky130_fd_sc_hd__and3_4
XANTENNA__20556__A _20556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18235_ _18235_/A VGND VGND VPWR VPWR _18236_/B sky130_fd_sc_hd__inv_2
XFILLER_50_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12659_ _12963_/A _12657_/X _12659_/C VGND VGND VPWR VPWR _12663_/B sky130_fd_sc_hd__and3_4
X_15447_ _15447_/A _23852_/Q VGND VGND VPWR VPWR _15448_/C sky130_fd_sc_hd__or2_4
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18026__A _18295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21267__A2 _21259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18166_ _17669_/X _18165_/X _17686_/X VGND VGND VPWR VPWR _18166_/X sky130_fd_sc_hd__o21a_4
X_15378_ _11797_/A _15362_/X _15378_/C VGND VGND VPWR VPWR _15378_/X sky130_fd_sc_hd__or3_4
XFILLER_102_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17117_ _13048_/A _17105_/X _19841_/A _17032_/B VGND VGND VPWR VPWR _17117_/X sky130_fd_sc_hd__o22a_4
X_14329_ _14322_/A _14327_/X _14328_/X VGND VGND VPWR VPWR _14329_/X sky130_fd_sc_hd__and3_4
X_18097_ _18097_/A _18174_/D _18093_/Y VGND VGND VPWR VPWR _18097_/X sky130_fd_sc_hd__and3_4
XANTENNA__12074__A _11993_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21387__A _21373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17048_ _17007_/X _17046_/B VGND VGND VPWR VPWR _17049_/B sky130_fd_sc_hd__and2_4
XANTENNA__12802__A _12802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21975__B1 _23517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21689__A2_N _21688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18999_ _18999_/A VGND VGND VPWR VPWR _18999_/X sky130_fd_sc_hd__buf_2
XFILLER_26_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12521__B _12640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20961_ _20849_/B _20400_/B VGND VGND VPWR VPWR _20961_/X sky130_fd_sc_hd__or2_4
XANTENNA__23886__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15832__B _15902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22700_ _22671_/A VGND VGND VPWR VPWR _22700_/X sky130_fd_sc_hd__buf_2
XFILLER_54_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23680_ _23073_/CLK _23680_/D VGND VGND VPWR VPWR _14912_/B sky130_fd_sc_hd__dfxtp_4
X_20892_ _20892_/A VGND VGND VPWR VPWR _21282_/A sky130_fd_sc_hd__buf_2
XFILLER_0_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20950__A1 _20493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22631_ _22406_/X _22629_/X _16131_/B _22626_/X VGND VGND VPWR VPWR _23127_/D sky130_fd_sc_hd__o22a_4
XFILLER_94_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12249__A _12695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23116__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22562_ _22460_/X _22557_/X _14863_/B _22518_/X VGND VGND VPWR VPWR _23168_/D sky130_fd_sc_hd__o22a_4
XFILLER_22_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24301_ _24301_/CLK _19174_/X HRESETn VGND VGND VPWR VPWR _19122_/A sky130_fd_sc_hd__dfrtp_4
X_21513_ _21512_/X _21508_/X _23771_/Q _21503_/X VGND VGND VPWR VPWR _23771_/D sky130_fd_sc_hd__o22a_4
X_22493_ _22486_/A VGND VGND VPWR VPWR _22493_/X sky130_fd_sc_hd__buf_2
X_24232_ _24203_/CLK _19345_/X HRESETn VGND VGND VPWR VPWR _20792_/A sky130_fd_sc_hd__dfrtp_4
X_21444_ _21289_/X _21440_/X _23809_/Q _21401_/X VGND VGND VPWR VPWR _23809_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22455__B2 _22447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24163_ _24162_/CLK _19870_/X HRESETn VGND VGND VPWR VPWR _11584_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_119_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21375_ _21256_/X _21369_/X _23855_/Q _21373_/X VGND VGND VPWR VPWR _23855_/D sky130_fd_sc_hd__o22a_4
X_23114_ _23561_/CLK _22649_/X VGND VGND VPWR VPWR _13966_/B sky130_fd_sc_hd__dfxtp_4
X_20326_ _20325_/X VGND VGND VPWR VPWR _20497_/A sky130_fd_sc_hd__buf_2
XFILLER_107_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24094_ _23485_/CLK _24094_/D VGND VGND VPWR VPWR _24094_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23045_ _22898_/A _23045_/B VGND VGND VPWR VPWR HADDR[28] sky130_fd_sc_hd__nor2_4
XFILLER_81_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13808__A _13620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15295__A _12531_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20257_ _18761_/X _20257_/B VGND VGND VPWR VPWR _20471_/A sky130_fd_sc_hd__or2_4
XFILLER_115_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12712__A _12198_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20188_ _24094_/Q VGND VGND VPWR VPWR _20188_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12431__B _12430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11961_ _16150_/A VGND VGND VPWR VPWR _16139_/A sky130_fd_sc_hd__buf_2
XANTENNA__23017__A _18162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23947_ _23915_/CLK _23947_/D VGND VGND VPWR VPWR _23947_/Q sky130_fd_sc_hd__dfxtp_4
X_13700_ _13700_/A VGND VGND VPWR VPWR _13765_/A sky130_fd_sc_hd__buf_2
X_14680_ _14666_/X _14680_/B VGND VGND VPWR VPWR _14681_/C sky130_fd_sc_hd__or2_4
XFILLER_79_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11892_ _15041_/A VGND VGND VPWR VPWR _15023_/A sky130_fd_sc_hd__buf_2
X_23878_ _23494_/CLK _23878_/D VGND VGND VPWR VPWR _14301_/B sky130_fd_sc_hd__dfxtp_4
X_13631_ _13631_/A _13631_/B _13631_/C VGND VGND VPWR VPWR _13638_/B sky130_fd_sc_hd__and3_4
X_22829_ _17477_/Y _22825_/X _22862_/A _22828_/X VGND VGND VPWR VPWR _22830_/A sky130_fd_sc_hd__a211o_4
XFILLER_73_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12159__A _11803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13562_ _13562_/A _23855_/Q VGND VGND VPWR VPWR _13563_/C sky130_fd_sc_hd__or2_4
X_16350_ _16364_/A _16282_/B VGND VGND VPWR VPWR _16350_/X sky130_fd_sc_hd__or2_4
XANTENNA__21497__A2 _21470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22694__B2 _22690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20376__A _20212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12513_ _13032_/A _12623_/B VGND VGND VPWR VPWR _12514_/C sky130_fd_sc_hd__or2_4
X_15301_ _14737_/A _15299_/X _15300_/X VGND VGND VPWR VPWR _15302_/C sky130_fd_sc_hd__and3_4
X_16281_ _15936_/A _16279_/X _16280_/X VGND VGND VPWR VPWR _16281_/X sky130_fd_sc_hd__and3_4
X_13493_ _11842_/X _11618_/X _13461_/X _11596_/X _13492_/X VGND VGND VPWR VPWR _13493_/X
+ sky130_fd_sc_hd__a32o_4
X_18020_ _18019_/X VGND VGND VPWR VPWR _18020_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12444_ _12444_/A _12571_/B VGND VGND VPWR VPWR _12444_/X sky130_fd_sc_hd__or2_4
X_15232_ _14243_/A _15224_/X _15231_/X VGND VGND VPWR VPWR _15232_/X sky130_fd_sc_hd__and3_4
XFILLER_51_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14093__B _24009_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15163_ _14096_/X _23809_/Q VGND VGND VPWR VPWR _15163_/X sky130_fd_sc_hd__or2_4
XFILLER_60_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_HCLK_A clkbuf_2_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12375_ _12419_/A _12276_/B VGND VGND VPWR VPWR _12376_/C sky130_fd_sc_hd__or2_4
XANTENNA__23759__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14114_ _15011_/A VGND VGND VPWR VPWR _14165_/A sky130_fd_sc_hd__buf_2
XFILLER_4_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15094_ _12341_/A _23103_/Q VGND VGND VPWR VPWR _15096_/B sky130_fd_sc_hd__or2_4
X_19971_ _19971_/A VGND VGND VPWR VPWR _19971_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14045_ _14045_/A _24042_/Q VGND VGND VPWR VPWR _14046_/C sky130_fd_sc_hd__or2_4
X_18922_ _11533_/D VGND VGND VPWR VPWR _18927_/A sky130_fd_sc_hd__inv_2
XFILLER_69_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18853_ _13918_/X _18848_/X _24391_/Q _18849_/X VGND VGND VPWR VPWR _24391_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21935__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21421__A2 _21419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17804_ _17804_/A VGND VGND VPWR VPWR _17804_/X sky130_fd_sc_hd__buf_2
XFILLER_94_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15933__A _15939_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18784_ _12990_/X _18781_/X _20520_/A _18782_/X VGND VGND VPWR VPWR _18784_/X sky130_fd_sc_hd__o22a_4
X_15996_ _15959_/A _23096_/Q VGND VGND VPWR VPWR _15998_/B sky130_fd_sc_hd__or2_4
X_17735_ _17735_/A _17117_/X VGND VGND VPWR VPWR _17735_/X sky130_fd_sc_hd__and2_4
XANTENNA__15652__B _15652_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14947_ _14937_/A _14873_/B VGND VGND VPWR VPWR _14947_/X sky130_fd_sc_hd__or2_4
XANTENNA__23139__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21185__B2 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13453__A _12462_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17666_ _16947_/Y VGND VGND VPWR VPWR _17667_/A sky130_fd_sc_hd__buf_2
X_14878_ _14995_/A _14874_/X _14878_/C VGND VGND VPWR VPWR _14878_/X sky130_fd_sc_hd__or3_4
XANTENNA__14268__B _14268_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19405_ _19403_/X _18613_/X _19403_/X _24197_/Q VGND VGND VPWR VPWR _24197_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16617_ _16617_/A _24028_/Q VGND VGND VPWR VPWR _16621_/B sky130_fd_sc_hd__or2_4
XANTENNA__13172__B _23953_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13829_ _13645_/A _13829_/B VGND VGND VPWR VPWR _13830_/C sky130_fd_sc_hd__or2_4
XANTENNA__24365__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17597_ _17387_/X VGND VGND VPWR VPWR _18567_/B sky130_fd_sc_hd__inv_2
XFILLER_56_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19336_ _19336_/A VGND VGND VPWR VPWR _19336_/X sky130_fd_sc_hd__buf_2
X_16548_ _16569_/A _16548_/B _16548_/C VGND VGND VPWR VPWR _16554_/B sky130_fd_sc_hd__and3_4
XFILLER_17_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22685__B2 _22683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_21_0_HCLK clkbuf_6_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19267_ _19220_/B VGND VGND VPWR VPWR _19267_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16479_ _16355_/X _16475_/X _16479_/C VGND VGND VPWR VPWR _16479_/X sky130_fd_sc_hd__or3_4
XANTENNA__14284__A _15533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18218_ _18155_/X VGND VGND VPWR VPWR _18218_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19198_ _19110_/A _19110_/B _19197_/Y VGND VGND VPWR VPWR _24289_/D sky130_fd_sc_hd__o21a_4
XFILLER_117_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18149_ _18274_/C _17591_/X _17589_/X VGND VGND VPWR VPWR _18217_/B sky130_fd_sc_hd__o21a_4
X_21160_ _21002_/X _21133_/A _15079_/B _21115_/X VGND VGND VPWR VPWR _21160_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21660__A2 _21655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22006__A _21985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20111_ _11538_/A VGND VGND VPWR VPWR _20111_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13628__A _12509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21091_ _20671_/X _21089_/X _15855_/B _21086_/X VGND VGND VPWR VPWR _21091_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12532__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16004__A _15929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20042_ _19994_/A VGND VGND VPWR VPWR _20042_/X sky130_fd_sc_hd__buf_2
XFILLER_8_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23801_ _23770_/CLK _23801_/D VGND VGND VPWR VPWR _16294_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15562__B _23371_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21993_ _21823_/X _21988_/X _23504_/Q _21992_/X VGND VGND VPWR VPWR _21993_/X sky130_fd_sc_hd__o22a_4
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14459__A _12459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22373__B1 _14279_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23732_ _24021_/CLK _23732_/D VGND VGND VPWR VPWR _12768_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24064__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20944_ _20943_/Y _20851_/X _20939_/B _20675_/X VGND VGND VPWR VPWR _20944_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22676__A _22668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_103_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR _23706_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _23983_/CLK _23663_/D VGND VGND VPWR VPWR _13530_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20875_ _20875_/A _20317_/B VGND VGND VPWR VPWR _20875_/X sky130_fd_sc_hd__or2_4
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16674__A _16652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22614_ _11810_/B VGND VGND VPWR VPWR _22614_/Y sky130_fd_sc_hd__inv_2
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21479__A2 _21477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23594_ _23819_/CLK _23594_/D VGND VGND VPWR VPWR _23594_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20196__A _20196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22545_ _22430_/X _22543_/X _15852_/B _22540_/X VGND VGND VPWR VPWR _23181_/D sky130_fd_sc_hd__o22a_4
XFILLER_22_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19985__A _19985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18601__A2_N _18600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12707__A _12235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22476_ _22476_/A VGND VGND VPWR VPWR _22476_/X sky130_fd_sc_hd__buf_2
X_24215_ _24239_/CLK _19375_/X HRESETn VGND VGND VPWR VPWR _24215_/Q sky130_fd_sc_hd__dfrtp_4
X_21427_ _21258_/X _21426_/X _15690_/B _21423_/X VGND VGND VPWR VPWR _21427_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14922__A _15063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16840__C _16840_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12160_ _11717_/X _23837_/Q VGND VGND VPWR VPWR _12160_/X sky130_fd_sc_hd__or2_4
X_24146_ _24250_/CLK _24146_/D HRESETn VGND VGND VPWR VPWR _24146_/Q sky130_fd_sc_hd__dfrtp_4
X_21358_ _21227_/X _21355_/X _23867_/Q _21352_/X VGND VGND VPWR VPWR _21358_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21651__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20309_ _20308_/X VGND VGND VPWR VPWR _20309_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13538__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12091_ _12091_/A _23837_/Q VGND VGND VPWR VPWR _12092_/C sky130_fd_sc_hd__or2_4
X_24077_ _23922_/CLK _20672_/X VGND VGND VPWR VPWR _15829_/B sky130_fd_sc_hd__dfxtp_4
X_21289_ _21574_/A VGND VGND VPWR VPWR _21289_/X sky130_fd_sc_hd__buf_2
XANTENNA__12442__A _12850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23028_ _18087_/X _23017_/B VGND VGND VPWR VPWR _23029_/C sky130_fd_sc_hd__or2_4
XANTENNA__21755__A _21755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15753__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15850_ _13522_/A _15848_/X _15849_/X VGND VGND VPWR VPWR _15851_/C sky130_fd_sc_hd__and3_4
XFILLER_49_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18280__A1 _18216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16568__B _24060_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14801_ _11669_/A _14793_/X _14800_/X VGND VGND VPWR VPWR _14818_/B sky130_fd_sc_hd__and3_4
XFILLER_79_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15781_ _15778_/X VGND VGND VPWR VPWR _15782_/B sky130_fd_sc_hd__inv_2
X_12993_ _12924_/X _12991_/Y VGND VGND VPWR VPWR _12993_/X sky130_fd_sc_hd__or2_4
XFILLER_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21167__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22364__B1 _15403_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17520_ _18307_/A _17518_/X _17519_/Y VGND VGND VPWR VPWR _17520_/X sky130_fd_sc_hd__o21a_4
X_14732_ _14158_/A _14794_/B VGND VGND VPWR VPWR _14734_/B sky130_fd_sc_hd__or2_4
X_11944_ _11901_/X VGND VGND VPWR VPWR _11994_/A sky130_fd_sc_hd__buf_2
XANTENNA__22586__A _22586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17451_ _12752_/Y _17014_/A _17014_/A _17664_/B VGND VGND VPWR VPWR _17525_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23431__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11875_ _16143_/A VGND VGND VPWR VPWR _11875_/X sky130_fd_sc_hd__buf_2
X_14663_ _15107_/A _14661_/X _14663_/C VGND VGND VPWR VPWR _14663_/X sky130_fd_sc_hd__and3_4
XFILLER_92_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16594__A1 _11992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16584__A _16569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16402_ _16087_/X _16400_/X _16401_/X VGND VGND VPWR VPWR _16403_/C sky130_fd_sc_hd__and3_4
XFILLER_60_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13614_ _13614_/A _13702_/B VGND VGND VPWR VPWR _13614_/X sky130_fd_sc_hd__or2_4
X_17382_ _17382_/A _17382_/B _18405_/A _18428_/A VGND VGND VPWR VPWR _17382_/X sky130_fd_sc_hd__or4_4
X_14594_ _15037_/A VGND VGND VPWR VPWR _14763_/A sky130_fd_sc_hd__buf_2
X_19121_ _19121_/A _19177_/A VGND VGND VPWR VPWR _19122_/B sky130_fd_sc_hd__and2_4
XFILLER_41_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16333_ _16303_/X _16331_/X _16332_/X VGND VGND VPWR VPWR _16333_/X sky130_fd_sc_hd__and3_4
XFILLER_92_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19532__B2 _19531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13545_ _13507_/X _13541_/X _13545_/C VGND VGND VPWR VPWR _13545_/X sky130_fd_sc_hd__or3_4
XFILLER_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23581__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19052_ _18994_/A VGND VGND VPWR VPWR _19052_/X sky130_fd_sc_hd__buf_2
XFILLER_51_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13476_ _13448_/X _23471_/Q VGND VGND VPWR VPWR _13479_/B sky130_fd_sc_hd__or2_4
X_16264_ _11959_/X _23577_/Q VGND VGND VPWR VPWR _16264_/X sky130_fd_sc_hd__or2_4
XANTENNA__22419__B2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21890__A2 _21887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18003_ _18003_/A _18002_/X VGND VGND VPWR VPWR _18003_/X sky130_fd_sc_hd__and2_4
XFILLER_103_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12427_ _13572_/A _12417_/X _12427_/C VGND VGND VPWR VPWR _12428_/C sky130_fd_sc_hd__and3_4
X_15215_ _14190_/A _15211_/X _15215_/C VGND VGND VPWR VPWR _15216_/C sky130_fd_sc_hd__or3_4
X_16195_ _16219_/A _22307_/A VGND VGND VPWR VPWR _16195_/X sky130_fd_sc_hd__or2_4
XANTENNA__18304__A _18425_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12358_ _12421_/A VGND VGND VPWR VPWR _13243_/A sky130_fd_sc_hd__buf_2
X_15146_ _15146_/A _15146_/B VGND VGND VPWR VPWR _15146_/X sky130_fd_sc_hd__or2_4
XANTENNA__21642__A2 _21641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18126__A1_N _17762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13448__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15077_ _15115_/A _15077_/B _15076_/X VGND VGND VPWR VPWR _15077_/X sky130_fd_sc_hd__or3_4
X_19954_ _16935_/X _19364_/X _17006_/X _19953_/X VGND VGND VPWR VPWR _19954_/X sky130_fd_sc_hd__o22a_4
XFILLER_4_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12289_ _12725_/A _12289_/B VGND VGND VPWR VPWR _12289_/X sky130_fd_sc_hd__or2_4
X_14028_ _14046_/A _14025_/X _14027_/X VGND VGND VPWR VPWR _14028_/X sky130_fd_sc_hd__and3_4
X_18905_ _18898_/A VGND VGND VPWR VPWR _18905_/X sky130_fd_sc_hd__buf_2
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19885_ _24159_/Q VGND VGND VPWR VPWR _19885_/Y sky130_fd_sc_hd__inv_2
X_18836_ _17181_/X _18834_/X _24404_/Q _18835_/X VGND VGND VPWR VPWR _24404_/D sky130_fd_sc_hd__o22a_4
XFILLER_95_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15663__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15382__B _15381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18767_ _18789_/A VGND VGND VPWR VPWR _18782_/A sky130_fd_sc_hd__buf_2
X_15979_ _15994_/A _15977_/X _15978_/X VGND VGND VPWR VPWR _15980_/C sky130_fd_sc_hd__and3_4
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21158__B2 _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13183__A _12737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17718_ _18558_/A _17287_/X VGND VGND VPWR VPWR _17718_/X sky130_fd_sc_hd__or2_4
XFILLER_110_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18698_ _17326_/X _18696_/X _18486_/X _18697_/X VGND VGND VPWR VPWR _18698_/X sky130_fd_sc_hd__a211o_4
XFILLER_82_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19789__B _19789_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17649_ _17765_/A _17648_/A VGND VGND VPWR VPWR _17651_/A sky130_fd_sc_hd__or2_4
XANTENNA__24436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20660_ _20468_/X _20659_/Y _19218_/A _20562_/X VGND VGND VPWR VPWR _20660_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22658__B2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19319_ _19318_/X _18005_/X _19318_/X _24250_/Q VGND VGND VPWR VPWR _24250_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13630__B _13630_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20591_ _20591_/A VGND VGND VPWR VPWR _20591_/X sky130_fd_sc_hd__buf_2
XANTENNA__12527__A _12466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22330_ _14875_/B VGND VGND VPWR VPWR _22330_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22261_ _22081_/X _22258_/X _16749_/B _22255_/X VGND VGND VPWR VPWR _22261_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15838__A _12915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18214__A _17871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14742__A _15413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24000_ _24065_/CLK _24000_/D VGND VGND VPWR VPWR _14866_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_3_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21212_ _21212_/A _21212_/B VGND VGND VPWR VPWR _21213_/A sky130_fd_sc_hd__or2_4
XANTENNA__21094__B1 _24011_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22192_ _22134_/X _22186_/X _14473_/B _22190_/X VGND VGND VPWR VPWR _22192_/X sky130_fd_sc_hd__o22a_4
X_21143_ _20697_/X _21140_/X _15407_/B _21137_/X VGND VGND VPWR VPWR _21143_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_28_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR _24180_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12262__A _12743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15312__A2 _13595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23304__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21074_ _20394_/X _21068_/X _24025_/Q _21072_/X VGND VGND VPWR VPWR _21074_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20025_ _20025_/A VGND VGND VPWR VPWR _20025_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21149__A1 _20797_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21149__B2 _21144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18884__A _18891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22346__B1 _16253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22897__A1 _22886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21976_ _21795_/X _21974_/X _23516_/Q _21971_/X VGND VGND VPWR VPWR _23516_/D sky130_fd_sc_hd__o22a_4
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20927_ _20403_/A _20926_/X _24258_/Q _20736_/X VGND VGND VPWR VPWR _20927_/X sky130_fd_sc_hd__o22a_4
X_23715_ _23363_/CLK _23715_/D VGND VGND VPWR VPWR _14791_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13821__A _15432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11651_/A VGND VGND VPWR VPWR _11661_/A sky130_fd_sc_hd__buf_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _20858_/A VGND VGND VPWR VPWR _20858_/Y sky130_fd_sc_hd__inv_2
X_23646_ _23774_/CLK _21739_/X VGND VGND VPWR VPWR _23646_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22649__B2 _22647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24106__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _17083_/A _11579_/X _11591_/C _11591_/D VGND VGND VPWR VPWR _11622_/A sky130_fd_sc_hd__or4_4
X_23577_ _23514_/CLK _23577_/D VGND VGND VPWR VPWR _23577_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_70_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20789_ _20732_/X _20788_/X _24296_/Q _20739_/X VGND VGND VPWR VPWR _20790_/B sky130_fd_sc_hd__o22a_4
XFILLER_10_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21321__B2 _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _13303_/X _13328_/X _13329_/X VGND VGND VPWR VPWR _13330_/X sky130_fd_sc_hd__and3_4
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22528_ _22401_/X _22522_/X _16248_/B _22526_/X VGND VGND VPWR VPWR _23193_/D sky130_fd_sc_hd__o22a_4
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13242_/A _24081_/Q VGND VGND VPWR VPWR _13262_/C sky130_fd_sc_hd__or2_4
XFILLER_104_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15748__A _13130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22459_ _22458_/X _22452_/X _15125_/B _22386_/X VGND VGND VPWR VPWR _22459_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14652__A _14679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12212_ _12211_/X VGND VGND VPWR VPWR _13046_/A sky130_fd_sc_hd__buf_2
X_15000_ _14151_/A _23263_/Q VGND VGND VPWR VPWR _15000_/X sky130_fd_sc_hd__or2_4
XANTENNA__21085__B1 _24017_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13192_ _15820_/A _13187_/X _13191_/X VGND VGND VPWR VPWR _13192_/X sky130_fd_sc_hd__or3_4
XANTENNA__21624__A2 _21619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12143_ _12167_/A _23677_/Q VGND VGND VPWR VPWR _12145_/B sky130_fd_sc_hd__or2_4
X_24129_ _23522_/CLK _20013_/Y HRESETn VGND VGND VPWR VPWR _24129_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13268__A _12392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12074_ _11993_/A _23933_/Q VGND VGND VPWR VPWR _12074_/X sky130_fd_sc_hd__or2_4
X_16951_ _16951_/A VGND VGND VPWR VPWR _17680_/A sky130_fd_sc_hd__inv_2
XFILLER_81_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21388__A1 _21277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21388__B2 _21387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22585__B1 _23156_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15902_ _13562_/A _15902_/B VGND VGND VPWR VPWR _15903_/C sky130_fd_sc_hd__or2_4
X_19670_ _19485_/A VGND VGND VPWR VPWR _19670_/X sky130_fd_sc_hd__buf_2
XFILLER_46_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16882_ _16081_/X _16881_/X _16081_/X _16881_/X VGND VGND VPWR VPWR _16887_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12900__A _12528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18621_ _18137_/A _18621_/B VGND VGND VPWR VPWR _18621_/X sky130_fd_sc_hd__and2_4
X_15833_ _12493_/A _15831_/X _15832_/X VGND VGND VPWR VPWR _15834_/C sky130_fd_sc_hd__and3_4
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14099__A _14136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18552_ _18480_/X _18549_/X _18508_/X _18551_/X VGND VGND VPWR VPWR _18552_/X sky130_fd_sc_hd__o22a_4
X_15764_ _12777_/X _15762_/X _15763_/X VGND VGND VPWR VPWR _15768_/B sky130_fd_sc_hd__and3_4
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12976_ _12976_/A _12976_/B VGND VGND VPWR VPWR _12978_/B sky130_fd_sc_hd__or2_4
XFILLER_94_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17503_ _17502_/X VGND VGND VPWR VPWR _18281_/A sky130_fd_sc_hd__inv_2
XANTENNA__19753__A1 _20939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14715_ _15623_/A _14715_/B _14715_/C VGND VGND VPWR VPWR _14716_/C sky130_fd_sc_hd__and3_4
XFILLER_94_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11927_ _12301_/A VGND VGND VPWR VPWR _14752_/A sky130_fd_sc_hd__buf_2
X_18483_ _18097_/A _18350_/B _18481_/Y _18016_/A _22944_/B VGND VGND VPWR VPWR _18484_/A
+ sky130_fd_sc_hd__a32o_4
X_15695_ _15695_/A _15695_/B _15694_/X VGND VGND VPWR VPWR _15695_/X sky130_fd_sc_hd__or3_4
X_17434_ _15911_/X _17377_/B VGND VGND VPWR VPWR _17434_/Y sky130_fd_sc_hd__nand2_4
X_14646_ _11710_/A _14646_/B VGND VGND VPWR VPWR _14647_/C sky130_fd_sc_hd__or2_4
XFILLER_61_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11858_ _15449_/A VGND VGND VPWR VPWR _11859_/A sky130_fd_sc_hd__buf_2
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17365_ _17365_/A VGND VGND VPWR VPWR _17365_/X sky130_fd_sc_hd__buf_2
X_11789_ _11729_/X VGND VGND VPWR VPWR _11823_/A sky130_fd_sc_hd__buf_2
X_14577_ _15144_/A _14574_/X _14577_/C VGND VGND VPWR VPWR _14577_/X sky130_fd_sc_hd__and3_4
XFILLER_60_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12347__A _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19104_ _24319_/Q VGND VGND VPWR VPWR _19104_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16316_ _16366_/A _16316_/B _16316_/C VGND VGND VPWR VPWR _16316_/X sky130_fd_sc_hd__and3_4
X_13528_ _13507_/X _13528_/B _13528_/C VGND VGND VPWR VPWR _13528_/X sky130_fd_sc_hd__or3_4
X_17296_ _17605_/A _17295_/X VGND VGND VPWR VPWR _17336_/B sky130_fd_sc_hd__and2_4
XFILLER_70_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19035_ _19024_/X _19033_/X _19034_/Y _19027_/X VGND VGND VPWR VPWR _19035_/X sky130_fd_sc_hd__o22a_4
X_16247_ _16152_/A _16242_/X _16246_/X VGND VGND VPWR VPWR _16247_/X sky130_fd_sc_hd__or3_4
XANTENNA__15658__A _12556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13459_ _12528_/A _13455_/X _13459_/C VGND VGND VPWR VPWR _13460_/B sky130_fd_sc_hd__or3_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14562__A _11799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21615__A2 _21612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16178_ _16206_/A _16178_/B _16177_/X VGND VGND VPWR VPWR _16179_/C sky130_fd_sc_hd__and3_4
XANTENNA__13178__A _12728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15129_ _14089_/A _23713_/Q VGND VGND VPWR VPWR _15129_/X sky130_fd_sc_hd__or2_4
XFILLER_64_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19937_ _19936_/X VGND VGND VPWR VPWR _20176_/A sky130_fd_sc_hd__inv_2
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21379__B2 _21373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15393__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13906__A _13910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19868_ _19740_/A _19822_/A VGND VGND VPWR VPWR _19868_/X sky130_fd_sc_hd__and2_4
XFILLER_110_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22040__A2 _22038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18819_ _18841_/A VGND VGND VPWR VPWR _18842_/A sky130_fd_sc_hd__inv_2
X_19799_ _19798_/X VGND VGND VPWR VPWR _19799_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21830_ _21828_/X _21829_/X _15685_/B _21824_/X VGND VGND VPWR VPWR _23598_/D sky130_fd_sc_hd__o22a_4
XFILLER_83_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21761_ _21541_/X _21755_/X _13569_/B _21759_/X VGND VGND VPWR VPWR _23631_/D sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_4_3_0_HCLK_A clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14737__A _14737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20712_ _20704_/X _20711_/Y _19216_/A _20562_/X VGND VGND VPWR VPWR _20712_/X sky130_fd_sc_hd__o22a_4
X_23500_ _23692_/CLK _23500_/D VGND VGND VPWR VPWR _15455_/B sky130_fd_sc_hd__dfxtp_4
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13641__A _13641_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21692_ _21506_/X _21691_/X _23677_/Q _21688_/X VGND VGND VPWR VPWR _21692_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23431_ _23079_/CLK _23431_/D VGND VGND VPWR VPWR _13875_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20643_ _17068_/A VGND VGND VPWR VPWR _22855_/A sky130_fd_sc_hd__buf_2
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12257__A _12257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21303__B2 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23362_ _24066_/CLK _23362_/D VGND VGND VPWR VPWR _15292_/B sky130_fd_sc_hd__dfxtp_4
X_20574_ _20574_/A VGND VGND VPWR VPWR _20574_/X sky130_fd_sc_hd__buf_2
XFILLER_20_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21854__A2 _21853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22313_ _13157_/B VGND VGND VPWR VPWR _22313_/X sky130_fd_sc_hd__buf_2
X_23293_ _23293_/CLK _23293_/D VGND VGND VPWR VPWR _12132_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14472__A _13019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22244_ _22136_/X _22243_/X _14698_/B _22240_/X VGND VGND VPWR VPWR _22244_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21606__A2 _21605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17783__A _17782_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22175_ _22105_/X _22172_/X _13249_/B _22169_/X VGND VGND VPWR VPWR _23409_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21126_ _21133_/A VGND VGND VPWR VPWR _21126_/X sky130_fd_sc_hd__buf_2
X_21057_ _21002_/X _21030_/A _15023_/B _21012_/X VGND VGND VPWR VPWR _24031_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12720__A _12720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20008_ _20007_/X VGND VGND VPWR VPWR _20008_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21790__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12830_ _12830_/A _12830_/B _12830_/C VGND VGND VPWR VPWR _12830_/X sky130_fd_sc_hd__and3_4
XFILLER_55_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15750__B _15685_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12761_ _13130_/A VGND VGND VPWR VPWR _12816_/A sky130_fd_sc_hd__buf_2
XFILLER_76_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _21919_/A VGND VGND VPWR VPWR _21959_/X sky130_fd_sc_hd__buf_2
XANTENNA__14647__A _15114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18119__A _17874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21542__B2 _21539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _13887_/A VGND VGND VPWR VPWR _14500_/X sky130_fd_sc_hd__buf_2
XANTENNA__13551__A _12980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11712_ _13257_/A VGND VGND VPWR VPWR _12381_/A sky130_fd_sc_hd__buf_2
XFILLER_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12688_/A _12692_/B _12692_/C VGND VGND VPWR VPWR _12696_/B sky130_fd_sc_hd__and3_4
X_15480_ _15480_/A _23308_/Q VGND VGND VPWR VPWR _15482_/B sky130_fd_sc_hd__or2_4
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _15114_/A VGND VGND VPWR VPWR _12421_/A sky130_fd_sc_hd__buf_2
X_14431_ _14431_/A _14431_/B VGND VGND VPWR VPWR _14433_/B sky130_fd_sc_hd__or2_4
XFILLER_93_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ _23922_/CLK _21764_/X VGND VGND VPWR VPWR _15902_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17958__A _18066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _17150_/A VGND VGND VPWR VPWR _17251_/A sky130_fd_sc_hd__buf_2
XFILLER_50_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11574_ _20086_/A _20098_/B _20090_/B _20090_/A VGND VGND VPWR VPWR _20071_/A sky130_fd_sc_hd__or4_4
X_14362_ _14379_/A _14279_/B VGND VGND VPWR VPWR _14362_/X sky130_fd_sc_hd__or2_4
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16101_ _16100_/X VGND VGND VPWR VPWR _16146_/A sky130_fd_sc_hd__buf_2
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18710__A2 _16997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _12740_/A _13311_/X _13312_/X VGND VGND VPWR VPWR _13313_/X sky130_fd_sc_hd__and3_4
XFILLER_7_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15478__A _12585_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14293_ _15447_/A _14293_/B VGND VGND VPWR VPWR _14294_/C sky130_fd_sc_hd__or2_4
X_17081_ _17081_/A _17900_/A VGND VGND VPWR VPWR _17081_/X sky130_fd_sc_hd__and2_4
XFILLER_52_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13244_ _12367_/A _13240_/X _13244_/C VGND VGND VPWR VPWR _13252_/B sky130_fd_sc_hd__or3_4
X_16032_ _16048_/A _16032_/B _16032_/C VGND VGND VPWR VPWR _16036_/B sky130_fd_sc_hd__and3_4
XFILLER_87_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_14_0_HCLK_A clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13175_ _12730_/A _24049_/Q VGND VGND VPWR VPWR _13176_/C sky130_fd_sc_hd__or2_4
XFILLER_48_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22270__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12126_ _11773_/X _12123_/X _12126_/C VGND VGND VPWR VPWR _12127_/C sky130_fd_sc_hd__and3_4
X_17983_ _17926_/X _17981_/Y _17812_/X _17982_/Y VGND VGND VPWR VPWR _17983_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_7_11_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR _23907_/CLK sky130_fd_sc_hd__clkbuf_1
X_19722_ _19722_/A _19689_/A VGND VGND VPWR VPWR _19723_/B sky130_fd_sc_hd__or2_4
XFILLER_42_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_74_0_HCLK clkbuf_7_75_0_HCLK/A VGND VGND VPWR VPWR _23840_/CLK sky130_fd_sc_hd__clkbuf_1
X_12057_ _12086_/A _24029_/Q VGND VGND VPWR VPWR _12060_/B sky130_fd_sc_hd__or2_4
X_16934_ _18171_/A VGND VGND VPWR VPWR _16935_/A sky130_fd_sc_hd__buf_2
XANTENNA__13726__A _13726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12630__A _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19653_ _19486_/Y VGND VGND VPWR VPWR _19667_/A sky130_fd_sc_hd__buf_2
X_16865_ _16858_/X _16859_/X _16865_/C _16865_/D VGND VGND VPWR VPWR _16865_/X sky130_fd_sc_hd__or4_4
XFILLER_4_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18604_ _18603_/Y VGND VGND VPWR VPWR _18604_/X sky130_fd_sc_hd__buf_2
XANTENNA__21781__B2 _21737_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15816_ _12859_/A _15814_/X _15815_/X VGND VGND VPWR VPWR _15816_/X sky130_fd_sc_hd__and3_4
XFILLER_24_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19584_ _19537_/A _19579_/X _19581_/X _19583_/X VGND VGND VPWR VPWR _19584_/X sky130_fd_sc_hd__a211o_4
X_16796_ _16803_/A _23099_/Q VGND VGND VPWR VPWR _16796_/X sky130_fd_sc_hd__or2_4
XFILLER_34_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18535_ _18097_/A _18348_/B _18533_/Y _18016_/A _22932_/B VGND VGND VPWR VPWR _18536_/A
+ sky130_fd_sc_hd__a32o_4
X_15747_ _13129_/A _15747_/B VGND VGND VPWR VPWR _15749_/B sky130_fd_sc_hd__or2_4
XFILLER_59_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15660__B _15722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12959_ _12959_/A _23955_/Q VGND VGND VPWR VPWR _12960_/C sky130_fd_sc_hd__or2_4
XFILLER_94_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21533__A1 _21531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18029__A _18421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14557__A _11648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21533__B2 _21527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18466_ _18101_/A _18466_/B VGND VGND VPWR VPWR _18468_/C sky130_fd_sc_hd__nor2_4
X_15678_ _12744_/A _15678_/B _15678_/C VGND VGND VPWR VPWR _15678_/X sky130_fd_sc_hd__and3_4
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14276__B _14276_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17417_ _17414_/X VGND VGND VPWR VPWR _17427_/B sky130_fd_sc_hd__inv_2
X_14629_ _13603_/A _14629_/B _14628_/X VGND VGND VPWR VPWR _14630_/C sky130_fd_sc_hd__and3_4
X_18397_ _18418_/B _18396_/X VGND VGND VPWR VPWR _18397_/X sky130_fd_sc_hd__or2_4
X_17348_ _15648_/X _17348_/B VGND VGND VPWR VPWR _17349_/A sky130_fd_sc_hd__or2_4
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17279_ _17277_/X _17278_/B VGND VGND VPWR VPWR _17902_/B sky130_fd_sc_hd__or2_4
XANTENNA__16712__A1 _12036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12805__A _12753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19018_ _24335_/Q VGND VGND VPWR VPWR _19018_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21049__B1 _14305_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20290_ _20516_/A VGND VGND VPWR VPWR _20290_/X sky130_fd_sc_hd__buf_2
XFILLER_118_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15835__B _15835_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13636__A _13636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22013__A2 _22009_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23980_ _24044_/CLK _21143_/X VGND VGND VPWR VPWR _15407_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12540__A _12540_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22931_ _22931_/A VGND VGND VPWR VPWR HADDR[8] sky130_fd_sc_hd__inv_2
XFILLER_83_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21772__B2 _21766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15851__A _15889_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22862_ _22862_/A VGND VGND VPWR VPWR _22872_/A sky130_fd_sc_hd__buf_2
XFILLER_83_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15451__A1 _11977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21813_ _21811_/X _21805_/X _12525_/B _21812_/X VGND VGND VPWR VPWR _23605_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15570__B _15570_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22793_ _22779_/X VGND VGND VPWR VPWR _22794_/A sky130_fd_sc_hd__buf_2
XANTENNA__14467__A _12862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13371__A _12787_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21744_ _21512_/X _21741_/X _23643_/Q _21738_/X VGND VGND VPWR VPWR _23643_/D sky130_fd_sc_hd__o22a_4
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21675_ _21565_/X _21669_/X _14486_/B _21673_/X VGND VGND VPWR VPWR _23685_/D sky130_fd_sc_hd__o22a_4
X_24463_ _24126_/CLK _24463_/D HRESETn VGND VGND VPWR VPWR _20029_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21288__B1 _15273_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20626_ _20448_/X _20624_/X _24366_/Q _20625_/X VGND VGND VPWR VPWR _20626_/X sky130_fd_sc_hd__o22a_4
X_23414_ _23155_/CLK _22168_/X VGND VGND VPWR VPWR _12298_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24394_ _24365_/CLK _18850_/X HRESETn VGND VGND VPWR VPWR _24394_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21827__A2 _21817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23345_ _23217_/CLK _23345_/D VGND VGND VPWR VPWR _13140_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20557_ _24401_/Q _20595_/B VGND VGND VPWR VPWR _20557_/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23276_ _24044_/CLK _22364_/X VGND VGND VPWR VPWR _15403_/B sky130_fd_sc_hd__dfxtp_4
X_20488_ _20488_/A VGND VGND VPWR VPWR _20488_/X sky130_fd_sc_hd__buf_2
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22227_ _22107_/X _22222_/X _13328_/B _22226_/X VGND VGND VPWR VPWR _22227_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18456__B2 _18455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23792__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22158_ _22172_/A VGND VGND VPWR VPWR _22158_/X sky130_fd_sc_hd__buf_2
XFILLER_79_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21109_ _21002_/X _21075_/A _23999_/Q _21072_/A VGND VGND VPWR VPWR _23999_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13546__A _12965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22004__A2 _22002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14980_ _14644_/A _14905_/B VGND VGND VPWR VPWR _14980_/X sky130_fd_sc_hd__or2_4
X_22089_ _22101_/A VGND VGND VPWR VPWR _22089_/X sky130_fd_sc_hd__buf_2
XANTENNA__12450__A _12450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13931_ _13960_/A _23722_/Q VGND VGND VPWR VPWR _13932_/C sky130_fd_sc_hd__or2_4
XANTENNA__24148__CLK _24223_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15761__A _13102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21763__B2 _21759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16650_ _16662_/A _23612_/Q VGND VGND VPWR VPWR _16650_/X sky130_fd_sc_hd__or2_4
X_13862_ _13862_/A VGND VGND VPWR VPWR _13879_/A sky130_fd_sc_hd__buf_2
XFILLER_75_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15601_ _15601_/A _23147_/Q VGND VGND VPWR VPWR _15603_/B sky130_fd_sc_hd__or2_4
XANTENNA__24121__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12813_ _12813_/A _12811_/X _12813_/C VGND VGND VPWR VPWR _12814_/C sky130_fd_sc_hd__and3_4
XANTENNA__19708__B2 _19707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16581_ _16715_/A _16581_/B _16581_/C VGND VGND VPWR VPWR _16581_/X sky130_fd_sc_hd__and3_4
XFILLER_90_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13793_ _13624_/A _13793_/B _13792_/X VGND VGND VPWR VPWR _13793_/X sky130_fd_sc_hd__and3_4
X_18320_ _18266_/A _17490_/Y VGND VGND VPWR VPWR _18321_/D sky130_fd_sc_hd__and2_4
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24298__CLK _24299_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23172__CLK _23107_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13281__A _15654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15532_ _14283_/A _24011_/Q VGND VGND VPWR VPWR _15532_/X sky130_fd_sc_hd__or2_4
XFILLER_91_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12744_ _12744_/A _12742_/X _12743_/X VGND VGND VPWR VPWR _12748_/B sky130_fd_sc_hd__and3_4
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18251_ _17874_/A _18250_/X VGND VGND VPWR VPWR _18251_/Y sky130_fd_sc_hd__nor2_4
XFILLER_97_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15463_ _15487_/A _15463_/B VGND VGND VPWR VPWR _15463_/X sky130_fd_sc_hd__or2_4
X_12675_ _12674_/X VGND VGND VPWR VPWR _12675_/Y sky130_fd_sc_hd__inv_2
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16592__A _11924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _17175_/Y _17173_/X _15648_/X _17145_/X VGND VGND VPWR VPWR _17202_/X sky130_fd_sc_hd__o22a_4
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _15617_/A _14317_/B VGND VGND VPWR VPWR _14414_/X sky130_fd_sc_hd__or2_4
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12559__A2 _11618_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21279__B1 _14292_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _11625_/X VGND VGND VPWR VPWR _11626_/Y sky130_fd_sc_hd__inv_2
X_18182_ _17837_/X _17199_/X _17975_/X _17216_/X VGND VGND VPWR VPWR _18182_/X sky130_fd_sc_hd__o22a_4
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21818__A2 _21817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ _12861_/A _15394_/B _15394_/C VGND VGND VPWR VPWR _15394_/X sky130_fd_sc_hd__and3_4
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _17145_/A VGND VGND VPWR VPWR _17133_/X sky130_fd_sc_hd__buf_2
XFILLER_50_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ _14345_/A VGND VGND VPWR VPWR _15616_/A sky130_fd_sc_hd__buf_2
X_11557_ _24426_/Q IRQ[11] _11556_/X VGND VGND VPWR VPWR _11558_/B sky130_fd_sc_hd__a21o_4
XFILLER_89_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22491__A2 _22486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12625__A _12948_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15001__A _15028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17064_ _17145_/A VGND VGND VPWR VPWR _17157_/A sky130_fd_sc_hd__buf_2
XANTENNA__21938__A _21938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14276_ _12260_/X _14276_/B VGND VGND VPWR VPWR _14276_/X sky130_fd_sc_hd__or2_4
XFILLER_100_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16015_ _16025_/A VGND VGND VPWR VPWR _16047_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13227_ _12367_/A _13227_/B _13226_/X VGND VGND VPWR VPWR _13227_/X sky130_fd_sc_hd__or3_4
XFILLER_100_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19644__B1 _19481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13158_ _15707_/A VGND VGND VPWR VPWR _15697_/A sky130_fd_sc_hd__buf_2
XFILLER_83_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12109_ _12008_/A _23709_/Q VGND VGND VPWR VPWR _12111_/B sky130_fd_sc_hd__or2_4
XFILLER_111_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13456__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13089_ _13098_/A _13089_/B VGND VGND VPWR VPWR _13089_/X sky130_fd_sc_hd__or2_4
X_17966_ _17242_/A VGND VGND VPWR VPWR _17966_/X sky130_fd_sc_hd__buf_2
XFILLER_117_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15681__A1 _12682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16917_ _16891_/Y _16917_/B _16917_/C VGND VGND VPWR VPWR _16918_/C sky130_fd_sc_hd__and3_4
X_19705_ _19703_/A _19822_/A _19672_/C _19607_/X VGND VGND VPWR VPWR _19705_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21673__A _21659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17897_ _17896_/X VGND VGND VPWR VPWR _17897_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21754__B2 _21752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15671__A _12705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16848_ _15914_/C VGND VGND VPWR VPWR _16850_/A sky130_fd_sc_hd__inv_2
X_19636_ _19549_/X _19617_/X _19635_/X _17543_/A _19585_/X VGND VGND VPWR VPWR _19636_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_65_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_4_0_HCLK clkbuf_6_2_0_HCLK/X VGND VGND VPWR VPWR _24199_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19567_ _19566_/X VGND VGND VPWR VPWR _19629_/A sky130_fd_sc_hd__buf_2
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16779_ _16624_/X _16779_/B _16779_/C VGND VGND VPWR VPWR _16780_/C sky130_fd_sc_hd__and3_4
XANTENNA__14287__A _15536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13191__A _12849_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18518_ _18517_/X VGND VGND VPWR VPWR _18518_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11704__A _16071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19498_ _20650_/A _19496_/X _19497_/X HRDATA[14] VGND VGND VPWR VPWR _19498_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__19797__B _19796_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12519__B _12639_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23665__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18449_ _18401_/X VGND VGND VPWR VPWR _18449_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21460_ _21452_/X VGND VGND VPWR VPWR _21460_/X sky130_fd_sc_hd__buf_2
XFILLER_18_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22009__A _22002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20411_ _20321_/X _20410_/X _24312_/Q _20330_/X VGND VGND VPWR VPWR _20411_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21391_ _21282_/X _21390_/X _14635_/B _21387_/X VGND VGND VPWR VPWR _23844_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22482__A2 _22479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12535__A _12904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23130_ _23130_/CLK _22627_/X VGND VGND VPWR VPWR _16489_/B sky130_fd_sc_hd__dfxtp_4
X_20342_ _20342_/A _20342_/B VGND VGND VPWR VPWR _20342_/X sky130_fd_sc_hd__and2_4
XANTENNA__21848__A _21812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20752__A _18577_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23061_ _20194_/A _11634_/B _16929_/B _19933_/A VGND VGND VPWR VPWR _23062_/A sky130_fd_sc_hd__or4_4
XANTENNA__18438__A1 _18011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15846__A _12386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20273_ _20213_/X _20230_/X _20233_/X _20272_/Y VGND VGND VPWR VPWR _20273_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22234__A2 _22229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19318__A _19328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14750__A _13960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22012_ _21857_/X _22009_/X _15253_/B _22006_/X VGND VGND VPWR VPWR _23490_/D sky130_fd_sc_hd__o22a_4
XFILLER_118_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21993__A1 _21823_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21993__B2 _21992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12270__A _12235_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22679__A _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21583__A _21583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13085__B _13085_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23963_ _23515_/CLK _23963_/D VGND VGND VPWR VPWR _23963_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16677__A _16677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22914_ _22980_/A VGND VGND VPWR VPWR _23038_/B sky130_fd_sc_hd__buf_2
XFILLER_99_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23894_ _23920_/CLK _21315_/X VGND VGND VPWR VPWR _12285_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22845_ _12752_/Y _22824_/X _22831_/X _22844_/X VGND VGND VPWR VPWR _22846_/A sky130_fd_sc_hd__a211o_4
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18892__A _18892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22776_ _20194_/A _17032_/B _20196_/A VGND VGND VPWR VPWR _22777_/A sky130_fd_sc_hd__or3_4
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18374__B1 _17634_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22170__B2 _22169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21727_ _21567_/X _21726_/X _14679_/B _21723_/X VGND VGND VPWR VPWR _21727_/X sky130_fd_sc_hd__o22a_4
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12460_ _12460_/A VGND VGND VPWR VPWR _12891_/A sky130_fd_sc_hd__buf_2
X_21658_ _21536_/X _21655_/X _13196_/B _21652_/X VGND VGND VPWR VPWR _23697_/D sky130_fd_sc_hd__o22a_4
X_24446_ _24435_/CLK _18769_/X HRESETn VGND VGND VPWR VPWR _24446_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18126__B1 _17762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12391_ _11665_/X _12364_/X _12390_/X VGND VGND VPWR VPWR _12429_/B sky130_fd_sc_hd__or3_4
X_20609_ _24207_/Q _20512_/X _20608_/X VGND VGND VPWR VPWR _20610_/A sky130_fd_sc_hd__o21a_4
X_21589_ _21580_/Y _21588_/X _21504_/X _21588_/X VGND VGND VPWR VPWR _21589_/X sky130_fd_sc_hd__a2bb2o_4
X_24377_ _24435_/CLK _24377_/D HRESETn VGND VGND VPWR VPWR _18961_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__12445__A _15823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22473__A2 _22472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14130_ _11879_/A _23881_/Q VGND VGND VPWR VPWR _14132_/B sky130_fd_sc_hd__or2_4
X_23328_ _23104_/CLK _22298_/X VGND VGND VPWR VPWR _14859_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14061_ _14065_/A _14059_/X _14060_/X VGND VGND VPWR VPWR _14062_/C sky130_fd_sc_hd__and3_4
XANTENNA__22225__A2 _22222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23259_ _23260_/CLK _22397_/X VGND VGND VPWR VPWR _16744_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_3_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18132__A _18174_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13012_ _13031_/A _23666_/Q VGND VGND VPWR VPWR _13012_/X sky130_fd_sc_hd__or2_4
XFILLER_79_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_6_0_HCLK_A clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17820_ _17813_/X _17816_/X _17818_/X _17819_/X VGND VGND VPWR VPWR _17820_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_95_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21984__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17751_ _18459_/A _17346_/X _17703_/X _17750_/X VGND VGND VPWR VPWR _17751_/X sky130_fd_sc_hd__o22a_4
XFILLER_43_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24302__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14963_ _12582_/A _23808_/Q VGND VGND VPWR VPWR _14964_/C sky130_fd_sc_hd__or2_4
XFILLER_43_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16587__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16702_ _12044_/X _16702_/B _16702_/C VGND VGND VPWR VPWR _16703_/C sky130_fd_sc_hd__and3_4
XANTENNA__15491__A _15491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13914_ _12617_/A _13914_/B _13914_/C VGND VGND VPWR VPWR _13915_/C sky130_fd_sc_hd__and3_4
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17682_ _17757_/A _17680_/X _17758_/A VGND VGND VPWR VPWR _18286_/A sky130_fd_sc_hd__a21o_4
X_14894_ _13956_/A _14894_/B _14893_/X VGND VGND VPWR VPWR _14894_/X sky130_fd_sc_hd__or3_4
XFILLER_21_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19421_ _19462_/A VGND VGND VPWR VPWR _19458_/A sky130_fd_sc_hd__inv_2
X_16633_ _16670_/A _16559_/B VGND VGND VPWR VPWR _16634_/C sky130_fd_sc_hd__or2_4
XFILLER_74_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13845_ _13845_/A _23495_/Q VGND VGND VPWR VPWR _13846_/C sky130_fd_sc_hd__or2_4
XFILLER_112_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19898__A _22932_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19352_ _19350_/X _18654_/X _19350_/X _24227_/Q VGND VGND VPWR VPWR _19352_/X sky130_fd_sc_hd__a2bb2o_4
X_16564_ _16538_/A _23900_/Q VGND VGND VPWR VPWR _16566_/B sky130_fd_sc_hd__or2_4
X_13776_ _13776_/A _13775_/Y VGND VGND VPWR VPWR _13776_/X sky130_fd_sc_hd__or2_4
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20837__A _22446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18303_ _18040_/X _17851_/X _17868_/X VGND VGND VPWR VPWR _18304_/B sky130_fd_sc_hd__o21ai_4
XFILLER_108_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22161__B2 _22155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15515_ _11671_/A _15515_/B _15515_/C VGND VGND VPWR VPWR _15515_/X sky130_fd_sc_hd__and3_4
XFILLER_17_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12727_ _15664_/A _12727_/B _12727_/C VGND VGND VPWR VPWR _12732_/B sky130_fd_sc_hd__and3_4
X_19283_ _19212_/B VGND VGND VPWR VPWR _19283_/Y sky130_fd_sc_hd__inv_2
X_16495_ _16355_/X _16491_/X _16495_/C VGND VGND VPWR VPWR _16496_/C sky130_fd_sc_hd__or3_4
X_18234_ _18234_/A _18234_/B VGND VGND VPWR VPWR _18235_/A sky130_fd_sc_hd__and2_4
X_15446_ _12203_/A _15504_/B VGND VGND VPWR VPWR _15448_/B sky130_fd_sc_hd__or2_4
X_12658_ _12643_/A _12658_/B VGND VGND VPWR VPWR _12659_/C sky130_fd_sc_hd__or2_4
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11609_ _14101_/A VGND VGND VPWR VPWR _11610_/A sky130_fd_sc_hd__buf_2
X_18165_ _18285_/C _17760_/X _17684_/X VGND VGND VPWR VPWR _18165_/X sky130_fd_sc_hd__o21a_4
X_15377_ _13991_/A _15369_/X _15377_/C VGND VGND VPWR VPWR _15378_/C sky130_fd_sc_hd__and3_4
X_12589_ _11740_/A VGND VGND VPWR VPWR _13731_/A sky130_fd_sc_hd__buf_2
XANTENNA__12355__A _12826_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17116_ _21583_/A VGND VGND VPWR VPWR _19841_/A sky130_fd_sc_hd__inv_2
X_14328_ _15574_/A _14328_/B VGND VGND VPWR VPWR _14328_/X sky130_fd_sc_hd__or2_4
X_18096_ _16999_/C VGND VGND VPWR VPWR _18174_/D sky130_fd_sc_hd__buf_2
XANTENNA__12074__B _23933_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17047_ _17047_/A VGND VGND VPWR VPWR _17047_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15666__A _15685_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14259_ _11669_/A _14259_/B _14259_/C VGND VGND VPWR VPWR _14260_/C sky130_fd_sc_hd__and3_4
XANTENNA__22216__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24325__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21975__B2 _21971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13186__A _12739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18840__A1 _17194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18998_ _24371_/Q VGND VGND VPWR VPWR _18998_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_44_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_44_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17949_ _17888_/X _17948_/X _19971_/A _17888_/X VGND VGND VPWR VPWR _24475_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21727__B2 _21723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20960_ _20846_/B HRDATA[17] VGND VGND VPWR VPWR _20960_/X sky130_fd_sc_hd__or2_4
XFILLER_54_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19619_ _19424_/A _19618_/X HRDATA[2] _19439_/X VGND VGND VPWR VPWR _19645_/A sky130_fd_sc_hd__o22a_4
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20891_ _24196_/Q _20873_/X _20890_/Y VGND VGND VPWR VPWR _20892_/A sky130_fd_sc_hd__o21a_4
XFILLER_80_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22630_ _22403_/X _22629_/X _15981_/B _22626_/X VGND VGND VPWR VPWR _23128_/D sky130_fd_sc_hd__o22a_4
XFILLER_59_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20747__A _20747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22561_ _22458_/X _22557_/X _15132_/B _22518_/X VGND VGND VPWR VPWR _23169_/D sky130_fd_sc_hd__o22a_4
XFILLER_35_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14745__A _13600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21512_ _21797_/A VGND VGND VPWR VPWR _21512_/X sky130_fd_sc_hd__buf_2
X_24300_ _24301_/CLK _24300_/D HRESETn VGND VGND VPWR VPWR _19121_/A sky130_fd_sc_hd__dfrtp_4
X_22492_ _22425_/X _22486_/X _13568_/B _22490_/X VGND VGND VPWR VPWR _23215_/D sky130_fd_sc_hd__o22a_4
X_21443_ _21287_/X _21440_/X _15290_/B _21437_/X VGND VGND VPWR VPWR _23810_/D sky130_fd_sc_hd__o22a_4
X_24231_ _24202_/CLK _24231_/D HRESETn VGND VGND VPWR VPWR _24231_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22455__A2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12265__A _12706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24162_ _24162_/CLK _19875_/X HRESETn VGND VGND VPWR VPWR _11633_/A sky130_fd_sc_hd__dfrtp_4
X_21374_ _21253_/X _21369_/X _13344_/B _21373_/X VGND VGND VPWR VPWR _23856_/D sky130_fd_sc_hd__o22a_4
X_20325_ _20301_/A VGND VGND VPWR VPWR _20325_/X sky130_fd_sc_hd__buf_2
X_23113_ _23433_/CLK _23113_/D VGND VGND VPWR VPWR _23113_/Q sky130_fd_sc_hd__dfxtp_4
X_24093_ _23485_/CLK _20316_/X VGND VGND VPWR VPWR _24093_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14480__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23044_ _22886_/X _23042_/X _17766_/A _23043_/X VGND VGND VPWR VPWR _23045_/B sky130_fd_sc_hd__o22a_4
Xclkbuf_7_126_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR _23157_/CLK sky130_fd_sc_hd__clkbuf_1
X_20256_ _18813_/X VGND VGND VPWR VPWR _20257_/B sky130_fd_sc_hd__inv_2
XFILLER_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18831__A1 _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20187_ _20187_/A VGND VGND VPWR VPWR _24109_/D sky130_fd_sc_hd__inv_2
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21718__B2 _21716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13824__A _15436_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11960_ _11959_/X VGND VGND VPWR VPWR _16150_/A sky130_fd_sc_hd__buf_2
X_23946_ _23915_/CLK _23946_/D VGND VGND VPWR VPWR _23946_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16200__A _11666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11891_ _12880_/A VGND VGND VPWR VPWR _15041_/A sky130_fd_sc_hd__buf_2
X_23877_ _23973_/CLK _23877_/D VGND VGND VPWR VPWR _14532_/B sky130_fd_sc_hd__dfxtp_4
X_13630_ _13630_/A _13630_/B VGND VGND VPWR VPWR _13631_/C sky130_fd_sc_hd__or2_4
XANTENNA__19511__A _19877_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22828_ _15051_/X _22826_/X _22827_/X VGND VGND VPWR VPWR _22828_/X sky130_fd_sc_hd__o21a_4
XFILLER_77_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23033__A _18050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13561_ _13561_/A _13487_/B VGND VGND VPWR VPWR _13561_/X sky130_fd_sc_hd__or2_4
XFILLER_53_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22759_ _22730_/Y _22758_/B VGND VGND VPWR VPWR _22759_/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22694__A2 _22693_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14655__A _14673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15300_ _14763_/A _15300_/B VGND VGND VPWR VPWR _15300_/X sky130_fd_sc_hd__or2_4
X_12512_ _12512_/A VGND VGND VPWR VPWR _13032_/A sky130_fd_sc_hd__buf_2
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16280_ _16252_/X _16280_/B VGND VGND VPWR VPWR _16280_/X sky130_fd_sc_hd__or2_4
XFILLER_9_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13492_ _11980_/X _13468_/X _13475_/X _13483_/X _13491_/X VGND VGND VPWR VPWR _13492_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_13_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15231_ _14190_/A _15227_/X _15230_/X VGND VGND VPWR VPWR _15231_/X sky130_fd_sc_hd__or3_4
X_12443_ _12443_/A _12564_/B VGND VGND VPWR VPWR _12443_/X sky130_fd_sc_hd__or2_4
X_24429_ _24334_/CLK _24429_/D HRESETn VGND VGND VPWR VPWR _20656_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_60_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20457__A1 _18162_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15162_ _14138_/X _15225_/B VGND VGND VPWR VPWR _15162_/X sky130_fd_sc_hd__or2_4
XANTENNA__21488__A _21467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21654__B1 _12827_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12374_ _12926_/A VGND VGND VPWR VPWR _12419_/A sky130_fd_sc_hd__buf_2
X_14113_ _14113_/A _14217_/B VGND VGND VPWR VPWR _14113_/X sky130_fd_sc_hd__or2_4
X_15093_ _15115_/A _15089_/X _15092_/X VGND VGND VPWR VPWR _15093_/X sky130_fd_sc_hd__or3_4
X_19970_ _19994_/A VGND VGND VPWR VPWR _19970_/X sky130_fd_sc_hd__buf_2
XFILLER_10_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23360__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12903__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21406__B1 _23837_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14044_ _14031_/A _23594_/Q VGND VGND VPWR VPWR _14044_/X sky130_fd_sc_hd__or2_4
X_18921_ _24350_/Q VGND VGND VPWR VPWR _20268_/A sky130_fd_sc_hd__inv_2
XANTENNA__21957__B2 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18852_ _17178_/X _18848_/X _24392_/Q _18849_/X VGND VGND VPWR VPWR _18852_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18822__A1 _11837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17803_ _17815_/A VGND VGND VPWR VPWR _17804_/A sky130_fd_sc_hd__buf_2
X_18783_ _17181_/X _18781_/X _24436_/Q _18782_/X VGND VGND VPWR VPWR _24436_/D sky130_fd_sc_hd__o22a_4
XFILLER_114_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15933__B _23256_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15995_ _16130_/A _15995_/B _15994_/X VGND VGND VPWR VPWR _15995_/X sky130_fd_sc_hd__or3_4
XFILLER_23_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22112__A _22112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17734_ _17734_/A _17111_/X VGND VGND VPWR VPWR _17734_/X sky130_fd_sc_hd__and2_4
XANTENNA__13734__A _15495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14946_ _14970_/A _14872_/B VGND VGND VPWR VPWR _14946_/X sky130_fd_sc_hd__or2_4
XFILLER_94_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21185__A2 _21183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17665_ _17665_/A _17685_/A VGND VGND VPWR VPWR _17665_/X sky130_fd_sc_hd__or2_4
X_14877_ _13985_/A _14875_/X _14877_/C VGND VGND VPWR VPWR _14878_/C sky130_fd_sc_hd__and3_4
X_16616_ _16616_/A _16614_/X _16615_/X VGND VGND VPWR VPWR _16616_/X sky130_fd_sc_hd__and3_4
X_19404_ _19403_/X _18598_/X _19403_/X _24198_/Q VGND VGND VPWR VPWR _19404_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13828_ _15443_/A _23079_/Q VGND VGND VPWR VPWR _13828_/X sky130_fd_sc_hd__or2_4
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17596_ _17409_/A VGND VGND VPWR VPWR _17601_/A sky130_fd_sc_hd__inv_2
XFILLER_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16547_ _16565_/A _23996_/Q VGND VGND VPWR VPWR _16548_/C sky130_fd_sc_hd__or2_4
X_19335_ _19317_/A VGND VGND VPWR VPWR _19336_/A sky130_fd_sc_hd__buf_2
XANTENNA__18889__A1 _12430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13759_ _12650_/A _13759_/B VGND VGND VPWR VPWR _13759_/X sky130_fd_sc_hd__or2_4
XFILLER_56_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22685__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14565__A _14563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19266_ _19220_/A _19220_/B _19265_/Y VGND VGND VPWR VPWR _24271_/D sky130_fd_sc_hd__o21a_4
X_16478_ _16203_/A _16478_/B _16477_/X VGND VGND VPWR VPWR _16479_/C sky130_fd_sc_hd__and3_4
XANTENNA__14284__B _14379_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18217_ _17446_/X _18217_/B VGND VGND VPWR VPWR _18217_/X sky130_fd_sc_hd__or2_4
X_15429_ _15429_/A _15493_/B VGND VGND VPWR VPWR _15429_/X sky130_fd_sc_hd__or2_4
X_19197_ _19197_/A VGND VGND VPWR VPWR _19197_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16780__A _16045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18148_ _17961_/X _18141_/Y _18076_/X _18147_/Y VGND VGND VPWR VPWR _18148_/X sky130_fd_sc_hd__a211o_4
XFILLER_7_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15396__A _13620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18079_ _17871_/A _18078_/Y VGND VGND VPWR VPWR _18079_/X sky130_fd_sc_hd__and2_4
XFILLER_102_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13909__A _13909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12813__A _12813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20110_ _11572_/X VGND VGND VPWR VPWR _20110_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21090_ _20637_/X _21089_/X _15724_/B _21086_/X VGND VGND VPWR VPWR _21090_/X sky130_fd_sc_hd__o22a_4
XFILLER_28_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23853__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21948__B2 _21942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20041_ _20041_/A VGND VGND VPWR VPWR _20041_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20620__A1 _20285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23800_ _24088_/CLK _23800_/D VGND VGND VPWR VPWR _23800_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13644__A _15443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17116__A _21583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21992_ _21985_/A VGND VGND VPWR VPWR _21992_/X sky130_fd_sc_hd__buf_2
XFILLER_2_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22373__B2 _22372_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23731_ _23986_/CLK _21606_/X VGND VGND VPWR VPWR _12929_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21861__A _21291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20943_ HRDATA[2] VGND VGND VPWR VPWR _20943_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _23342_/CLK _23662_/D VGND VGND VPWR VPWR _15737_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _20844_/A _20490_/B VGND VGND VPWR VPWR _20874_/X sky130_fd_sc_hd__or2_4
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22613_ _22462_/X _22586_/A _23135_/Q _22576_/A VGND VGND VPWR VPWR _23135_/D sky130_fd_sc_hd__o22a_4
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23593_ _23910_/CLK _21842_/X VGND VGND VPWR VPWR _23593_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14475__A _12533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20687__A1 _20494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22544_ _22427_/X _22543_/X _15659_/B _22540_/X VGND VGND VPWR VPWR _22544_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20687__B2 _20686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12707__B _23924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17786__A _18421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22475_ _22396_/X _22472_/X _16806_/B _22469_/X VGND VGND VPWR VPWR _23227_/D sky130_fd_sc_hd__o22a_4
X_24214_ _24239_/CLK _19376_/X HRESETn VGND VGND VPWR VPWR _24214_/Q sky130_fd_sc_hd__dfrtp_4
X_21426_ _21419_/A VGND VGND VPWR VPWR _21426_/X sky130_fd_sc_hd__buf_2
XFILLER_107_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18501__B1 _18500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21357_ _21225_/X _21355_/X _23868_/Q _21352_/X VGND VGND VPWR VPWR _23868_/D sky130_fd_sc_hd__o22a_4
X_24145_ _24250_/CLK _19920_/X HRESETn VGND VGND VPWR VPWR _24145_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12723__A _15664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20308_ _17636_/X _20578_/A _20290_/X _20307_/Y VGND VGND VPWR VPWR _20308_/X sky130_fd_sc_hd__a211o_4
X_12090_ _12086_/A _12159_/B VGND VGND VPWR VPWR _12092_/B sky130_fd_sc_hd__or2_4
X_21288_ _21287_/X _21283_/X _15273_/B _21278_/X VGND VGND VPWR VPWR _23906_/D sky130_fd_sc_hd__o22a_4
X_24076_ _23794_/CLK _20698_/X VGND VGND VPWR VPWR _15437_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21939__A1 _21816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21939__B2 _21935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20239_ _20516_/A VGND VGND VPWR VPWR _20492_/A sky130_fd_sc_hd__buf_2
X_23027_ _23027_/A _23027_/B VGND VGND VPWR VPWR _23027_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__18804__A1 _14564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24371__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23028__A _18087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14800_ _13706_/A _14796_/X _14799_/X VGND VGND VPWR VPWR _14800_/X sky130_fd_sc_hd__or3_4
XANTENNA__13554__A _13554_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15780_ _15713_/Y _15780_/B VGND VGND VPWR VPWR _15783_/A sky130_fd_sc_hd__and2_4
X_12992_ _12991_/Y VGND VGND VPWR VPWR _12992_/X sky130_fd_sc_hd__buf_2
XFILLER_57_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18568__B1 _18063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22364__A1 _22117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22364__B2 _22358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14369__B _14293_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14731_ _12531_/A _14727_/X _14731_/C VGND VGND VPWR VPWR _14731_/X sky130_fd_sc_hd__or3_4
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11943_ _11943_/A _24030_/Q VGND VGND VPWR VPWR _11946_/B sky130_fd_sc_hd__or2_4
X_23929_ _23770_/CLK _21233_/X VGND VGND VPWR VPWR _16263_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_40_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20914__A2 _20873_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17450_ _17037_/Y _17449_/X _17042_/A VGND VGND VPWR VPWR _17664_/B sky130_fd_sc_hd__o21a_4
X_14662_ _14672_/A _14662_/B VGND VGND VPWR VPWR _14663_/C sky130_fd_sc_hd__or2_4
XFILLER_72_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11874_ _16147_/A VGND VGND VPWR VPWR _16143_/A sky130_fd_sc_hd__buf_2
XFILLER_45_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16401_ _16397_/X _16401_/B VGND VGND VPWR VPWR _16401_/X sky130_fd_sc_hd__or2_4
XANTENNA__22116__B2 _22108_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13613_ _13606_/A VGND VGND VPWR VPWR _13614_/A sky130_fd_sc_hd__buf_2
X_17381_ _18418_/B VGND VGND VPWR VPWR _18428_/A sky130_fd_sc_hd__inv_2
XFILLER_92_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14593_ _12439_/A _14682_/B VGND VGND VPWR VPWR _14596_/B sky130_fd_sc_hd__or2_4
X_19120_ _19120_/A _19120_/B VGND VGND VPWR VPWR _19177_/A sky130_fd_sc_hd__and2_4
X_16332_ _16323_/A _23993_/Q VGND VGND VPWR VPWR _16332_/X sky130_fd_sc_hd__or2_4
XANTENNA__23726__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11802__A _16231_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13544_ _13511_/X _13544_/B _13543_/X VGND VGND VPWR VPWR _13545_/C sky130_fd_sc_hd__and3_4
XFILLER_9_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21875__B1 _23580_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19051_ _19046_/X _19050_/X _19046_/X _24330_/Q VGND VGND VPWR VPWR _24330_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16263_ _16090_/A _16263_/B VGND VGND VPWR VPWR _16263_/X sky130_fd_sc_hd__or2_4
X_13475_ _11861_/X _13471_/X _13475_/C VGND VGND VPWR VPWR _13475_/X sky130_fd_sc_hd__or3_4
XANTENNA__22419__A2 _22416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_8_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18002_ _17659_/X _17660_/X _17762_/X VGND VGND VPWR VPWR _18002_/X sky130_fd_sc_hd__or3_4
X_15214_ _14206_/A _15212_/X _15214_/C VGND VGND VPWR VPWR _15215_/C sky130_fd_sc_hd__and3_4
XANTENNA__21627__B1 _14654_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12426_ _15882_/A _12420_/X _12426_/C VGND VGND VPWR VPWR _12427_/C sky130_fd_sc_hd__or3_4
X_16194_ _16194_/A _16194_/B _16194_/C VGND VGND VPWR VPWR _16198_/B sky130_fd_sc_hd__and3_4
XANTENNA__22107__A _20590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23876__CLK _23107_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21011__A _21015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15145_ _14145_/A _15141_/X _15144_/X VGND VGND VPWR VPWR _15145_/X sky130_fd_sc_hd__or3_4
XFILLER_86_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13729__A _15497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12357_ _15743_/A _12355_/X _12357_/C VGND VGND VPWR VPWR _12363_/B sky130_fd_sc_hd__and3_4
XFILLER_5_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12633__A _12622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15076_ _15114_/A _15076_/B _15075_/X VGND VGND VPWR VPWR _15076_/X sky130_fd_sc_hd__and3_4
X_19953_ _19940_/X _19945_/Y _19947_/X _19951_/X _19952_/Y VGND VGND VPWR VPWR _19953_/X
+ sky130_fd_sc_hd__a32o_4
X_12288_ _12688_/A _12288_/B _12288_/C VGND VGND VPWR VPWR _12292_/B sky130_fd_sc_hd__and3_4
XANTENNA__12352__B _12224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14027_ _14035_/A _14027_/B VGND VGND VPWR VPWR _14027_/X sky130_fd_sc_hd__or2_4
X_18904_ _15646_/X _18898_/X _24363_/Q _18899_/X VGND VGND VPWR VPWR _24363_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23106__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15944__A _15939_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19416__A _22978_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19884_ _19379_/X VGND VGND VPWR VPWR _19884_/X sky130_fd_sc_hd__buf_2
XANTENNA__18320__A _18266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16759__B _16759_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18835_ _18835_/A VGND VGND VPWR VPWR _18835_/X sky130_fd_sc_hd__buf_2
XANTENNA__15663__B _15725_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13464__A _11913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15978_ _15957_/A _24056_/Q VGND VGND VPWR VPWR _15978_/X sky130_fd_sc_hd__or2_4
X_18766_ _18788_/A VGND VGND VPWR VPWR _18789_/A sky130_fd_sc_hd__inv_2
XFILLER_83_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22355__A1 _22100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21158__A2 _21154_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22355__B2 _22351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14279__B _14279_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14929_ _13998_/A _14929_/B _14929_/C VGND VGND VPWR VPWR _14934_/B sky130_fd_sc_hd__and3_4
X_17717_ _16969_/A _17385_/X _17713_/X VGND VGND VPWR VPWR _17747_/B sky130_fd_sc_hd__a21bo_4
XFILLER_58_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18697_ _18697_/A _17610_/Y VGND VGND VPWR VPWR _18697_/X sky130_fd_sc_hd__and2_4
XANTENNA__17231__B1 _14565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17648_ _17648_/A _17647_/X VGND VGND VPWR VPWR _17648_/Y sky130_fd_sc_hd__nor2_4
X_17579_ _17132_/Y _17781_/B _17271_/Y _17578_/X VGND VGND VPWR VPWR _18746_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22658__A2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11712__A _13257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20669__A1 _24205_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19318_ _19328_/A VGND VGND VPWR VPWR _19318_/X sky130_fd_sc_hd__buf_2
X_20590_ _20590_/A VGND VGND VPWR VPWR _20591_/A sky130_fd_sc_hd__buf_2
XANTENNA__24476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19249_ _19249_/A VGND VGND VPWR VPWR _19249_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22260_ _22079_/X _22258_/X _16608_/B _22255_/X VGND VGND VPWR VPWR _22260_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15838__B _15838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21211_ _23934_/Q VGND VGND VPWR VPWR _21211_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13639__A _12302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22191_ _22131_/X _22186_/X _23398_/Q _22190_/X VGND VGND VPWR VPWR _22191_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21094__B2 _21093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22291__B1 _14271_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21142_ _20671_/X _21140_/X _15799_/B _21137_/X VGND VGND VPWR VPWR _23981_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21073_ _20373_/X _21068_/X _16390_/B _21072_/X VGND VGND VPWR VPWR _24026_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15854__A _12413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20024_ _20000_/A VGND VGND VPWR VPWR _20024_/X sky130_fd_sc_hd__buf_2
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22594__B2 _22590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16669__B _23484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15573__B _15573_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21149__A2 _21147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_14_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21591__A _21605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21975_ _21791_/X _21974_/X _23517_/Q _21971_/X VGND VGND VPWR VPWR _23517_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20919__B _20358_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23714_ _24066_/CLK _23714_/D VGND VGND VPWR VPWR _15256_/B sky130_fd_sc_hd__dfxtp_4
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _20255_/A _20925_/X _19094_/A _18870_/X VGND VGND VPWR VPWR _20926_/X sky130_fd_sc_hd__o22a_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17773__B2 _11629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _23515_/CLK _21742_/X VGND VGND VPWR VPWR _23645_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19996__A _19996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20109__B1 _19380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ _20654_/X _20854_/Y _20856_/X _19079_/Y _20709_/X VGND VGND VPWR VPWR _20858_/A
+ sky130_fd_sc_hd__a32o_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22649__A2 _22643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20000__A _20000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12718__A _12284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11622__A _11622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ _17262_/A _17273_/A _17040_/A _17028_/A VGND VGND VPWR VPWR _11591_/D sky130_fd_sc_hd__or4_4
X_23576_ _23539_/CLK _21881_/X VGND VGND VPWR VPWR _23576_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20788_ _20733_/X _20787_/X _24328_/Q _20686_/X VGND VGND VPWR VPWR _20788_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21321__A2 _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22527_ _22398_/X _22522_/X _16387_/B _22526_/X VGND VGND VPWR VPWR _23194_/D sky130_fd_sc_hd__o22a_4
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14933__A _15063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13260_ _13260_/A _23473_/Q VGND VGND VPWR VPWR _13262_/B sky130_fd_sc_hd__or2_4
XANTENNA__24146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22458_ _22458_/A VGND VGND VPWR VPWR _22458_/X sky130_fd_sc_hd__buf_2
XANTENNA__15748__B _15748_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12211_ _12211_/A VGND VGND VPWR VPWR _12211_/X sky130_fd_sc_hd__buf_2
XFILLER_109_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21409_ _21401_/X VGND VGND VPWR VPWR _21409_/X sky130_fd_sc_hd__buf_2
XANTENNA__13549__A _13548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21085__B2 _21079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22282__B1 _15458_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13191_ _12849_/A _13188_/X _13190_/X VGND VGND VPWR VPWR _13191_/X sky130_fd_sc_hd__and3_4
XANTENNA__12453__A _12850_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22389_ _22382_/Y _22387_/X _22388_/X _22387_/X VGND VGND VPWR VPWR _22389_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20832__A1 _18594_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12142_ _11747_/X _12138_/X _12141_/X VGND VGND VPWR VPWR _12142_/X sky130_fd_sc_hd__or3_4
X_24128_ _24066_/CLK _24128_/D HRESETn VGND VGND VPWR VPWR _24128_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21766__A _21752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20670__A _20670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15764__A _12777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22034__B1 _12312_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12073_ _12096_/A _12073_/B _12073_/C VGND VGND VPWR VPWR _12073_/X sky130_fd_sc_hd__or3_4
X_16950_ _24126_/Q VGND VGND VPWR VPWR _17681_/A sky130_fd_sc_hd__inv_2
X_24059_ _24059_/CLK _21019_/X VGND VGND VPWR VPWR _24059_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22585__A1 _22413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21388__A2 _21383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22585__B2 _22583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16579__B _23484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15901_ _13561_/A _15831_/B VGND VGND VPWR VPWR _15901_/X sky130_fd_sc_hd__or2_4
XFILLER_81_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23279__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16881_ _15928_/X _16239_/B _16236_/X VGND VGND VPWR VPWR _16881_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15832_ _12874_/A _15902_/B VGND VGND VPWR VPWR _15832_/X sky130_fd_sc_hd__or2_4
X_18620_ _18714_/A _17605_/A _17782_/Y VGND VGND VPWR VPWR _18620_/X sky130_fd_sc_hd__a21o_4
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22597__A _22583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15763_ _15751_/A _15763_/B VGND VGND VPWR VPWR _15763_/X sky130_fd_sc_hd__or2_4
X_18551_ _17716_/X _18550_/X _17716_/X _18550_/X VGND VGND VPWR VPWR _18551_/X sky130_fd_sc_hd__a2bb2o_4
X_12975_ _12951_/A _12975_/B _12975_/C VGND VGND VPWR VPWR _12979_/B sky130_fd_sc_hd__and3_4
X_14714_ _14714_/A _14714_/B VGND VGND VPWR VPWR _14715_/C sky130_fd_sc_hd__or2_4
X_17502_ _17500_/Y _17501_/X VGND VGND VPWR VPWR _17502_/X sky130_fd_sc_hd__or2_4
X_11926_ _11925_/Y VGND VGND VPWR VPWR _12301_/A sky130_fd_sc_hd__buf_2
X_18482_ _18349_/A _16972_/B _18460_/Y VGND VGND VPWR VPWR _22944_/B sky130_fd_sc_hd__a21oi_4
X_15694_ _12705_/A _15692_/X _15694_/C VGND VGND VPWR VPWR _15694_/X sky130_fd_sc_hd__and3_4
XFILLER_72_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17433_ _17382_/B _17431_/Y _17432_/X VGND VGND VPWR VPWR _17433_/X sky130_fd_sc_hd__o21a_4
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14645_ _15105_/A _14569_/B VGND VGND VPWR VPWR _14645_/X sky130_fd_sc_hd__or2_4
XFILLER_72_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11857_ _13972_/A VGND VGND VPWR VPWR _15449_/A sky130_fd_sc_hd__buf_2
XFILLER_61_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15004__A _15023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17364_ _17364_/A VGND VGND VPWR VPWR _17364_/X sky130_fd_sc_hd__buf_2
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14576_ _14575_/X _14654_/B VGND VGND VPWR VPWR _14577_/C sky130_fd_sc_hd__or2_4
X_11788_ _12169_/A _11788_/B _11787_/X VGND VGND VPWR VPWR _11793_/B sky130_fd_sc_hd__and3_4
Xclkbuf_7_34_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR _23845_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_41_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12347__B _12213_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16315_ _16188_/A _16249_/B VGND VGND VPWR VPWR _16316_/C sky130_fd_sc_hd__or2_4
X_19103_ _18971_/A _19101_/Y _24320_/Q _19102_/X VGND VGND VPWR VPWR _24320_/D sky130_fd_sc_hd__a2bb2o_4
X_13527_ _12754_/X _13527_/B _13527_/C VGND VGND VPWR VPWR _13528_/C sky130_fd_sc_hd__and3_4
XANTENNA__15939__A _15939_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_97_0_HCLK clkbuf_6_48_0_HCLK/X VGND VGND VPWR VPWR _23130_/CLK sky130_fd_sc_hd__clkbuf_1
X_17295_ _14564_/X _17295_/B VGND VGND VPWR VPWR _17295_/X sky130_fd_sc_hd__or2_4
XFILLER_105_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14843__A _12575_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19034_ _24365_/Q VGND VGND VPWR VPWR _19034_/Y sky130_fd_sc_hd__inv_2
X_16246_ _16151_/A _16244_/X _16245_/X VGND VGND VPWR VPWR _16246_/X sky130_fd_sc_hd__and3_4
X_13458_ _12870_/A _13458_/B _13458_/C VGND VGND VPWR VPWR _13459_/C sky130_fd_sc_hd__and3_4
XFILLER_16_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12409_ _12418_/A _12328_/B VGND VGND VPWR VPWR _12409_/X sky130_fd_sc_hd__or2_4
XFILLER_115_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13459__A _12528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21076__B2 _21072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16177_ _16193_/A _16103_/B VGND VGND VPWR VPWR _16177_/X sky130_fd_sc_hd__or2_4
XFILLER_115_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13389_ _11681_/X _13389_/B _13389_/C VGND VGND VPWR VPWR _13389_/X sky130_fd_sc_hd__or3_4
XANTENNA__12363__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15128_ _14083_/A _15128_/B VGND VGND VPWR VPWR _15128_/X sky130_fd_sc_hd__or2_4
XANTENNA__21676__A _21636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__15674__A _12240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15059_ _14037_/A _15054_/X _15058_/X VGND VGND VPWR VPWR _15068_/B sky130_fd_sc_hd__or3_4
X_19936_ _19936_/A VGND VGND VPWR VPWR _19936_/X sky130_fd_sc_hd__buf_2
XANTENNA__21379__A2 _21376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16489__B _16489_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15393__B _15455_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19867_ _19793_/A _19867_/B _19867_/C _19880_/B VGND VGND VPWR VPWR _19867_/X sky130_fd_sc_hd__and4_4
XFILLER_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20587__B1 _20586_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13194__A _12315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18818_ _18834_/A VGND VGND VPWR VPWR _18818_/X sky130_fd_sc_hd__buf_2
XANTENNA__19992__A2 _16985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19798_ _19449_/X _19793_/X _19797_/Y _16907_/C _19490_/X VGND VGND VPWR VPWR _19798_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_110_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18749_ _18745_/Y _18747_/X _18744_/X _18748_/X VGND VGND VPWR VPWR _18750_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21000__A1 _24191_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21760_ _21538_/X _21755_/X _13337_/B _21759_/X VGND VGND VPWR VPWR _23632_/D sky130_fd_sc_hd__o22a_4
XFILLER_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20711_ _20710_/X VGND VGND VPWR VPWR _20711_/Y sky130_fd_sc_hd__inv_2
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21691_ _21705_/A VGND VGND VPWR VPWR _21691_/X sky130_fd_sc_hd__buf_2
XANTENNA__12538__A _12497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23430_ _23781_/CLK _23430_/D VGND VGND VPWR VPWR _14296_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20642_ _20641_/X VGND VGND VPWR VPWR _20642_/X sky130_fd_sc_hd__buf_2
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17507__A1 _17504_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17507__B2 _17506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20573_ _20573_/A VGND VGND VPWR VPWR _20574_/A sky130_fd_sc_hd__buf_2
X_23361_ _24032_/CLK _23361_/D VGND VGND VPWR VPWR _15228_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15849__A _13548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14753__A _11976_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22312_ _23314_/Q VGND VGND VPWR VPWR _22312_/X sky130_fd_sc_hd__buf_2
X_23292_ _23100_/CLK _22342_/X VGND VGND VPWR VPWR _16620_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_30_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22243_ _22207_/A VGND VGND VPWR VPWR _22243_/X sky130_fd_sc_hd__buf_2
XANTENNA__22264__B1 _16244_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12273__A _12233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22174_ _22103_/X _22172_/X _13039_/B _22169_/X VGND VGND VPWR VPWR _22174_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21586__A _21590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20490__A _20342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21125_ _20394_/X _21119_/X _23993_/Q _21123_/X VGND VGND VPWR VPWR _23993_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21056_ _20982_/X _21051_/X _14892_/B _21012_/X VGND VGND VPWR VPWR _21056_/X sky130_fd_sc_hd__o22a_4
XFILLER_101_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20007_ _19994_/X _16946_/Y _20000_/X _20006_/X VGND VGND VPWR VPWR _20007_/X sky130_fd_sc_hd__o22a_4
XFILLER_115_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11617__A _13595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17304__A _17297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12760_ _13065_/A VGND VGND VPWR VPWR _13130_/A sky130_fd_sc_hd__buf_2
XFILLER_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _21850_/X _21952_/X _14450_/B _21956_/X VGND VGND VPWR VPWR _21958_/X sky130_fd_sc_hd__o22a_4
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21542__A2 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _12373_/A VGND VGND VPWR VPWR _13257_/A sky130_fd_sc_hd__buf_2
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _18664_/X _20291_/X _20758_/X _20908_/Y VGND VGND VPWR VPWR _20910_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24398__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12691_/A _12774_/B VGND VGND VPWR VPWR _12692_/C sky130_fd_sc_hd__or2_4
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _21819_/X _21887_/X _13085_/B _21884_/X VGND VGND VPWR VPWR _21889_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12448__A _14748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14427_/Y _14430_/B VGND VGND VPWR VPWR _14430_/X sky130_fd_sc_hd__or2_4
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11642_/A VGND VGND VPWR VPWR _15114_/A sky130_fd_sc_hd__buf_2
X_23628_ _23564_/CLK _23628_/D VGND VGND VPWR VPWR _15512_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _13844_/A VGND VGND VPWR VPWR _14379_/A sky130_fd_sc_hd__buf_2
XANTENNA__15759__A _12765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11573_ _11569_/X _11570_/X _11572_/X VGND VGND VPWR VPWR _20090_/A sky130_fd_sc_hd__or3_4
X_23559_ _23591_/CLK _23559_/D VGND VGND VPWR VPWR _23559_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24077__CLK _23922_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18135__A _18205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14663__A _15107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16100_ _13283_/X VGND VGND VPWR VPWR _16100_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _15697_/A _13312_/B VGND VGND VPWR VPWR _13312_/X sky130_fd_sc_hd__or2_4
XFILLER_35_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17080_ _18025_/A VGND VGND VPWR VPWR _17900_/A sky130_fd_sc_hd__inv_2
X_14292_ _13678_/A _14292_/B VGND VGND VPWR VPWR _14292_/X sky130_fd_sc_hd__or2_4
XFILLER_10_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16031_ _16047_/A _23576_/Q VGND VGND VPWR VPWR _16032_/C sky130_fd_sc_hd__or2_4
X_13243_ _13243_/A _13243_/B _13243_/C VGND VGND VPWR VPWR _13244_/C sky130_fd_sc_hd__and3_4
XFILLER_109_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12183__A _16077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13174_ _12728_/A _13174_/B VGND VGND VPWR VPWR _13174_/X sky130_fd_sc_hd__or2_4
XANTENNA__17693__B _17367_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12125_ _12168_/A _23741_/Q VGND VGND VPWR VPWR _12126_/C sky130_fd_sc_hd__or2_4
XFILLER_69_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15494__A _15494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22007__B1 _14269_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17982_ _17911_/X _17848_/X _17912_/X _17841_/X VGND VGND VPWR VPWR _17982_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__12911__A _12497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22558__B2 _22554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19721_ _19740_/B VGND VGND VPWR VPWR _19721_/Y sky130_fd_sc_hd__inv_2
X_12056_ _11943_/A VGND VGND VPWR VPWR _12086_/A sky130_fd_sc_hd__buf_2
X_16933_ _16933_/A VGND VGND VPWR VPWR _18171_/A sky130_fd_sc_hd__buf_2
X_19652_ _19447_/X _19651_/X _17299_/Y _19493_/X VGND VGND VPWR VPWR _19652_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__19974__A2 _17766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16864_ _15388_/X _14568_/Y _16863_/Y _14567_/X VGND VGND VPWR VPWR _16865_/D sky130_fd_sc_hd__o22a_4
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21781__A2 _21776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18603_ _20077_/D VGND VGND VPWR VPWR _18603_/Y sky130_fd_sc_hd__inv_2
X_15815_ _12444_/A _15815_/B VGND VGND VPWR VPWR _15815_/X sky130_fd_sc_hd__or2_4
X_16795_ _16624_/X _16787_/X _16795_/C VGND VGND VPWR VPWR _16795_/X sky130_fd_sc_hd__and3_4
X_19583_ _19582_/Y _19766_/A VGND VGND VPWR VPWR _19583_/X sky130_fd_sc_hd__and2_4
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14838__A _14845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22120__A _22108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13742__A _13697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15746_ _12957_/A _15746_/B _15745_/X VGND VGND VPWR VPWR _15746_/X sky130_fd_sc_hd__or3_4
X_18534_ _18533_/A _16970_/B _18515_/Y VGND VGND VPWR VPWR _22932_/B sky130_fd_sc_hd__a21oi_4
XFILLER_34_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12958_ _12958_/A _23891_/Q VGND VGND VPWR VPWR _12958_/X sky130_fd_sc_hd__or2_4
XFILLER_59_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21533__A2 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20852__A1_N _19699_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11909_ _11909_/A VGND VGND VPWR VPWR _15578_/A sky130_fd_sc_hd__buf_2
X_15677_ _12743_/A _15677_/B VGND VGND VPWR VPWR _15678_/C sky130_fd_sc_hd__or2_4
X_18465_ _18295_/A _17348_/B VGND VGND VPWR VPWR _18468_/B sky130_fd_sc_hd__nor2_4
X_12889_ _13029_/A _23443_/Q VGND VGND VPWR VPWR _12890_/C sky130_fd_sc_hd__or2_4
XANTENNA__12358__A _12421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14628_ _12883_/A _14714_/B VGND VGND VPWR VPWR _14628_/X sky130_fd_sc_hd__or2_4
X_17416_ _17416_/A VGND VGND VPWR VPWR _18525_/B sky130_fd_sc_hd__inv_2
X_18396_ _17592_/X _18395_/X VGND VGND VPWR VPWR _18396_/X sky130_fd_sc_hd__and2_4
XFILLER_33_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17347_ _17339_/Y _17340_/X _17020_/A _17346_/X VGND VGND VPWR VPWR _17348_/B sky130_fd_sc_hd__o22a_4
XANTENNA__15669__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14559_ _13699_/A _14557_/X _14559_/C VGND VGND VPWR VPWR _14560_/C sky130_fd_sc_hd__and3_4
XANTENNA__22494__B1 _15699_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14573__A _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17278_ _17277_/X _17278_/B VGND VGND VPWR VPWR _17278_/X sky130_fd_sc_hd__and2_4
XANTENNA__22790__A _17283_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23444__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14292__B _14292_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16229_ _16229_/A _16229_/B _16228_/X VGND VGND VPWR VPWR _16230_/C sky130_fd_sc_hd__or3_4
X_19017_ _19002_/X _19015_/X _19016_/X _24336_/Q VGND VGND VPWR VPWR _19017_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13189__A _15707_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21049__B2 _21048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13917__A _11799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23594__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12821__A _12753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22549__B2 _22547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19919_ _19916_/X _24146_/Q _19917_/X _20895_/B VGND VGND VPWR VPWR _24146_/D sky130_fd_sc_hd__o22a_4
XFILLER_69_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22930_ _22924_/X _16998_/A _22887_/X _22929_/X VGND VGND VPWR VPWR _22931_/A sky130_fd_sc_hd__a211o_4
XFILLER_60_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17976__B2 _17827_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21772__A2 _21769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22861_ _22813_/X _22861_/B VGND VGND VPWR VPWR HWDATA[25] sky130_fd_sc_hd__nor2_4
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14748__A _14748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13652__A _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21812_ _21812_/A VGND VGND VPWR VPWR _21812_/X sky130_fd_sc_hd__buf_2
X_22792_ _22862_/A VGND VGND VPWR VPWR _22792_/X sky130_fd_sc_hd__buf_2
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21743_ _21510_/X _21741_/X _23644_/Q _21738_/X VGND VGND VPWR VPWR _23644_/D sky130_fd_sc_hd__o22a_4
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12268__A _12267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24462_ _24126_/CLK _24462_/D HRESETn VGND VGND VPWR VPWR _24462_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21674_ _21562_/X _21669_/X _14330_/B _21673_/X VGND VGND VPWR VPWR _23686_/D sky130_fd_sc_hd__o22a_4
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23413_ _23635_/CLK _22170_/X VGND VGND VPWR VPWR _12653_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20625_ _20407_/A VGND VGND VPWR VPWR _20625_/X sky130_fd_sc_hd__buf_2
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15579__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21288__B2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24393_ _24365_/CLK _18851_/X HRESETn VGND VGND VPWR VPWR _24393_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14483__A _13614_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11900__A _15956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23344_ _23920_/CLK _23344_/D VGND VGND VPWR VPWR _13287_/B sky130_fd_sc_hd__dfxtp_4
X_20556_ _20556_/A VGND VGND VPWR VPWR _20595_/B sky130_fd_sc_hd__buf_2
Xclkbuf_7_80_0_HCLK clkbuf_6_40_0_HCLK/X VGND VGND VPWR VPWR _24425_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23275_ _24011_/CLK _23275_/D VGND VGND VPWR VPWR _23275_/Q sky130_fd_sc_hd__dfxtp_4
X_20487_ _20487_/A VGND VGND VPWR VPWR _20487_/X sky130_fd_sc_hd__buf_2
XFILLER_69_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22226_ _22219_/A VGND VGND VPWR VPWR _22226_/X sky130_fd_sc_hd__buf_2
XFILLER_118_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22205__A _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14930__B _14866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13827__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22157_ _22153_/A VGND VGND VPWR VPWR _22172_/A sky130_fd_sc_hd__buf_2
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16203__A _16203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12731__A _12705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21108_ _20982_/X _21103_/X _14866_/B _21072_/A VGND VGND VPWR VPWR _24000_/D sky130_fd_sc_hd__o22a_4
X_22088_ _20418_/A VGND VGND VPWR VPWR _22088_/X sky130_fd_sc_hd__buf_2
XFILLER_59_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13930_ _15036_/A _23338_/Q VGND VGND VPWR VPWR _13932_/B sky130_fd_sc_hd__or2_4
XFILLER_87_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21039_ _20671_/X _21037_/X _15818_/B _21034_/X VGND VGND VPWR VPWR _21039_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21763__A2 _21762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13861_ _14810_/A VGND VGND VPWR VPWR _13862_/A sky130_fd_sc_hd__buf_2
XFILLER_21_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15600_ _15616_/A _15600_/B _15599_/X VGND VGND VPWR VPWR _15600_/X sky130_fd_sc_hd__and3_4
X_12812_ _12800_/A _24052_/Q VGND VGND VPWR VPWR _12813_/C sky130_fd_sc_hd__or2_4
X_16580_ _16583_/A _24092_/Q VGND VGND VPWR VPWR _16581_/C sky130_fd_sc_hd__or2_4
X_13792_ _15430_/A _13792_/B VGND VGND VPWR VPWR _13792_/X sky130_fd_sc_hd__or2_4
XFILLER_28_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22712__A1 _21291_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15531_ _12307_/A _15529_/X _15530_/X VGND VGND VPWR VPWR _15531_/X sky130_fd_sc_hd__and3_4
XANTENNA__22712__B2 _22668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12743_ _12743_/A _23796_/Q VGND VGND VPWR VPWR _12743_/X sky130_fd_sc_hd__or2_4
XFILLER_16_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18250_ _17796_/X _17984_/X _17964_/X VGND VGND VPWR VPWR _18250_/X sky130_fd_sc_hd__o21a_4
X_15462_ _15486_/A _15462_/B VGND VGND VPWR VPWR _15462_/X sky130_fd_sc_hd__or2_4
XFILLER_19_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12674_ _12673_/X VGND VGND VPWR VPWR _12674_/X sky130_fd_sc_hd__buf_2
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17688__B _17688_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17201_/A VGND VGND VPWR VPWR _17256_/A sky130_fd_sc_hd__buf_2
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _13847_/A VGND VGND VPWR VPWR _15617_/A sky130_fd_sc_hd__buf_2
XANTENNA__21279__A1 _21277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _11625_/A _11624_/X VGND VGND VPWR VPWR _11625_/X sky130_fd_sc_hd__and2_4
X_18181_ _18180_/X VGND VGND VPWR VPWR _18181_/Y sky130_fd_sc_hd__inv_2
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15489__A _13735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21279__B2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _15393_/A _15455_/B VGND VGND VPWR VPWR _15394_/C sky130_fd_sc_hd__or2_4
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17701__A2_N _17354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17132_ _16678_/X VGND VGND VPWR VPWR _17132_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11810__A _11803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ _15623_/A _14341_/X _14344_/C VGND VGND VPWR VPWR _14344_/X sky130_fd_sc_hd__and3_4
XFILLER_11_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _20762_/A IRQ[10] VGND VGND VPWR VPWR _11556_/X sky130_fd_sc_hd__and2_4
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17063_ _17063_/A VGND VGND VPWR VPWR _17145_/A sky130_fd_sc_hd__inv_2
X_14275_ _12257_/A _14275_/B VGND VGND VPWR VPWR _14275_/X sky130_fd_sc_hd__or2_4
XANTENNA__22779__A1 _18720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16014_ _16019_/A _23352_/Q VGND VGND VPWR VPWR _16014_/X sky130_fd_sc_hd__or2_4
X_13226_ _13243_/A _13224_/X _13226_/C VGND VGND VPWR VPWR _13226_/X sky130_fd_sc_hd__and3_4
XANTENNA__22115__A _20670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13737__A _13737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13157_ _15696_/A _13157_/B VGND VGND VPWR VPWR _13157_/X sky130_fd_sc_hd__or2_4
XFILLER_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12641__A _12982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16113__A _16113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12108_ _16541_/A _12108_/B _12108_/C VGND VGND VPWR VPWR _12108_/X sky130_fd_sc_hd__and3_4
XFILLER_97_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13456__B _13456_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13088_ _13088_/A VGND VGND VPWR VPWR _13098_/A sky130_fd_sc_hd__buf_2
X_17965_ _17962_/X _17963_/X _17964_/X VGND VGND VPWR VPWR _17965_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__12360__B _12236_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19704_ _19663_/A _19703_/X _19877_/A VGND VGND VPWR VPWR _19704_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__20006__A2 _19985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12039_ _11888_/A VGND VGND VPWR VPWR _16713_/A sky130_fd_sc_hd__buf_2
X_16916_ _16916_/A _16916_/B _17083_/A _16890_/X VGND VGND VPWR VPWR _16917_/C sky130_fd_sc_hd__or4_4
XANTENNA__21203__B2 _21201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22400__B1 _16380_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17896_ _17896_/A _17895_/Y VGND VGND VPWR VPWR _17896_/X sky130_fd_sc_hd__and2_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21754__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19635_ _19612_/A _19624_/Y _19627_/Y _19634_/X VGND VGND VPWR VPWR _19635_/X sky130_fd_sc_hd__or4_4
XFILLER_77_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16847_ _13280_/B _16832_/X _13280_/B _16832_/X VGND VGND VPWR VPWR _16847_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20962__B1 HRDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13472__A _13448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19566_ _19517_/A _19511_/B _19729_/C VGND VGND VPWR VPWR _19566_/X sky130_fd_sc_hd__or3_4
XANTENNA__24242__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16778_ _16598_/X _16778_/B _16777_/X VGND VGND VPWR VPWR _16779_/C sky130_fd_sc_hd__or3_4
XFILLER_111_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_5_23_0_HCLK_A clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22785__A _17115_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22703__B2 _22697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18517_ _18097_/A _18349_/B _18514_/Y _18016_/A _22939_/B VGND VGND VPWR VPWR _18517_/X
+ sky130_fd_sc_hd__a32o_4
X_15729_ _15724_/A _15729_/B VGND VGND VPWR VPWR _15729_/X sky130_fd_sc_hd__or2_4
X_19497_ _19712_/A VGND VGND VPWR VPWR _19497_/X sky130_fd_sc_hd__buf_2
XFILLER_34_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16783__A _11823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24348__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18448_ _18466_/B _18395_/C VGND VGND VPWR VPWR _18448_/X sky130_fd_sc_hd__or2_4
XFILLER_37_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18379_ _18340_/X _18376_/X _18377_/X _18378_/X VGND VGND VPWR VPWR _18379_/X sky130_fd_sc_hd__o22a_4
XFILLER_18_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20410_ _20322_/X _20409_/X _24344_/Q _20247_/X VGND VGND VPWR VPWR _20410_/X sky130_fd_sc_hd__o22a_4
X_21390_ _21383_/A VGND VGND VPWR VPWR _21390_/X sky130_fd_sc_hd__buf_2
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18686__A2 _17111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20341_ _18757_/X VGND VGND VPWR VPWR _20342_/A sky130_fd_sc_hd__buf_2
XANTENNA__18503__A _18697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20272_ _20272_/A VGND VGND VPWR VPWR _20272_/Y sky130_fd_sc_hd__inv_2
X_23060_ _23060_/A VGND VGND VPWR VPWR HADDR[31] sky130_fd_sc_hd__inv_2
XANTENNA__15846__B _23501_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22011_ _21855_/X _22009_/X _14788_/B _22006_/X VGND VGND VPWR VPWR _23491_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13647__A _13647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12551__A _13032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21442__B2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21993__A2 _21988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15862__A _13522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23962_ _23632_/CLK _21174_/X VGND VGND VPWR VPWR _23962_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13683__A1 _11977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22913_ _23051_/A _22913_/B _22912_/X VGND VGND VPWR VPWR _22917_/B sky130_fd_sc_hd__or3_4
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23893_ _23315_/CLK _23893_/D VGND VGND VPWR VPWR _12639_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14478__A _13054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22844_ _17298_/Y _22778_/Y _22794_/A VGND VGND VPWR VPWR _22844_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17789__A _17779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22775_ _22774_/X VGND VGND VPWR VPWR _24103_/D sky130_fd_sc_hd__inv_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22170__A2 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21726_ _21690_/A VGND VGND VPWR VPWR _21726_/X sky130_fd_sc_hd__buf_2
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20181__B2 _19929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24445_ _24435_/CLK _24445_/D HRESETn VGND VGND VPWR VPWR _20297_/A sky130_fd_sc_hd__dfrtp_4
X_21657_ _21534_/X _21655_/X _13122_/B _21652_/X VGND VGND VPWR VPWR _21657_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12726__A _12726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20608_ _20534_/A _20607_/X VGND VGND VPWR VPWR _20608_/X sky130_fd_sc_hd__or2_4
XFILLER_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12390_ _13557_/A _12390_/B _12390_/C VGND VGND VPWR VPWR _12390_/X sky130_fd_sc_hd__and3_4
X_24376_ _24435_/CLK _18887_/X HRESETn VGND VGND VPWR VPWR _24376_/Q sky130_fd_sc_hd__dfstp_4
X_21588_ _21595_/A VGND VGND VPWR VPWR _21588_/X sky130_fd_sc_hd__buf_2
XANTENNA__20943__A HRDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23327_ _23487_/CLK _23327_/D VGND VGND VPWR VPWR _15056_/B sky130_fd_sc_hd__dfxtp_4
X_20539_ _20285_/X _20539_/B VGND VGND VPWR VPWR _20539_/X sky130_fd_sc_hd__and2_4
XANTENNA__21681__B2 _21637_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14941__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14060_ _14035_/A _23850_/Q VGND VGND VPWR VPWR _14060_/X sky130_fd_sc_hd__or2_4
X_23258_ _23354_/CLK _22400_/X VGND VGND VPWR VPWR _16380_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_101_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24115__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13011_ _12891_/A _13007_/X _13011_/C VGND VGND VPWR VPWR _13011_/X sky130_fd_sc_hd__or3_4
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18132__B _18174_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22209_ _22075_/X _22208_/X _12162_/B _22205_/X VGND VGND VPWR VPWR _22209_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13557__A _13557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17029__A _17040_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22630__B1 _15981_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23189_ _23987_/CLK _22534_/X VGND VGND VPWR VPWR _12462_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12461__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15772__A _12792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14962_ _12340_/A _14962_/B VGND VGND VPWR VPWR _14962_/X sky130_fd_sc_hd__or2_4
X_17750_ _17706_/X _17710_/X _17748_/X _17705_/Y _17749_/Y VGND VGND VPWR VPWR _17750_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_88_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16701_ _12091_/A _23547_/Q VGND VGND VPWR VPWR _16702_/C sky130_fd_sc_hd__or2_4
XFILLER_75_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13913_ _13718_/A _13825_/B VGND VGND VPWR VPWR _13914_/C sky130_fd_sc_hd__or2_4
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14893_ _13982_/A _14891_/X _14892_/X VGND VGND VPWR VPWR _14893_/X sky130_fd_sc_hd__and3_4
X_17681_ _17681_/A _17487_/X VGND VGND VPWR VPWR _17758_/A sky130_fd_sc_hd__and2_4
XANTENNA__20944__B1 _20939_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19420_ _16996_/A _19430_/B VGND VGND VPWR VPWR _19462_/A sky130_fd_sc_hd__or2_4
XFILLER_21_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11805__A _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13844_ _13844_/A VGND VGND VPWR VPWR _13845_/A sky130_fd_sc_hd__buf_2
X_16632_ _16618_/X VGND VGND VPWR VPWR _16670_/A sky130_fd_sc_hd__buf_2
XFILLER_74_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19351_ _19347_/X _18648_/X _19350_/X _20888_/A VGND VGND VPWR VPWR _19351_/X sky130_fd_sc_hd__a2bb2o_4
X_13775_ _13774_/X VGND VGND VPWR VPWR _13775_/Y sky130_fd_sc_hd__inv_2
X_16563_ _16741_/A _16533_/X _16542_/X _16554_/X _16562_/X VGND VGND VPWR VPWR _16563_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18302_ _18301_/X VGND VGND VPWR VPWR _18446_/B sky130_fd_sc_hd__inv_2
X_12726_ _12726_/A _23828_/Q VGND VGND VPWR VPWR _12727_/C sky130_fd_sc_hd__or2_4
X_15514_ _12613_/A _15514_/B _15514_/C VGND VGND VPWR VPWR _15515_/C sky130_fd_sc_hd__or3_4
X_16494_ _16506_/A _16494_/B _16493_/X VGND VGND VPWR VPWR _16495_/C sky130_fd_sc_hd__and3_4
X_19282_ _19212_/A _19212_/B _19281_/Y VGND VGND VPWR VPWR _19282_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17640__A2_N _17044_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15445_ _13677_/A _15443_/X _15445_/C VGND VGND VPWR VPWR _15449_/B sky130_fd_sc_hd__and3_4
X_18233_ _24126_/Q _18233_/B VGND VGND VPWR VPWR _18234_/B sky130_fd_sc_hd__and2_4
X_12657_ _12604_/A _12657_/B VGND VGND VPWR VPWR _12657_/X sky130_fd_sc_hd__or2_4
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12636__A _13118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ _11608_/A VGND VGND VPWR VPWR _12860_/A sky130_fd_sc_hd__buf_2
X_15376_ _14008_/A _15372_/X _15376_/C VGND VGND VPWR VPWR _15377_/C sky130_fd_sc_hd__or3_4
X_18164_ _18164_/A VGND VGND VPWR VPWR _18285_/C sky130_fd_sc_hd__buf_2
XANTENNA__21949__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12588_ _12655_/A _12572_/X _12587_/X VGND VGND VPWR VPWR _12588_/X sky130_fd_sc_hd__or3_4
XANTENNA__21121__B1 _23996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19865__B2 _19531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12355__B _12228_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ _15543_/A _14327_/B VGND VGND VPWR VPWR _14327_/X sky130_fd_sc_hd__or2_4
X_17115_ _15185_/X VGND VGND VPWR VPWR _17115_/Y sky130_fd_sc_hd__inv_2
X_11539_ _20966_/A IRQ[1] VGND VGND VPWR VPWR _11539_/X sky130_fd_sc_hd__and2_4
X_18095_ _18342_/A VGND VGND VPWR VPWR _18097_/A sky130_fd_sc_hd__buf_2
XANTENNA__15947__A _13442_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21672__B2 _21666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17046_ _17007_/X _17046_/B VGND VGND VPWR VPWR _17047_/A sky130_fd_sc_hd__or2_4
XFILLER_67_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14258_ _14367_/A _14253_/X _14257_/X VGND VGND VPWR VPWR _14259_/C sky130_fd_sc_hd__or3_4
XANTENNA__19617__A1 _20754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13209_ _13239_/A _13141_/B VGND VGND VPWR VPWR _13210_/C sky130_fd_sc_hd__or2_4
XANTENNA__13467__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21424__B2 _21423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14189_ _14206_/A _14189_/B _14189_/C VGND VGND VPWR VPWR _14190_/C sky130_fd_sc_hd__and3_4
XFILLER_63_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12371__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21975__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13186__B _24081_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18997_ _18995_/Y _18996_/Y _11524_/X VGND VGND VPWR VPWR _18997_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15682__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17948_ _16927_/X _17945_/X _17639_/X _17947_/X VGND VGND VPWR VPWR _17948_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21727__A2 _21726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17879_ _17270_/X _17875_/X _17878_/X VGND VGND VPWR VPWR _17879_/X sky130_fd_sc_hd__o21a_4
XFILLER_22_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14298__A _12459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20935__B1 _20934_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19618_ _24144_/Q _19435_/X HRDATA[18] _19432_/X VGND VGND VPWR VPWR _19618_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11715__A _11715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20890_ _20282_/A _20889_/X VGND VGND VPWR VPWR _20890_/Y sky130_fd_sc_hd__nand2_4
X_19549_ _19449_/A VGND VGND VPWR VPWR _19549_/X sky130_fd_sc_hd__buf_2
XFILLER_81_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18356__A1 _17893_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13930__A _15036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22560_ _22456_/X _22557_/X _15259_/B _22554_/X VGND VGND VPWR VPWR _23170_/D sky130_fd_sc_hd__o22a_4
XFILLER_74_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21511_ _21510_/X _21508_/X _23772_/Q _21503_/X VGND VGND VPWR VPWR _21511_/X sky130_fd_sc_hd__o22a_4
X_22491_ _22422_/X _22486_/X _13336_/B _22490_/X VGND VGND VPWR VPWR _23216_/D sky130_fd_sc_hd__o22a_4
XFILLER_37_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12546__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24230_ _24230_/CLK _19348_/X HRESETn VGND VGND VPWR VPWR _20833_/A sky130_fd_sc_hd__dfrtp_4
X_21442_ _21285_/X _21440_/X _23811_/Q _21437_/X VGND VGND VPWR VPWR _21442_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21859__A _21574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19856__A1 _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24161_ _24165_/CLK _19879_/Y HRESETn VGND VGND VPWR VPWR _16919_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15857__A _13529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20466__A2 _20844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21373_ _21373_/A VGND VGND VPWR VPWR _21373_/X sky130_fd_sc_hd__buf_2
XANTENNA__21663__B2 _21659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23112_ _23816_/CLK _22652_/X VGND VGND VPWR VPWR _13660_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20324_ _20255_/X _20323_/X _24380_/Q _18872_/B VGND VGND VPWR VPWR _20324_/X sky130_fd_sc_hd__o22a_4
X_24092_ _24092_/CLK _24092_/D VGND VGND VPWR VPWR _24092_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15576__B _23691_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14480__B _14480_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23043_ _19901_/X _17891_/B _22899_/X VGND VGND VPWR VPWR _23043_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21415__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22612__B1 _14882_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20255_ _20255_/A VGND VGND VPWR VPWR _20255_/X sky130_fd_sc_hd__buf_2
XANTENNA__12281__A _11596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20186_ _19379_/X _17737_/A _19313_/A _20185_/X VGND VGND VPWR VPWR _20187_/A sky130_fd_sc_hd__o22a_4
XFILLER_103_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15592__A _15592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21179__B1 _12287_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21718__A2 _21712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23945_ _23494_/CLK _23945_/D VGND VGND VPWR VPWR _23945_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19792__B1 _16630_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11890_ _11890_/A VGND VGND VPWR VPWR _12880_/A sky130_fd_sc_hd__buf_2
X_23876_ _23107_/CLK _23876_/D VGND VGND VPWR VPWR _14688_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14001__A _14021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22827_ _22779_/X VGND VGND VPWR VPWR _22827_/X sky130_fd_sc_hd__buf_2
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13560_ _13511_/X _13558_/X _13560_/C VGND VGND VPWR VPWR _13560_/X sky130_fd_sc_hd__and3_4
XFILLER_25_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17312__A _14429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22758_ _22756_/Y _22758_/B _22754_/X VGND VGND VPWR VPWR _24098_/D sky130_fd_sc_hd__and3_4
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12511_ _13623_/A VGND VGND VPWR VPWR _12512_/A sky130_fd_sc_hd__buf_2
XFILLER_38_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21709_ _21702_/A VGND VGND VPWR VPWR _21709_/X sky130_fd_sc_hd__buf_2
XFILLER_16_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24331__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13491_ _13491_/A _13491_/B VGND VGND VPWR VPWR _13491_/X sky130_fd_sc_hd__and2_4
X_22689_ _20574_/A _22686_/X _13193_/B _22683_/X VGND VGND VPWR VPWR _22689_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12456__A _12865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15230_ _15203_/A _15228_/X _15229_/X VGND VGND VPWR VPWR _15230_/X sky130_fd_sc_hd__and3_4
X_12442_ _12850_/A VGND VGND VPWR VPWR _12443_/A sky130_fd_sc_hd__buf_2
X_24428_ _24334_/CLK _18793_/X HRESETn VGND VGND VPWR VPWR _24428_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15581__A1 _11977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21769__A _21740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20673__A _20444_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16870__B _16870_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15161_ _14136_/A _15161_/B _15160_/X VGND VGND VPWR VPWR _15161_/X sky130_fd_sc_hd__or3_4
XFILLER_103_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15767__A _15743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12373_ _12373_/A VGND VGND VPWR VPWR _12926_/A sky130_fd_sc_hd__buf_2
X_24359_ _24330_/CLK _24359_/D HRESETn VGND VGND VPWR VPWR _19068_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__21654__B2 _21652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14671__A _14679_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23505__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_50_0_HCLK clkbuf_5_25_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14112_ _15019_/A VGND VGND VPWR VPWR _14113_/A sky130_fd_sc_hd__buf_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15092_ _15104_/A _15090_/X _15091_/X VGND VGND VPWR VPWR _15092_/X sky130_fd_sc_hd__and3_4
XFILLER_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14390__B _14301_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14043_ _14815_/A _14041_/X _14042_/X VGND VGND VPWR VPWR _14043_/X sky130_fd_sc_hd__and3_4
X_18920_ _15119_/X _18891_/A _24351_/Q _18892_/A VGND VGND VPWR VPWR _24351_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21406__A1 _21221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21406__B2 _21402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12191__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21957__A2 _21952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18851_ _14261_/X _18848_/X _24393_/Q _18849_/X VGND VGND VPWR VPWR _18851_/X sky130_fd_sc_hd__o22a_4
XFILLER_84_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16598__A _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17802_ _17826_/A VGND VGND VPWR VPWR _17802_/X sky130_fd_sc_hd__buf_2
XFILLER_0_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18782_ _18782_/A VGND VGND VPWR VPWR _18782_/X sky130_fd_sc_hd__buf_2
X_15994_ _15994_/A _15992_/X _15994_/C VGND VGND VPWR VPWR _15994_/X sky130_fd_sc_hd__and3_4
XFILLER_114_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17733_ _16965_/C _17106_/X _17729_/X VGND VGND VPWR VPWR _17743_/B sky130_fd_sc_hd__a21bo_4
X_14945_ _11645_/A VGND VGND VPWR VPWR _14970_/A sky130_fd_sc_hd__buf_2
XFILLER_85_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19783__B1 _16652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15007__A _15030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19702__A _19706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17664_ _24130_/Q _17664_/B VGND VGND VPWR VPWR _17685_/A sky130_fd_sc_hd__and2_4
X_14876_ _14906_/A _23520_/Q VGND VGND VPWR VPWR _14877_/C sky130_fd_sc_hd__or2_4
XFILLER_63_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18050__A3 _18044_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19403_ _19302_/X VGND VGND VPWR VPWR _19403_/X sky130_fd_sc_hd__buf_2
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16615_ _16610_/A _23772_/Q VGND VGND VPWR VPWR _16615_/X sky130_fd_sc_hd__or2_4
XFILLER_78_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13827_ _15442_/A _13827_/B _13826_/X VGND VGND VPWR VPWR _13827_/X sky130_fd_sc_hd__or3_4
XFILLER_56_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17595_ _18395_/A _17361_/X _17372_/X _18418_/B VGND VGND VPWR VPWR _17595_/X sky130_fd_sc_hd__or4_4
XANTENNA__14846__A _12599_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18338__B2 _18337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13750__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19334_ _19332_/X _18378_/X _19332_/X _24239_/Q VGND VGND VPWR VPWR _24239_/D sky130_fd_sc_hd__a2bb2o_4
X_13758_ _15495_/A _13756_/X _13757_/X VGND VGND VPWR VPWR _13762_/B sky130_fd_sc_hd__and3_4
X_16546_ _16567_/A _23676_/Q VGND VGND VPWR VPWR _16548_/B sky130_fd_sc_hd__or2_4
X_12709_ _12709_/A _12707_/X _12709_/C VGND VGND VPWR VPWR _12709_/X sky130_fd_sc_hd__and3_4
XFILLER_17_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19265_ _19220_/X VGND VGND VPWR VPWR _19265_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21893__A1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13689_ _14207_/A VGND VGND VPWR VPWR _13690_/A sky130_fd_sc_hd__buf_2
X_16477_ _16159_/X _16401_/B VGND VGND VPWR VPWR _16477_/X sky130_fd_sc_hd__or2_4
XANTENNA__12366__A _11740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21893__B2 _21891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18216_ _18216_/A VGND VGND VPWR VPWR _18216_/X sky130_fd_sc_hd__buf_2
X_15428_ _15442_/A _15424_/X _15428_/C VGND VGND VPWR VPWR _15428_/X sky130_fd_sc_hd__or3_4
XFILLER_34_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19196_ _19111_/A _19197_/A _19195_/Y VGND VGND VPWR VPWR _19196_/X sky130_fd_sc_hd__o21a_4
XFILLER_89_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15359_ _14810_/A _15293_/B VGND VGND VPWR VPWR _15359_/X sky130_fd_sc_hd__or2_4
X_18147_ _18392_/A _18146_/X VGND VGND VPWR VPWR _18147_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15677__A _12743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18053__A _18224_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18078_ _17862_/X _18077_/X _17869_/X VGND VGND VPWR VPWR _18078_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__15396__B _15459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18988__A _19002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13197__A _15707_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17029_ _17040_/A VGND VGND VPWR VPWR _18864_/C sky130_fd_sc_hd__inv_2
XFILLER_119_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20040_ _20018_/X _17699_/X _20024_/X _20039_/X VGND VGND VPWR VPWR _20041_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21948__A2 _21945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13925__A _13925_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20620__A2 HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21991_ _21821_/X _21988_/X _13138_/B _21985_/X VGND VGND VPWR VPWR _21991_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22373__A2 _22368_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23730_ _23314_/CLK _21607_/X VGND VGND VPWR VPWR _23730_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20942_ _20841_/X _20941_/X VGND VGND VPWR VPWR _20942_/X sky130_fd_sc_hd__and2_4
XFILLER_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20384__A1 _20293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _23826_/CLK _21714_/X VGND VGND VPWR VPWR _15798_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _20512_/A VGND VGND VPWR VPWR _20873_/X sky130_fd_sc_hd__buf_2
XFILLER_53_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18228__A _18129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22612_ _22460_/X _22607_/X _14882_/B _22576_/A VGND VGND VPWR VPWR _23136_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13660__A _15429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23592_ _23368_/CLK _23592_/D VGND VGND VPWR VPWR _23592_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22543_ _22536_/A VGND VGND VPWR VPWR _22543_/X sky130_fd_sc_hd__buf_2
XANTENNA__12276__A _12711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23528__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22474_ _22394_/X _22472_/X _16672_/B _22469_/X VGND VGND VPWR VPWR _23228_/D sky130_fd_sc_hd__o22a_4
XANTENNA__20493__A _20493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24213_ _24239_/CLK _19381_/X HRESETn VGND VGND VPWR VPWR _24213_/Q sky130_fd_sc_hd__dfrtp_4
X_21425_ _21256_/X _21419_/X _23823_/Q _21423_/X VGND VGND VPWR VPWR _21425_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18501__A1 _18499_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24144_ _24230_/CLK _24144_/D HRESETn VGND VGND VPWR VPWR _24144_/Q sky130_fd_sc_hd__dfrtp_4
X_21356_ _21221_/X _21355_/X _23869_/Q _21352_/X VGND VGND VPWR VPWR _21356_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18898__A _18898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20307_ _20291_/X _20306_/X VGND VGND VPWR VPWR _20307_/Y sky130_fd_sc_hd__nor2_4
X_24075_ _23688_/CLK _24075_/D VGND VGND VPWR VPWR _24075_/Q sky130_fd_sc_hd__dfxtp_4
X_21287_ _21287_/A VGND VGND VPWR VPWR _21287_/X sky130_fd_sc_hd__buf_2
XFILLER_2_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20940__B _20754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21939__A2 _21938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23026_ _22967_/A VGND VGND VPWR VPWR _23026_/X sky130_fd_sc_hd__buf_2
XFILLER_104_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20238_ _20447_/A VGND VGND VPWR VPWR _20238_/X sky130_fd_sc_hd__buf_2
XANTENNA__22061__B2 _22056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13835__A _15450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20169_ _20134_/Y _20169_/B VGND VGND VPWR VPWR _20169_/X sky130_fd_sc_hd__and2_4
XFILLER_77_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16211__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12991_ _12990_/X VGND VGND VPWR VPWR _12991_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22364__A2 _22361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11942_ _11983_/A VGND VGND VPWR VPWR _11943_/A sky130_fd_sc_hd__buf_2
X_14730_ _14734_/A _14728_/X _14730_/C VGND VGND VPWR VPWR _14731_/C sky130_fd_sc_hd__and3_4
XANTENNA__19522__A _19866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23928_ _24088_/CLK _23928_/D VGND VGND VPWR VPWR _23928_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20668__A _20534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20375__B2 _20374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14661_ _15105_/A _14661_/B VGND VGND VPWR VPWR _14661_/X sky130_fd_sc_hd__or2_4
X_11873_ _11872_/X VGND VGND VPWR VPWR _16147_/A sky130_fd_sc_hd__buf_2
X_23859_ _23859_/CLK _21370_/X VGND VGND VPWR VPWR _23859_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14666__A _14252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18138__A _18266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22116__A2 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13612_ _13800_/A VGND VGND VPWR VPWR _15424_/A sky130_fd_sc_hd__buf_2
X_16400_ _16400_/A _22304_/A VGND VGND VPWR VPWR _16400_/X sky130_fd_sc_hd__or2_4
XFILLER_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13570__A _12754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14592_ _14737_/A _14590_/X _14591_/X VGND VGND VPWR VPWR _14592_/X sky130_fd_sc_hd__and3_4
X_17380_ _17380_/A _17380_/B VGND VGND VPWR VPWR _18418_/B sky130_fd_sc_hd__or2_4
XANTENNA__22883__A _22882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13543_ _13559_/A _13466_/B VGND VGND VPWR VPWR _13543_/X sky130_fd_sc_hd__or2_4
X_16331_ _16322_/A _16256_/B VGND VGND VPWR VPWR _16331_/X sky130_fd_sc_hd__or2_4
X_16262_ _16095_/A _16258_/X _16261_/X VGND VGND VPWR VPWR _16262_/X sky130_fd_sc_hd__or3_4
X_19050_ _19024_/X _19048_/Y _19049_/Y _19027_/X VGND VGND VPWR VPWR _19050_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21499__A _21112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13474_ _11913_/X _13474_/B _13474_/C VGND VGND VPWR VPWR _13475_/C sky130_fd_sc_hd__and3_4
X_15213_ _14210_/A _15213_/B VGND VGND VPWR VPWR _15214_/C sky130_fd_sc_hd__or2_4
X_18001_ _17950_/X _17953_/X _17006_/X _18000_/X VGND VGND VPWR VPWR _18001_/X sky130_fd_sc_hd__o22a_4
X_12425_ _13550_/A _12423_/X _12425_/C VGND VGND VPWR VPWR _12426_/C sky130_fd_sc_hd__and3_4
XFILLER_16_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15497__A _15497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16193_ _16193_/A _23991_/Q VGND VGND VPWR VPWR _16194_/C sky130_fd_sc_hd__or2_4
XFILLER_103_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21627__B2 _21623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12914__A _12914_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15144_ _15144_/A _15144_/B _15143_/X VGND VGND VPWR VPWR _15144_/X sky130_fd_sc_hd__and3_4
X_12356_ _12828_/A _12229_/B VGND VGND VPWR VPWR _12357_/C sky130_fd_sc_hd__or2_4
XFILLER_99_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15075_ _15110_/A _23423_/Q VGND VGND VPWR VPWR _15075_/X sky130_fd_sc_hd__or2_4
X_19952_ _18745_/Y _19950_/X _17998_/X VGND VGND VPWR VPWR _19952_/Y sky130_fd_sc_hd__a21oi_4
X_12287_ _12286_/X _12287_/B VGND VGND VPWR VPWR _12288_/C sky130_fd_sc_hd__or2_4
XFILLER_107_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14026_ _14026_/A VGND VGND VPWR VPWR _14035_/A sky130_fd_sc_hd__buf_2
X_18903_ _17191_/X _18898_/X _24364_/Q _18899_/X VGND VGND VPWR VPWR _24364_/D sky130_fd_sc_hd__o22a_4
XFILLER_64_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19883_ _19447_/X _19882_/X _17079_/A _19493_/X VGND VGND VPWR VPWR _19883_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__19416__B _19416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15944__B _16019_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18834_ _18834_/A VGND VGND VPWR VPWR _18834_/X sky130_fd_sc_hd__buf_2
XANTENNA__13745__A _12937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20602__A2 _20601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16121__A _16121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_57_0_HCLK clkbuf_6_28_0_HCLK/X VGND VGND VPWR VPWR _23564_/CLK sky130_fd_sc_hd__clkbuf_1
X_18765_ _18781_/A VGND VGND VPWR VPWR _18765_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15977_ _15984_/A _23608_/Q VGND VGND VPWR VPWR _15977_/X sky130_fd_sc_hd__or2_4
XFILLER_76_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22355__A2 _22354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17716_ _17716_/A _17712_/X VGND VGND VPWR VPWR _17716_/X sky130_fd_sc_hd__or2_4
X_14928_ _12582_/A _14864_/B VGND VGND VPWR VPWR _14929_/C sky130_fd_sc_hd__or2_4
XFILLER_97_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18696_ _18499_/X _17325_/X _18500_/X VGND VGND VPWR VPWR _18696_/X sky130_fd_sc_hd__a21o_4
XANTENNA__17231__A1 _17165_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17647_ _17647_/A VGND VGND VPWR VPWR _17647_/X sky130_fd_sc_hd__buf_2
X_14859_ _13983_/A _14859_/B VGND VGND VPWR VPWR _14859_/X sky130_fd_sc_hd__or2_4
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18048__A _18048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19508__B1 HRDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13480__A _13448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17578_ _16814_/B _17278_/B _17282_/Y _17577_/X VGND VGND VPWR VPWR _17578_/X sky130_fd_sc_hd__o22a_4
XFILLER_95_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12808__B _23892_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19317_ _19317_/A VGND VGND VPWR VPWR _19328_/A sky130_fd_sc_hd__buf_2
X_16529_ _16541_/A _16527_/X _16529_/C VGND VGND VPWR VPWR _16533_/B sky130_fd_sc_hd__and3_4
XFILLER_32_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20669__A2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12096__A _12096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19248_ _24280_/Q _19249_/A _19247_/Y VGND VGND VPWR VPWR _24280_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21618__B2 _21616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19179_ _19120_/B VGND VGND VPWR VPWR _19179_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21210_ _21002_/X _21183_/A _15088_/B _21165_/X VGND VGND VPWR VPWR _23935_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22017__B _22017_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21094__A2 _21089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22190_ _22169_/A VGND VGND VPWR VPWR _22190_/X sky130_fd_sc_hd__buf_2
XANTENNA__22291__B2 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21141_ _20637_/X _21140_/X _15667_/B _21137_/X VGND VGND VPWR VPWR _23982_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22043__A1 _21823_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21072_ _21072_/A VGND VGND VPWR VPWR _21072_/X sky130_fd_sc_hd__buf_2
XFILLER_67_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22043__B2 _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18798__A1 _14261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22594__A2 _22593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20023_ _20023_/A VGND VGND VPWR VPWR _20023_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17127__A _17126_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13655__A _13794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22968__A _22968_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17470__A1 _17466_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21872__A _21901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17470__B2 _17469_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15870__A _13551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21974_ _21988_/A VGND VGND VPWR VPWR _21974_/X sky130_fd_sc_hd__buf_2
XANTENNA__20488__A _20488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23713_ _23819_/CLK _21630_/X VGND VGND VPWR VPWR _23713_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17222__A1 _18728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20925_ _24386_/Q _20405_/A _24418_/Q _20449_/A VGND VGND VPWR VPWR _20925_/X sky130_fd_sc_hd__o22a_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14486__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11903__A _11903_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13390__A _12822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23644_ _23867_/CLK _23644_/D VGND VGND VPWR VPWR _23644_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20856_ _20855_/Y _20708_/B VGND VGND VPWR VPWR _20856_/X sky130_fd_sc_hd__or2_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21306__B1 _23901_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12718__B _23892_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23575_ _23699_/CLK _23575_/D VGND VGND VPWR VPWR _23575_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20787_ _20622_/X _20786_/X _19213_/A _20736_/X VGND VGND VPWR VPWR _20787_/X sky130_fd_sc_hd__o22a_4
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18722__B2 _22824_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22526_ _22518_/X VGND VGND VPWR VPWR _22526_/X sky130_fd_sc_hd__buf_2
XANTENNA__23059__B1 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22208__A _22222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21112__A _21112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22457_ _22456_/X _22452_/X _15252_/B _22447_/X VGND VGND VPWR VPWR _23234_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12734__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _13635_/A VGND VGND VPWR VPWR _12211_/A sky130_fd_sc_hd__buf_2
X_21408_ _21227_/X _21405_/X _23835_/Q _21402_/X VGND VGND VPWR VPWR _23835_/D sky130_fd_sc_hd__o22a_4
XFILLER_87_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22282__A1 _22117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21085__A2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13190_ _15785_/A _13190_/B VGND VGND VPWR VPWR _13190_/X sky130_fd_sc_hd__or2_4
XANTENNA__13549__B _23823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22388_ _20276_/A VGND VGND VPWR VPWR _22388_/X sky130_fd_sc_hd__buf_2
XFILLER_109_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22282__B2 _22276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12141_ _11820_/A _12139_/X _12141_/C VGND VGND VPWR VPWR _12141_/X sky130_fd_sc_hd__and3_4
X_24127_ _23522_/CLK _20023_/Y HRESETn VGND VGND VPWR VPWR _18234_/A sky130_fd_sc_hd__dfrtp_4
X_21339_ _21280_/X _21333_/X _14532_/B _21337_/X VGND VGND VPWR VPWR _23877_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19517__A _19517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24186__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18421__A _18421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18238__B1 _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12072_ _12068_/X _12069_/X _12072_/C VGND VGND VPWR VPWR _12073_/C sky130_fd_sc_hd__and3_4
X_24058_ _23472_/CLK _21021_/X VGND VGND VPWR VPWR _16417_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22034__B2 _22028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15900_ _13522_/A _15900_/B _15900_/C VGND VGND VPWR VPWR _15904_/B sky130_fd_sc_hd__and3_4
X_23009_ _22980_/A VGND VGND VPWR VPWR _23017_/B sky130_fd_sc_hd__buf_2
XANTENNA__13565__A _13551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22585__A2 _22579_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16880_ _16525_/X _16816_/X _16525_/X _16816_/X VGND VGND VPWR VPWR _16887_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15831_ _12872_/A _15831_/B VGND VGND VPWR VPWR _15831_/X sky130_fd_sc_hd__or2_4
XANTENNA__15780__A _15713_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19738__B1 _12101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18550_ _17746_/X _17747_/B _17713_/X VGND VGND VPWR VPWR _18550_/X sky130_fd_sc_hd__o21a_4
X_12974_ _12974_/A _12974_/B VGND VGND VPWR VPWR _12975_/C sky130_fd_sc_hd__or2_4
X_15762_ _15750_/A _15762_/B VGND VGND VPWR VPWR _15762_/X sky130_fd_sc_hd__or2_4
XFILLER_59_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20398__A _20512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21545__B1 _15722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17501_ _17175_/Y _17498_/X VGND VGND VPWR VPWR _17501_/X sky130_fd_sc_hd__and2_4
XANTENNA__17213__A1 _12676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14713_ _14341_/A _14627_/B VGND VGND VPWR VPWR _14715_/B sky130_fd_sc_hd__or2_4
X_11925_ _12529_/A VGND VGND VPWR VPWR _11925_/Y sky130_fd_sc_hd__inv_2
X_18481_ _18349_/A _18349_/B VGND VGND VPWR VPWR _18481_/Y sky130_fd_sc_hd__nand2_4
X_15693_ _15693_/A _15758_/B VGND VGND VPWR VPWR _15694_/C sky130_fd_sc_hd__or2_4
XFILLER_75_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17432_ _17192_/Y _17432_/B VGND VGND VPWR VPWR _17432_/X sky130_fd_sc_hd__or2_4
X_11856_ _13986_/A VGND VGND VPWR VPWR _13972_/A sky130_fd_sc_hd__buf_2
X_14644_ _14644_/A VGND VGND VPWR VPWR _15105_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14575_ _14997_/A VGND VGND VPWR VPWR _14575_/X sky130_fd_sc_hd__buf_2
X_17363_ _17363_/A VGND VGND VPWR VPWR _17506_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15004__B _15079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11787_ _11819_/A _21110_/A VGND VGND VPWR VPWR _11787_/X sky130_fd_sc_hd__or2_4
XFILLER_109_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19102_ _24319_/Q _18999_/A _18935_/X VGND VGND VPWR VPWR _19102_/X sky130_fd_sc_hd__a21o_4
XANTENNA__20845__B _20650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16314_ _16185_/A _16248_/B VGND VGND VPWR VPWR _16316_/B sky130_fd_sc_hd__or2_4
X_13526_ _13562_/A _13457_/B VGND VGND VPWR VPWR _13527_/C sky130_fd_sc_hd__or2_4
X_17294_ _14565_/Y _17294_/B VGND VGND VPWR VPWR _17605_/A sky130_fd_sc_hd__or2_4
XANTENNA__15939__B _23352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19033_ _19031_/Y _19032_/Y _11519_/B VGND VGND VPWR VPWR _19033_/X sky130_fd_sc_hd__o21a_4
X_13457_ _12477_/X _13457_/B VGND VGND VPWR VPWR _13458_/C sky130_fd_sc_hd__or2_4
X_16245_ _16150_/A _16245_/B VGND VGND VPWR VPWR _16245_/X sky130_fd_sc_hd__or2_4
XANTENNA__12644__A _12963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12408_ _11671_/A VGND VGND VPWR VPWR _13572_/A sky130_fd_sc_hd__buf_2
XANTENNA__15020__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22273__A1 _22100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13388_ _13388_/A _13388_/B _13387_/X VGND VGND VPWR VPWR _13389_/C sky130_fd_sc_hd__and3_4
X_16176_ _13378_/X VGND VGND VPWR VPWR _16193_/A sky130_fd_sc_hd__buf_2
XANTENNA__22273__B2 _22269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_20_0_HCLK clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12339_ _11645_/A VGND VGND VPWR VPWR _12340_/A sky130_fd_sc_hd__buf_2
X_15127_ _12196_/A _15125_/X _15127_/C VGND VGND VPWR VPWR _15127_/X sky130_fd_sc_hd__and3_4
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15058_ _11723_/A _15058_/B _15058_/C VGND VGND VPWR VPWR _15058_/X sky130_fd_sc_hd__and3_4
X_19935_ _22888_/A _19927_/X VGND VGND VPWR VPWR _19936_/A sky130_fd_sc_hd__or2_4
XFILLER_64_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15674__B _15674_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14009_ _14009_/A VGND VGND VPWR VPWR _14815_/A sky130_fd_sc_hd__buf_2
XANTENNA__13475__A _11861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19866_ _19454_/A _19866_/B VGND VGND VPWR VPWR _19866_/X sky130_fd_sc_hd__or2_4
XFILLER_64_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22788__A _17298_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18817_ _18841_/A VGND VGND VPWR VPWR _18834_/A sky130_fd_sc_hd__buf_2
XFILLER_56_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19797_ _19667_/A _19796_/X VGND VGND VPWR VPWR _19797_/Y sky130_fd_sc_hd__nand2_4
XFILLER_95_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14266__A1 _14174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15690__A _12722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18748_ _17057_/A _19941_/B _17057_/A _19941_/B VGND VGND VPWR VPWR _18748_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16007__A2 _11619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18679_ _18487_/X _18671_/X _18672_/Y _18674_/X _18678_/Y VGND VGND VPWR VPWR _18679_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_97_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12819__A _12803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20710_ _20654_/X _20705_/Y _20708_/X _19044_/Y _20709_/X VGND VGND VPWR VPWR _20710_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12029__B1 _11598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21690_ _21690_/A VGND VGND VPWR VPWR _21705_/A sky130_fd_sc_hd__buf_2
XFILLER_63_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20641_ _11579_/X VGND VGND VPWR VPWR _20641_/X sky130_fd_sc_hd__buf_2
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21839__B2 _21836_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23360_ _24032_/CLK _23360_/D VGND VGND VPWR VPWR _14898_/B sky130_fd_sc_hd__dfxtp_4
X_20572_ _24209_/Q _20512_/X _20571_/X VGND VGND VPWR VPWR _20573_/A sky130_fd_sc_hd__o21a_4
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22028__A _22020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22311_ _22311_/A VGND VGND VPWR VPWR _23315_/D sky130_fd_sc_hd__buf_2
X_23291_ _23293_/CLK _23291_/D VGND VGND VPWR VPWR _16759_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12554__A _13046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22242_ _22134_/X _22236_/X _14472_/B _22240_/X VGND VGND VPWR VPWR _23365_/D sky130_fd_sc_hd__o22a_4
XFILLER_30_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11555__A2 IRQ[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15865__A _13511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22173_ _22100_/X _22172_/X _23411_/Q _22169_/X VGND VGND VPWR VPWR _22173_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20490__B _20490_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21124_ _20373_/X _21119_/X _16398_/B _21123_/X VGND VGND VPWR VPWR _21124_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15584__B _23499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13385__A _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21055_ _20958_/X _21051_/X _15159_/B _21012_/X VGND VGND VPWR VPWR _21055_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21775__B1 _14480_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20006_ _18227_/X _19985_/X _20005_/Y _19996_/X VGND VGND VPWR VPWR _20006_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17443__A1 _17439_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18640__B1 _17998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17443__B2 _17667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_40_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR _23816_/CLK sky130_fd_sc_hd__clkbuf_1
X_21957_ _21847_/X _21952_/X _14289_/B _21956_/X VGND VGND VPWR VPWR _23526_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12729__A _12743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A VGND VGND VPWR VPWR _12373_/A sky130_fd_sc_hd__buf_2
XFILLER_76_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20715_/A _20908_/B VGND VGND VPWR VPWR _20908_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15105__A _15105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12690_ _12221_/X _12773_/B VGND VGND VPWR VPWR _12692_/B sky130_fd_sc_hd__or2_4
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _21816_/X _21887_/X _12943_/B _21884_/X VGND VGND VPWR VPWR _21888_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _14177_/A VGND VGND VPWR VPWR _11642_/A sky130_fd_sc_hd__buf_2
X_23627_ _23688_/CLK _23627_/D VGND VGND VPWR VPWR _15570_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_42_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _20488_/A VGND VGND VPWR VPWR _20839_/X sky130_fd_sc_hd__buf_2
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _15598_/A _14278_/B VGND VGND VPWR VPWR _14360_/X sky130_fd_sc_hd__or2_4
XFILLER_11_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _24444_/Q IRQ[29] _20166_/A VGND VGND VPWR VPWR _11572_/X sky130_fd_sc_hd__a21o_4
X_23558_ _23845_/CLK _23558_/D VGND VGND VPWR VPWR _14293_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _15696_/A _13311_/B VGND VGND VPWR VPWR _13311_/X sky130_fd_sc_hd__or2_4
XFILLER_89_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22509_ _22454_/X _22507_/X _14772_/B _22504_/X VGND VGND VPWR VPWR _22509_/X sky130_fd_sc_hd__o22a_4
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14291_ _11859_/A _14285_/X _14290_/X VGND VGND VPWR VPWR _14291_/X sky130_fd_sc_hd__or3_4
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23489_ _23391_/CLK _22013_/X VGND VGND VPWR VPWR _15126_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_11_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12464__A _12464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13242_ _13242_/A _24049_/Q VGND VGND VPWR VPWR _13243_/C sky130_fd_sc_hd__or2_4
X_16030_ _16019_/A _23928_/Q VGND VGND VPWR VPWR _16032_/B sky130_fd_sc_hd__or2_4
XFILLER_109_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23246__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20681__A _20253_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11546__A2 IRQ[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13173_ _12255_/X _13171_/X _13173_/C VGND VGND VPWR VPWR _13173_/X sky130_fd_sc_hd__and3_4
XANTENNA__15775__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12124_ _16072_/A VGND VGND VPWR VPWR _12168_/A sky130_fd_sc_hd__buf_2
XANTENNA__22007__B2 _22006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17981_ _17801_/X _17842_/X _17807_/X _17838_/X VGND VGND VPWR VPWR _17981_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_46_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12911__B _12983_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19720_ _19873_/B _19720_/B VGND VGND VPWR VPWR _19740_/B sky130_fd_sc_hd__or2_4
XANTENNA__13295__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22558__A2 _22557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12055_ _11875_/X VGND VGND VPWR VPWR _12088_/A sky130_fd_sc_hd__buf_2
X_16932_ _16931_/X VGND VGND VPWR VPWR _16933_/A sky130_fd_sc_hd__inv_2
X_19651_ _19554_/X _19644_/Y _19648_/Y _19445_/X _19650_/Y VGND VGND VPWR VPWR _19651_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18631__B1 _18424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16863_ _15388_/X VGND VGND VPWR VPWR _16863_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22401__A _20393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18602_ _24453_/Q VGND VGND VPWR VPWR _18602_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15814_ _12443_/A _23885_/Q VGND VGND VPWR VPWR _15814_/X sky130_fd_sc_hd__or2_4
XFILLER_20_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19582_ _19582_/A VGND VGND VPWR VPWR _19582_/Y sky130_fd_sc_hd__inv_2
X_16794_ _16598_/X _16790_/X _16793_/X VGND VGND VPWR VPWR _16795_/C sky130_fd_sc_hd__or3_4
XFILLER_59_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14838__B _14780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18533_ _18533_/A _18174_/D VGND VGND VPWR VPWR _18533_/Y sky130_fd_sc_hd__nand2_4
XFILLER_59_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15745_ _13102_/A _15735_/X _15744_/X VGND VGND VPWR VPWR _15745_/X sky130_fd_sc_hd__and3_4
X_12957_ _12957_/A _12957_/B _12957_/C VGND VGND VPWR VPWR _12957_/X sky130_fd_sc_hd__or3_4
XFILLER_73_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12639__A _12591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15015__A _15015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11908_ _14998_/A VGND VGND VPWR VPWR _11909_/A sky130_fd_sc_hd__buf_2
X_18464_ _18418_/A _18395_/A VGND VGND VPWR VPWR _18464_/X sky130_fd_sc_hd__or2_4
XFILLER_33_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19710__A _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15676_ _12742_/A _15732_/B VGND VGND VPWR VPWR _15678_/B sky130_fd_sc_hd__or2_4
X_12888_ _12518_/A _12945_/B VGND VGND VPWR VPWR _12888_/X sky130_fd_sc_hd__or2_4
X_17415_ _14263_/X _17414_/X VGND VGND VPWR VPWR _17416_/A sky130_fd_sc_hd__or2_4
XFILLER_21_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14627_ _13606_/A _14627_/B VGND VGND VPWR VPWR _14629_/B sky130_fd_sc_hd__or2_4
X_11839_ _11838_/Y VGND VGND VPWR VPWR _11839_/X sky130_fd_sc_hd__buf_2
X_18395_ _18395_/A _17361_/X _18395_/C VGND VGND VPWR VPWR _18395_/X sky130_fd_sc_hd__or3_4
X_17346_ _17363_/A _17345_/X VGND VGND VPWR VPWR _17346_/X sky130_fd_sc_hd__or2_4
XFILLER_53_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14558_ _13697_/X _14480_/B VGND VGND VPWR VPWR _14559_/C sky130_fd_sc_hd__or2_4
XFILLER_14_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22494__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13509_ _15884_/A _13435_/B VGND VGND VPWR VPWR _13510_/C sky130_fd_sc_hd__or2_4
X_17277_ _16812_/X VGND VGND VPWR VPWR _17277_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12374__A _12926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14489_ _15435_/A _14485_/X _14489_/C VGND VGND VPWR VPWR _14490_/B sky130_fd_sc_hd__or3_4
X_19016_ _19002_/A VGND VGND VPWR VPWR _19016_/X sky130_fd_sc_hd__buf_2
X_16228_ _16206_/A _16226_/X _16228_/C VGND VGND VPWR VPWR _16228_/X sky130_fd_sc_hd__and3_4
XANTENNA__21687__A _21702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21049__A2 _21044_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22246__B2 _22240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12093__B _12162_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24171__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11537__A2 IRQ[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15685__A _15685_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16159_ _13397_/X VGND VGND VPWR VPWR _16159_/X sky130_fd_sc_hd__buf_2
XANTENNA__17122__B1 _21007_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22549__A2 _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11718__A _11717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19918_ _19916_/X _24147_/Q _19917_/X _20490_/B VGND VGND VPWR VPWR _24147_/D sky130_fd_sc_hd__o22a_4
XFILLER_111_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19849_ _19678_/A _19845_/X _19848_/Y _21007_/A _19531_/A VGND VGND VPWR VPWR _19849_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18622__B1 _18063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13933__A _14782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_27_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_54_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22860_ _16008_/Y _22814_/X _22853_/X _22859_/X VGND VGND VPWR VPWR _22861_/B sky130_fd_sc_hd__o22a_4
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21509__B1 _23773_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20980__A1 _24192_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21811_ _20487_/A VGND VGND VPWR VPWR _21811_/X sky130_fd_sc_hd__buf_2
XANTENNA__19717__A3 _19716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22791_ _22777_/X VGND VGND VPWR VPWR _22862_/A sky130_fd_sc_hd__buf_2
XANTENNA__12549__A _12914_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21742_ _21506_/X _21741_/X _23645_/Q _21738_/X VGND VGND VPWR VPWR _21742_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24461_ _24126_/CLK _18434_/X HRESETn VGND VGND VPWR VPWR _24461_/Q sky130_fd_sc_hd__dfrtp_4
X_21673_ _21659_/A VGND VGND VPWR VPWR _21673_/X sky130_fd_sc_hd__buf_2
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18236__A _17672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23412_ _23635_/CLK _23412_/D VGND VGND VPWR VPWR _12819_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20624_ _24398_/Q _20623_/X _24430_/Q _20449_/X VGND VGND VPWR VPWR _20624_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22485__A1 _22413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21288__A2 _21283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24392_ _24365_/CLK _18852_/X HRESETn VGND VGND VPWR VPWR _24392_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22981__A _18334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22485__B2 _22483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23343_ _23827_/CLK _23343_/D VGND VGND VPWR VPWR _13502_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20555_ _20422_/X _20939_/B _20286_/A VGND VGND VPWR VPWR _20555_/X sky130_fd_sc_hd__a21o_4
XANTENNA__24460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12284__A _12496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23274_ _24011_/CLK _23274_/D VGND VGND VPWR VPWR _13939_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22237__B2 _22233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13099__B _23538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20486_ _20486_/A VGND VGND VPWR VPWR _20487_/A sky130_fd_sc_hd__buf_2
X_22225_ _22105_/X _22222_/X _13181_/B _22219_/X VGND VGND VPWR VPWR _23377_/D sky130_fd_sc_hd__o22a_4
XFILLER_101_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21996__B1 _15715_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22156_ _22149_/Y _22155_/X _22073_/X _22155_/X VGND VGND VPWR VPWR _22156_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_109_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR _23920_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21107_ _20958_/X _21103_/X _15196_/B _21072_/A VGND VGND VPWR VPWR _24001_/D sky130_fd_sc_hd__o22a_4
XFILLER_47_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22087_ _22086_/X _22077_/X _16267_/B _22084_/X VGND VGND VPWR VPWR _23449_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19405__A2_N _18613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14004__A _14845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21038_ _20637_/X _21037_/X _15686_/B _21034_/X VGND VGND VPWR VPWR _24046_/D sky130_fd_sc_hd__o22a_4
XFILLER_75_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14939__A _11645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13860_ _14002_/A VGND VGND VPWR VPWR _14810_/A sky130_fd_sc_hd__buf_2
XFILLER_47_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12811_ _12799_/A _23604_/Q VGND VGND VPWR VPWR _12811_/X sky130_fd_sc_hd__or2_4
XFILLER_16_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13791_ _15429_/A _13791_/B VGND VGND VPWR VPWR _13793_/B sky130_fd_sc_hd__or2_4
X_22989_ _22989_/A _22989_/B _22988_/X VGND VGND VPWR VPWR _22989_/X sky130_fd_sc_hd__and3_4
XANTENNA__12459__A _12459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18916__A1 _14851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22712__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15530_ _12260_/X _15530_/B VGND VGND VPWR VPWR _15530_/X sky130_fd_sc_hd__or2_4
X_12742_ _12742_/A _12823_/B VGND VGND VPWR VPWR _12742_/X sky130_fd_sc_hd__or2_4
XFILLER_70_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12178__B _23645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20676__A HRDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23052__A _17636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12673_ _12989_/A _12673_/B _12673_/C VGND VGND VPWR VPWR _12673_/X sky130_fd_sc_hd__and3_4
X_15461_ _13738_/A _15456_/X _15460_/X VGND VGND VPWR VPWR _15461_/X sky130_fd_sc_hd__or3_4
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17863_/A _17169_/X _17845_/A _17199_/X VGND VGND VPWR VPWR _17200_/X sky130_fd_sc_hd__o22a_4
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _24383_/Q _11576_/X NMI _20076_/A VGND VGND VPWR VPWR _11624_/X sky130_fd_sc_hd__a211o_4
X_14412_ _15611_/A _14408_/X _14412_/C VGND VGND VPWR VPWR _14421_/B sky130_fd_sc_hd__or3_4
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18180_ _18180_/A _18180_/B _18180_/C _18180_/D VGND VGND VPWR VPWR _18180_/X sky130_fd_sc_hd__or4_4
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21279__A2 _21271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _15392_/A _15454_/B VGND VGND VPWR VPWR _15394_/B sky130_fd_sc_hd__or2_4
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22891__A _23015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14393__B _14304_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ _17173_/A VGND VGND VPWR VPWR _17131_/X sky130_fd_sc_hd__buf_2
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19341__B2 _24235_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11555_ _24424_/Q IRQ[9] _11554_/X VGND VGND VPWR VPWR _11558_/A sky130_fd_sc_hd__a21o_4
X_14343_ _15584_/A _14269_/B VGND VGND VPWR VPWR _14344_/C sky130_fd_sc_hd__or2_4
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14274_ _15412_/A _14270_/X _14273_/X VGND VGND VPWR VPWR _14274_/X sky130_fd_sc_hd__or3_4
X_17062_ _17062_/A _17058_/X _17061_/X VGND VGND VPWR VPWR _17063_/A sky130_fd_sc_hd__and3_4
XANTENNA__24130__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22228__B2 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13225_ _13257_/A _13166_/B VGND VGND VPWR VPWR _13226_/C sky130_fd_sc_hd__or2_4
X_16013_ _16023_/A VGND VGND VPWR VPWR _16019_/A sky130_fd_sc_hd__buf_2
XANTENNA__12922__A _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13156_ _15706_/A VGND VGND VPWR VPWR _15696_/A sky130_fd_sc_hd__buf_2
XFILLER_88_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12107_ _11971_/A _23805_/Q VGND VGND VPWR VPWR _12108_/C sky130_fd_sc_hd__or2_4
XFILLER_112_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13087_ _13087_/A VGND VGND VPWR VPWR _13109_/A sky130_fd_sc_hd__buf_2
X_17964_ _17868_/A VGND VGND VPWR VPWR _17964_/X sky130_fd_sc_hd__buf_2
X_19703_ _19703_/A _19690_/X VGND VGND VPWR VPWR _19703_/X sky130_fd_sc_hd__or2_4
X_12038_ _11875_/X VGND VGND VPWR VPWR _16718_/A sky130_fd_sc_hd__buf_2
X_16915_ _16907_/X _16915_/B _16914_/X VGND VGND VPWR VPWR _16917_/B sky130_fd_sc_hd__and3_4
XANTENNA__21203__A2 _21197_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15952__B _15952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17895_ _17951_/A _17894_/X _18342_/A VGND VGND VPWR VPWR _17895_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_113_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22131__A _22446_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14849__A _14040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19634_ _19499_/A _19633_/X VGND VGND VPWR VPWR _19634_/X sky130_fd_sc_hd__and2_4
XANTENNA__13753__A _12638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16846_ _15928_/X _16239_/B _15928_/X _16239_/B VGND VGND VPWR VPWR _16851_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21970__A _21985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19565_ _19471_/A _19559_/A _19621_/A VGND VGND VPWR VPWR _19729_/C sky130_fd_sc_hd__or3_4
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16777_ _16747_/X _16775_/X _16777_/C VGND VGND VPWR VPWR _16777_/X sky130_fd_sc_hd__and3_4
X_13989_ _11839_/X _11615_/X _13958_/X _11592_/X _13988_/X VGND VGND VPWR VPWR _13989_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_59_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18907__A1 _17171_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22164__B1 _16283_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22703__A2 _22700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18516_ _16957_/A _18515_/Y _16972_/B VGND VGND VPWR VPWR _22939_/B sky130_fd_sc_hd__o21a_4
X_15728_ _13133_/A _15720_/X _15728_/C VGND VGND VPWR VPWR _15746_/B sky130_fd_sc_hd__and3_4
XFILLER_34_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19496_ _19545_/A VGND VGND VPWR VPWR _19496_/X sky130_fd_sc_hd__buf_2
XANTENNA__21911__B1 _15274_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18447_ _17794_/A _18304_/B _17933_/X _18446_/X VGND VGND VPWR VPWR _18447_/X sky130_fd_sc_hd__a211o_4
X_15659_ _12284_/X _15659_/B VGND VGND VPWR VPWR _15661_/B sky130_fd_sc_hd__or2_4
XANTENNA__24289__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18056__A _18129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14584__A _14149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18378_ _18285_/C _17759_/X _18285_/C _17759_/X VGND VGND VPWR VPWR _18378_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15399__B _15462_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17329_ _15121_/X _17220_/A VGND VGND VPWR VPWR _17329_/X sky130_fd_sc_hd__or2_4
XANTENNA__19883__A2 _19882_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20340_ _20280_/X _20339_/X _24092_/Q _20203_/X VGND VGND VPWR VPWR _24092_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13928__A _14778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20271_ _19953_/X _20238_/X _20240_/X _20270_/X VGND VGND VPWR VPWR _20272_/A sky130_fd_sc_hd__a211o_4
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12832__A _12802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16304__A _16185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22010_ _21852_/X _22009_/X _14646_/B _22006_/X VGND VGND VPWR VPWR _23492_/D sky130_fd_sc_hd__o22a_4
XFILLER_66_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21442__A2 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12551__B _12658_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23961_ _23514_/CLK _21175_/X VGND VGND VPWR VPWR _16273_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14759__A _12883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13663__A _15431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22912_ _17726_/X _18642_/A _17724_/X VGND VGND VPWR VPWR _22912_/X sky130_fd_sc_hd__o21a_4
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23892_ _23315_/CLK _21318_/X VGND VGND VPWR VPWR _23892_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_83_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21880__A _21887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22843_ _22843_/A VGND VGND VPWR VPWR HWDATA[20] sky130_fd_sc_hd__inv_2
XFILLER_83_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12279__A _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19350__A _19336_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22774_ _22773_/A _22773_/B _24095_/D _22773_/Y VGND VGND VPWR VPWR _22774_/X sky130_fd_sc_hd__a211o_4
XANTENNA__11614__C _12860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21725_ _21565_/X _21719_/X _14523_/B _21723_/X VGND VGND VPWR VPWR _21725_/X sky130_fd_sc_hd__o22a_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11911__A _11911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21656_ _21531_/X _21655_/X _12976_/B _21652_/X VGND VGND VPWR VPWR _23699_/D sky130_fd_sc_hd__o22a_4
X_24444_ _24277_/CLK _18771_/X HRESETn VGND VGND VPWR VPWR _24444_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23904__CLK _23840_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20607_ _24239_/Q _20421_/X _20606_/X VGND VGND VPWR VPWR _20607_/X sky130_fd_sc_hd__o21a_4
XFILLER_71_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24375_ _24277_/CLK _18888_/X HRESETn VGND VGND VPWR VPWR _18975_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__15102__B _23071_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21587_ _21602_/A VGND VGND VPWR VPWR _21595_/A sky130_fd_sc_hd__buf_2
XANTENNA__19874__A2 _19706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23326_ _23326_/CLK _23326_/D VGND VGND VPWR VPWR _11790_/B sky130_fd_sc_hd__dfxtp_4
X_20538_ _20511_/X _20537_/X _12909_/B _20488_/X VGND VGND VPWR VPWR _20538_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21681__A2 _21676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23257_ _23130_/CLK _23257_/D VGND VGND VPWR VPWR _16240_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13838__A _13690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20469_ _20469_/A _20519_/B VGND VGND VPWR VPWR _20469_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12742__A _12742_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16214__A _16198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13010_ _12917_/A _13010_/B _13010_/C VGND VGND VPWR VPWR _13011_/C sky130_fd_sc_hd__and3_4
XFILLER_84_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22208_ _22222_/A VGND VGND VPWR VPWR _22208_/X sky130_fd_sc_hd__buf_2
XANTENNA__17637__B2 _17636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23188_ _23987_/CLK _23188_/D VGND VGND VPWR VPWR _12773_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_106_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22139_ _20915_/A VGND VGND VPWR VPWR _22139_/X sky130_fd_sc_hd__buf_2
XFILLER_79_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23047__A _17880_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14961_ _14658_/A _14961_/B _14960_/X VGND VGND VPWR VPWR _14969_/B sky130_fd_sc_hd__or3_4
XANTENNA__15772__B _15699_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24354__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14669__A _15115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16700_ _12086_/A _16775_/B VGND VGND VPWR VPWR _16702_/B sky130_fd_sc_hd__or2_4
XANTENNA__13573__A _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13912_ _13909_/A _13824_/B VGND VGND VPWR VPWR _13914_/B sky130_fd_sc_hd__or2_4
X_17680_ _17680_/A _17479_/X VGND VGND VPWR VPWR _17680_/X sky130_fd_sc_hd__or2_4
X_14892_ _14867_/X _14892_/B VGND VGND VPWR VPWR _14892_/X sky130_fd_sc_hd__or2_4
XFILLER_74_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22886__A _22985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16631_ _16630_/X _16631_/B VGND VGND VPWR VPWR _16634_/B sky130_fd_sc_hd__or2_4
Xclkbuf_6_10_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_10_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13843_ _14218_/A VGND VGND VPWR VPWR _13844_/A sky130_fd_sc_hd__buf_2
XFILLER_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12189__A _11842_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22146__B1 _14883_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19350_ _19336_/A VGND VGND VPWR VPWR _19350_/X sky130_fd_sc_hd__buf_2
X_16562_ _11982_/X _16562_/B VGND VGND VPWR VPWR _16562_/X sky130_fd_sc_hd__and2_4
X_13774_ _13685_/Y _13772_/X VGND VGND VPWR VPWR _13774_/X sky130_fd_sc_hd__or2_4
X_18301_ _17862_/A _18300_/X _18183_/X _17867_/X VGND VGND VPWR VPWR _18301_/X sky130_fd_sc_hd__o22a_4
X_15513_ _13087_/A _15511_/X _15513_/C VGND VGND VPWR VPWR _15514_/C sky130_fd_sc_hd__and3_4
XFILLER_95_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12725_ _12725_/A _23124_/Q VGND VGND VPWR VPWR _12727_/B sky130_fd_sc_hd__or2_4
X_19281_ _19213_/B VGND VGND VPWR VPWR _19281_/Y sky130_fd_sc_hd__inv_2
X_16493_ _16473_/X _16424_/B VGND VGND VPWR VPWR _16493_/X sky130_fd_sc_hd__or2_4
XANTENNA__12917__A _12917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18232_ _17889_/A _16999_/C _18231_/Y VGND VGND VPWR VPWR _18233_/B sky130_fd_sc_hd__and3_4
XANTENNA__11821__A _11821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15444_ _13635_/A _23788_/Q VGND VGND VPWR VPWR _15445_/C sky130_fd_sc_hd__or2_4
XFILLER_31_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24311__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12656_ _13118_/A _12656_/B _12655_/X VGND VGND VPWR VPWR _12656_/X sky130_fd_sc_hd__and3_4
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ _15015_/A VGND VGND VPWR VPWR _11608_/A sky130_fd_sc_hd__buf_2
X_18163_ _17950_/X _18133_/X _18022_/X _18162_/X VGND VGND VPWR VPWR _18163_/X sky130_fd_sc_hd__o22a_4
XANTENNA__11540__B IRQ[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12587_ _12970_/A _12580_/X _12587_/C VGND VGND VPWR VPWR _12587_/X sky130_fd_sc_hd__and3_4
X_15375_ _12598_/A _15373_/X _15375_/C VGND VGND VPWR VPWR _15376_/C sky130_fd_sc_hd__and3_4
XFILLER_8_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21121__B2 _21116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17114_ _17114_/A VGND VGND VPWR VPWR _17863_/A sky130_fd_sc_hd__buf_2
XFILLER_15_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14326_ _12460_/A _14321_/X _14325_/X VGND VGND VPWR VPWR _14326_/X sky130_fd_sc_hd__or3_4
X_11538_ _11538_/A _11538_/B VGND VGND VPWR VPWR _11538_/X sky130_fd_sc_hd__or2_4
X_18094_ _16943_/A _18093_/Y _16985_/X VGND VGND VPWR VPWR _23021_/B sky130_fd_sc_hd__o21a_4
XANTENNA__21672__A2 _21669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21030__A _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17045_ _12116_/Y _17016_/X _17023_/X _17044_/Y VGND VGND VPWR VPWR _17046_/B sky130_fd_sc_hd__o22a_4
XFILLER_99_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13748__A _11648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14257_ _14371_/A _14257_/B _14257_/C VGND VGND VPWR VPWR _14257_/X sky130_fd_sc_hd__and3_4
XANTENNA__12652__A _12652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13208_ _12373_/A VGND VGND VPWR VPWR _13239_/A sky130_fd_sc_hd__buf_2
XANTENNA__21424__A2 _21419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14188_ _14205_/A _23721_/Q VGND VGND VPWR VPWR _14189_/C sky130_fd_sc_hd__or2_4
XFILLER_67_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15963__A _16095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13139_ _15654_/A _13137_/X _13139_/C VGND VGND VPWR VPWR _13139_/X sky130_fd_sc_hd__and3_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18996_ _18996_/A VGND VGND VPWR VPWR _18996_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17947_ _17765_/X _17946_/X _17765_/X _17946_/X VGND VGND VPWR VPWR _17947_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21188__B2 _21187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13483__A _13483_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17878_ _18390_/A VGND VGND VPWR VPWR _17878_/X sky130_fd_sc_hd__buf_2
XFILLER_66_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16829_ _15928_/X _16239_/X _16521_/Y VGND VGND VPWR VPWR _16829_/X sky130_fd_sc_hd__o21a_4
X_19617_ _20754_/A _19551_/X _19615_/X _19616_/X VGND VGND VPWR VPWR _19617_/X sky130_fd_sc_hd__a211o_4
XFILLER_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12099__A _12068_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19548_ _19447_/X _19547_/X _18760_/C _19493_/X VGND VGND VPWR VPWR _19548_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__22688__A1 _21249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22688__B2 _22683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19479_ _19561_/A _19526_/B _19481_/B VGND VGND VPWR VPWR _19536_/A sky130_fd_sc_hd__a21oi_4
XFILLER_107_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20163__A2 IRQ[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21360__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21510_ _21795_/A VGND VGND VPWR VPWR _21510_/X sky130_fd_sc_hd__buf_2
XANTENNA__11731__A _16071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15203__A _15203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22490_ _22483_/A VGND VGND VPWR VPWR _22490_/X sky130_fd_sc_hd__buf_2
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18108__A2 _17913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12546__B _12667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21441_ _21282_/X _21440_/X _14696_/B _21437_/X VGND VGND VPWR VPWR _23812_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24160_ _24165_/CLK _19883_/Y HRESETn VGND VGND VPWR VPWR _17030_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_33_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21372_ _21251_/X _21369_/X _13257_/B _21366_/X VGND VGND VPWR VPWR _23857_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22860__A1 _16008_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21663__A2 _21662_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23111_ _23816_/CLK _23111_/D VGND VGND VPWR VPWR _13814_/B sky130_fd_sc_hd__dfxtp_4
X_20323_ _24412_/Q _18814_/X _24444_/Q _20260_/X VGND VGND VPWR VPWR _20323_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13658__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24091_ _24026_/CLK _20357_/X VGND VGND VPWR VPWR _24091_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12562__A _13908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23042_ _19901_/X _16939_/A _16988_/X _17944_/X _22889_/X VGND VGND VPWR VPWR _23042_/X
+ sky130_fd_sc_hd__o32a_4
X_20254_ _20253_/X VGND VGND VPWR VPWR _20255_/A sky130_fd_sc_hd__buf_2
XANTENNA__21415__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22612__B2 _22576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15873__A _13494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18292__A1 _17674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20185_ _18755_/X _20057_/X _20184_/Y _19929_/X VGND VGND VPWR VPWR _20185_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14489__A _15435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21179__B2 _21173_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23944_ _24008_/CLK _21199_/X VGND VGND VPWR VPWR _13652_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20926__A1 _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11625__B _11624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23875_ _23494_/CLK _21342_/X VGND VGND VPWR VPWR _14819_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22826_ _22778_/Y VGND VGND VPWR VPWR _22826_/X sky130_fd_sc_hd__buf_2
XFILLER_38_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14936__B _14879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21115__A _21130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22757_ _22756_/A _22755_/B VGND VGND VPWR VPWR _22758_/B sky130_fd_sc_hd__or2_4
XFILLER_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12737__A _12737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11641__A _14177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12510_ _13641_/A VGND VGND VPWR VPWR _13623_/A sky130_fd_sc_hd__buf_2
XANTENNA__15113__A _11710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13490_ _12876_/A _13486_/X _13490_/C VGND VGND VPWR VPWR _13491_/B sky130_fd_sc_hd__or3_4
X_21708_ _21536_/X _21705_/X _13153_/B _21702_/X VGND VGND VPWR VPWR _23665_/D sky130_fd_sc_hd__o22a_4
X_22688_ _21249_/A _22686_/X _13119_/B _22683_/X VGND VGND VPWR VPWR _22688_/X sky130_fd_sc_hd__o22a_4
XFILLER_51_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12456__B _12586_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12441_ _12441_/A VGND VGND VPWR VPWR _12850_/A sky130_fd_sc_hd__buf_2
X_21639_ _21633_/Y _21638_/X _21504_/X _21638_/X VGND VGND VPWR VPWR _23710_/D sky130_fd_sc_hd__a2bb2o_4
X_24427_ _24334_/CLK _24427_/D HRESETn VGND VGND VPWR VPWR _20706_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18424__A _18107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16870__C _16868_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13592__A1 _13493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12372_ _12418_/A _12274_/B VGND VGND VPWR VPWR _12372_/X sky130_fd_sc_hd__or2_4
X_15160_ _14098_/A _15158_/X _15159_/X VGND VGND VPWR VPWR _15160_/X sky130_fd_sc_hd__and3_4
X_24358_ _24330_/CLK _24358_/D HRESETn VGND VGND VPWR VPWR _19072_/A sky130_fd_sc_hd__dfstp_4
XFILLER_5_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22851__A1 _12338_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21654__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_1_0_HCLK clkbuf_4_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14111_ _15010_/A VGND VGND VPWR VPWR _15019_/A sky130_fd_sc_hd__buf_2
X_15091_ _15110_/A _15023_/B VGND VGND VPWR VPWR _15091_/X sky130_fd_sc_hd__or2_4
X_23309_ _23986_/CLK _22317_/X VGND VGND VPWR VPWR _23309_/Q sky130_fd_sc_hd__dfxtp_4
X_24289_ _24301_/CLK _24289_/D HRESETn VGND VGND VPWR VPWR _19110_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24232__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14042_ _12568_/A _23946_/Q VGND VGND VPWR VPWR _14042_/X sky130_fd_sc_hd__or2_4
XANTENNA__22603__B2 _22597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13287__B _13287_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18850_ _17171_/X _18848_/X _24394_/Q _18849_/X VGND VGND VPWR VPWR _18850_/X sky130_fd_sc_hd__o22a_4
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17801_ _17911_/A VGND VGND VPWR VPWR _17801_/X sky130_fd_sc_hd__buf_2
XFILLER_67_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18781_ _18781_/A VGND VGND VPWR VPWR _18781_/X sky130_fd_sc_hd__buf_2
XFILLER_114_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15993_ _16097_/A _23640_/Q VGND VGND VPWR VPWR _15994_/C sky130_fd_sc_hd__or2_4
XFILLER_48_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17732_ _17731_/Y _17732_/B VGND VGND VPWR VPWR _17743_/A sky130_fd_sc_hd__or2_4
X_14944_ _14658_/A _14938_/X _14943_/X VGND VGND VPWR VPWR _14953_/B sky130_fd_sc_hd__or3_4
XFILLER_94_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20917__A1 _20872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20917__B2 _20839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17663_ _24130_/Q _17664_/B VGND VGND VPWR VPWR _17665_/A sky130_fd_sc_hd__nor2_4
X_14875_ _14895_/A _14875_/B VGND VGND VPWR VPWR _14875_/X sky130_fd_sc_hd__or2_4
X_19402_ _19399_/X _18560_/X _19399_/X _24199_/Q VGND VGND VPWR VPWR _19402_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16614_ _16799_/A _16614_/B VGND VGND VPWR VPWR _16614_/X sky130_fd_sc_hd__or2_4
XFILLER_62_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13826_ _13631_/A _13826_/B _13826_/C VGND VGND VPWR VPWR _13826_/X sky130_fd_sc_hd__and3_4
X_17594_ _17594_/A VGND VGND VPWR VPWR _17594_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19333_ _19332_/X _18337_/X _19332_/X _24240_/Q VGND VGND VPWR VPWR _24240_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16545_ _16586_/A VGND VGND VPWR VPWR _16567_/A sky130_fd_sc_hd__buf_2
X_13757_ _15494_/A _13757_/B VGND VGND VPWR VPWR _13757_/X sky130_fd_sc_hd__or2_4
XANTENNA__12647__A _12591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21342__B2 _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15023__A _15023_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12708_ _12240_/A _23572_/Q VGND VGND VPWR VPWR _12709_/C sky130_fd_sc_hd__or2_4
X_19264_ _24272_/Q _19220_/X _19263_/Y VGND VGND VPWR VPWR _19264_/X sky130_fd_sc_hd__o21a_4
X_16476_ _16158_/A _22304_/A VGND VGND VPWR VPWR _16478_/B sky130_fd_sc_hd__or2_4
XANTENNA__21893__A2 _21887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13688_ _13688_/A VGND VGND VPWR VPWR _14207_/A sky130_fd_sc_hd__buf_2
X_18215_ _17794_/X _18212_/Y _18076_/X _18214_/X VGND VGND VPWR VPWR _18215_/X sky130_fd_sc_hd__a211o_4
X_15427_ _15431_/A _15425_/X _15427_/C VGND VGND VPWR VPWR _15428_/C sky130_fd_sc_hd__and3_4
Xclkbuf_7_17_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR _24250_/CLK sky130_fd_sc_hd__clkbuf_1
X_12639_ _12591_/X _12639_/B VGND VGND VPWR VPWR _12639_/X sky130_fd_sc_hd__or2_4
X_19195_ _19112_/B VGND VGND VPWR VPWR _19195_/Y sky130_fd_sc_hd__inv_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18146_ _17796_/X _18145_/X _17836_/X _18117_/X VGND VGND VPWR VPWR _18146_/X sky130_fd_sc_hd__o22a_4
X_15358_ _14010_/A _15292_/B VGND VGND VPWR VPWR _15360_/B sky130_fd_sc_hd__or2_4
XANTENNA__17849__B2 _17848_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22842__A1 _17439_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14309_ _15553_/A _14309_/B VGND VGND VPWR VPWR _14309_/X sky130_fd_sc_hd__or2_4
XANTENNA__13478__A _13477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18077_ _17864_/X _17235_/X _17866_/X VGND VGND VPWR VPWR _18077_/X sky130_fd_sc_hd__o21a_4
XFILLER_32_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15289_ _14149_/A _15289_/B VGND VGND VPWR VPWR _15289_/X sky130_fd_sc_hd__or2_4
X_17028_ _17028_/A _17561_/B VGND VGND VPWR VPWR _17028_/X sky130_fd_sc_hd__and2_4
XANTENNA__21695__A _21687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15693__A _15693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18979_ _24374_/Q VGND VGND VPWR VPWR _18979_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11726__A _15743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21990_ _21819_/X _21988_/X _23506_/Q _21985_/X VGND VGND VPWR VPWR _23506_/D sky130_fd_sc_hd__o22a_4
XFILLER_39_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20941_ _20842_/X _20939_/X _20940_/X HRDATA[10] _20847_/X VGND VGND VPWR VPWR _20941_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_27_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13941__A _12302_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20872_ _20279_/A VGND VGND VPWR VPWR _20872_/X sky130_fd_sc_hd__buf_2
X_23660_ _23404_/CLK _21715_/X VGND VGND VPWR VPWR _15406_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22611_ _22458_/X _22607_/X _15149_/B _22576_/A VGND VGND VPWR VPWR _23137_/D sky130_fd_sc_hd__o22a_4
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23591_ _23591_/CLK _21846_/X VGND VGND VPWR VPWR _23591_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_74_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12557__A _12922_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16029__A _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22530__B1 _16019_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22542_ _22425_/X _22536_/X _13434_/B _22540_/X VGND VGND VPWR VPWR _22542_/X sky130_fd_sc_hd__o22a_4
X_22473_ _22390_/X _22472_/X _12177_/B _22469_/X VGND VGND VPWR VPWR _22473_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15868__A _13548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14772__A _15443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18244__A _18244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21424_ _21253_/X _21419_/X _13326_/B _21423_/X VGND VGND VPWR VPWR _23824_/D sky130_fd_sc_hd__o22a_4
X_24212_ _24239_/CLK _19383_/X HRESETn VGND VGND VPWR VPWR _24212_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19376__A1_N _19374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21097__B1 _24009_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22833__A1 _13350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15587__B _23723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24143_ _24230_/CLK _24143_/D HRESETn VGND VGND VPWR VPWR _24143_/Q sky130_fd_sc_hd__dfrtp_4
X_21355_ _21369_/A VGND VGND VPWR VPWR _21355_/X sky130_fd_sc_hd__buf_2
XANTENNA__12292__A _15688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20306_ _20292_/X _20304_/X _19138_/A _20305_/X VGND VGND VPWR VPWR _20306_/X sky130_fd_sc_hd__o22a_4
X_24074_ _23819_/CLK _24074_/D VGND VGND VPWR VPWR _24074_/Q sky130_fd_sc_hd__dfxtp_4
X_21286_ _21285_/X _21283_/X _14802_/B _21278_/X VGND VGND VPWR VPWR _23907_/D sky130_fd_sc_hd__o22a_4
XFILLER_85_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23025_ _23025_/A VGND VGND VPWR VPWR HADDR[24] sky130_fd_sc_hd__inv_2
XFILLER_46_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20237_ _20424_/A VGND VGND VPWR VPWR _20447_/A sky130_fd_sc_hd__buf_2
XFILLER_2_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22061__A2 _22059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20168_ _11570_/X _20168_/B VGND VGND VPWR VPWR _20169_/B sky130_fd_sc_hd__or2_4
XFILLER_77_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16211__B _16211_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22349__B1 _16103_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15108__A _15108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19314__A1_N _19303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19803__A _19876_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12990_ _12989_/X VGND VGND VPWR VPWR _12990_/X sky130_fd_sc_hd__buf_2
X_20099_ _11559_/B VGND VGND VPWR VPWR _20099_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14012__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11941_ _16143_/A VGND VGND VPWR VPWR _11998_/A sky130_fd_sc_hd__buf_2
X_23927_ _23632_/CLK _21238_/X VGND VGND VPWR VPWR _16181_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18419__A _18295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17323__A _15379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14660_ _14925_/A VGND VGND VPWR VPWR _15107_/A sky130_fd_sc_hd__buf_2
X_11872_ _12493_/A VGND VGND VPWR VPWR _11872_/X sky130_fd_sc_hd__buf_2
X_23858_ _23794_/CLK _23858_/D VGND VGND VPWR VPWR _13123_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13611_ _13611_/A VGND VGND VPWR VPWR _13800_/A sky130_fd_sc_hd__buf_2
XFILLER_109_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22809_ _22792_/X _22809_/B VGND VGND VPWR VPWR HWDATA[11] sky130_fd_sc_hd__nor2_4
XFILLER_77_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14591_ _14161_/A _14680_/B VGND VGND VPWR VPWR _14591_/X sky130_fd_sc_hd__or2_4
XFILLER_60_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23789_ _23794_/CLK _23789_/D VGND VGND VPWR VPWR _15836_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12467__A _13651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21324__B2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16330_ _13422_/A _16330_/B _16330_/C VGND VGND VPWR VPWR _16338_/B sky130_fd_sc_hd__or3_4
X_13542_ _13558_/A _23599_/Q VGND VGND VPWR VPWR _13544_/B sky130_fd_sc_hd__or2_4
XFILLER_38_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16261_ _15976_/A _16259_/X _16260_/X VGND VGND VPWR VPWR _16261_/X sky130_fd_sc_hd__and3_4
XANTENNA__15778__A _12989_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13473_ _13450_/A _13554_/B VGND VGND VPWR VPWR _13474_/C sky130_fd_sc_hd__or2_4
XANTENNA__21499__B _21348_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18000_ _17954_/X _17960_/Y _17987_/X _17996_/X _17999_/Y VGND VGND VPWR VPWR _18000_/X
+ sky130_fd_sc_hd__a32o_4
X_15212_ _14251_/A _15212_/B VGND VGND VPWR VPWR _15212_/X sky130_fd_sc_hd__or2_4
XFILLER_16_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12424_ _12386_/X _12424_/B VGND VGND VPWR VPWR _12425_/C sky130_fd_sc_hd__or2_4
XANTENNA__21627__A2 _21626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16192_ _16223_/A _23671_/Q VGND VGND VPWR VPWR _16194_/B sky130_fd_sc_hd__or2_4
XFILLER_12_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15143_ _14143_/A _15213_/B VGND VGND VPWR VPWR _15143_/X sky130_fd_sc_hd__or2_4
XANTENNA__13298__A _12914_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12355_ _12826_/A _12228_/B VGND VGND VPWR VPWR _12355_/X sky130_fd_sc_hd__or2_4
X_12286_ _12211_/X VGND VGND VPWR VPWR _12286_/X sky130_fd_sc_hd__buf_2
X_15074_ _15074_/A VGND VGND VPWR VPWR _15110_/A sky130_fd_sc_hd__buf_2
X_19951_ _18745_/Y _19950_/X VGND VGND VPWR VPWR _19951_/X sky130_fd_sc_hd__or2_4
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22404__A _22416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14025_ _11647_/A _14025_/B VGND VGND VPWR VPWR _14025_/X sky130_fd_sc_hd__or2_4
X_18902_ _15911_/X _18898_/X _24365_/Q _18899_/X VGND VGND VPWR VPWR _18902_/X sky130_fd_sc_hd__o22a_4
X_19882_ _19554_/X _19880_/X _19881_/X _19581_/X _19808_/A VGND VGND VPWR VPWR _19882_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12930__A _12982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18833_ _12674_/X _18827_/X _20469_/A _18828_/X VGND VGND VPWR VPWR _24405_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13745__B _13745_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18764_ _18788_/A VGND VGND VPWR VPWR _18781_/A sky130_fd_sc_hd__buf_2
X_15976_ _15976_/A _15974_/X _15976_/C VGND VGND VPWR VPWR _15976_/X sky130_fd_sc_hd__and3_4
XFILLER_114_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17715_ _17748_/A VGND VGND VPWR VPWR _17716_/A sky130_fd_sc_hd__inv_2
X_14927_ _11646_/A _14863_/B VGND VGND VPWR VPWR _14929_/B sky130_fd_sc_hd__or2_4
XFILLER_49_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18695_ _17794_/A _17871_/B _17933_/X _18694_/X VGND VGND VPWR VPWR _18695_/X sky130_fd_sc_hd__a211o_4
XFILLER_35_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13761__A _13737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17646_ _17646_/A _17646_/B VGND VGND VPWR VPWR _17647_/A sky130_fd_sc_hd__or2_4
X_14858_ _13955_/A _14856_/X _14857_/X VGND VGND VPWR VPWR _14858_/X sky130_fd_sc_hd__and3_4
XFILLER_63_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14576__B _14654_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13809_ _15424_/A _13807_/X _13808_/X VGND VGND VPWR VPWR _13809_/X sky130_fd_sc_hd__and3_4
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13480__B _13568_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17577_ _17532_/Y _17569_/X _17576_/X VGND VGND VPWR VPWR _17577_/X sky130_fd_sc_hd__o21a_4
X_14789_ _13690_/A _14787_/X _14789_/C VGND VGND VPWR VPWR _14789_/X sky130_fd_sc_hd__and3_4
XANTENNA__12377__A _15882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21315__B2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19316_ _19313_/X _17947_/X _19313_/X _24251_/Q VGND VGND VPWR VPWR _19316_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16528_ _16536_/A _23516_/Q VGND VGND VPWR VPWR _16529_/C sky130_fd_sc_hd__or2_4
XFILLER_31_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18192__B1 _18048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16791__B _16791_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18731__A2 _18730_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19247_ _19247_/A VGND VGND VPWR VPWR _19247_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15688__A _15688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16459_ _16464_/A _16390_/B VGND VGND VPWR VPWR _16459_/X sky130_fd_sc_hd__or2_4
XANTENNA__14592__A _14737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16742__A1 _11992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18064__A _18205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19178_ _19120_/A _19120_/B _19177_/Y VGND VGND VPWR VPWR _24299_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21618__A2 _21612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18999__A _18999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12824__B _23796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18129_ _18129_/A VGND VGND VPWR VPWR _18129_/X sky130_fd_sc_hd__buf_2
XFILLER_8_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22291__A2 _22286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19692__B1 _19877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21140_ _21133_/A VGND VGND VPWR VPWR _21140_/X sky130_fd_sc_hd__buf_2
XANTENNA__13001__A _12879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21071_ _20356_/X _21068_/X _24027_/Q _21065_/X VGND VGND VPWR VPWR _24027_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13936__A _15037_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22043__A2 _22038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12840__A _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16312__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20022_ _20018_/X _17674_/A _20000_/X _20021_/X VGND VGND VPWR VPWR _20023_/A sky130_fd_sc_hd__o22a_4
XFILLER_100_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21003__B1 _24063_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21973_ _22002_/A VGND VGND VPWR VPWR _21988_/A sky130_fd_sc_hd__buf_2
XFILLER_39_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0_0_HCLK_A clkbuf_2_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14767__A _13800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21554__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13671__A _12233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23712_ _23073_/CLK _21631_/X VGND VGND VPWR VPWR _14860_/B sky130_fd_sc_hd__dfxtp_4
X_20924_ _20921_/X _20923_/X _20240_/X VGND VGND VPWR VPWR _20924_/Y sky130_fd_sc_hd__o21ai_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14486__B _14486_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _20855_/A VGND VGND VPWR VPWR _20855_/Y sky130_fd_sc_hd__inv_2
X_23643_ _23515_/CLK _23643_/D VGND VGND VPWR VPWR _23643_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12287__A _12286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21306__A1 _21221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21306__B2 _21302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20786_ _20681_/X _20785_/X _19062_/A _20625_/X VGND VGND VPWR VPWR _20786_/X sky130_fd_sc_hd__o22a_4
X_23574_ _23539_/CLK _23574_/D VGND VGND VPWR VPWR _12271_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22525_ _22396_/X _22522_/X _16754_/B _22519_/X VGND VGND VPWR VPWR _22525_/X sky130_fd_sc_hd__o22a_4
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22456_ _22456_/A VGND VGND VPWR VPWR _22456_/X sky130_fd_sc_hd__buf_2
XFILLER_6_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20009__A _19985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_63_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR _23826_/CLK sky130_fd_sc_hd__clkbuf_1
X_21407_ _21225_/X _21405_/X _23836_/Q _21402_/X VGND VGND VPWR VPWR _21407_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15110__B _24063_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22387_ _22386_/X VGND VGND VPWR VPWR _22387_/X sky130_fd_sc_hd__buf_2
XANTENNA__22282__A2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14007__A _11738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12140_ _11829_/A _12140_/B VGND VGND VPWR VPWR _12141_/C sky130_fd_sc_hd__or2_4
XFILLER_68_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21338_ _21277_/X _21333_/X _14301_/B _21337_/X VGND VGND VPWR VPWR _23878_/D sky130_fd_sc_hd__o22a_4
X_24126_ _24126_/CLK _20028_/Y HRESETn VGND VGND VPWR VPWR _24126_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12071_ _12098_/A _23549_/Q VGND VGND VPWR VPWR _12072_/C sky130_fd_sc_hd__or2_4
X_21269_ _21268_/X _21259_/X _23914_/Q _21266_/X VGND VGND VPWR VPWR _23914_/D sky130_fd_sc_hd__o22a_4
X_24057_ _23514_/CLK _24057_/D VGND VGND VPWR VPWR _24057_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16222__A _16198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23008_ _23003_/A _18172_/Y VGND VGND VPWR VPWR _23008_/Y sky130_fd_sc_hd__nand2_4
XFILLER_49_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15830_ _12522_/A _15828_/X _15829_/X VGND VGND VPWR VPWR _15834_/B sky130_fd_sc_hd__and3_4
XANTENNA__24155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15761_ _13102_/A _15753_/X _15760_/X VGND VGND VPWR VPWR _15761_/X sky130_fd_sc_hd__and3_4
XFILLER_64_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15780__B _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12973_ _12949_/A _23091_/Q VGND VGND VPWR VPWR _12975_/B sky130_fd_sc_hd__or2_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20348__A2 _20347_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17500_ _17499_/X VGND VGND VPWR VPWR _17500_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21545__B2 _21539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14712_ _14673_/A _14712_/B _14712_/C VGND VGND VPWR VPWR _14712_/X sky130_fd_sc_hd__and3_4
XFILLER_46_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11924_ _11924_/A _11904_/X _11923_/X VGND VGND VPWR VPWR _11924_/X sky130_fd_sc_hd__or3_4
X_18480_ _18198_/A VGND VGND VPWR VPWR _18480_/X sky130_fd_sc_hd__buf_2
X_15692_ _12735_/A _15757_/B VGND VGND VPWR VPWR _15692_/X sky130_fd_sc_hd__or2_4
XFILLER_45_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17431_ _15646_/X _17348_/B VGND VGND VPWR VPWR _17431_/Y sky130_fd_sc_hd__nand2_4
XFILLER_75_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14643_ _14197_/A VGND VGND VPWR VPWR _14644_/A sky130_fd_sc_hd__buf_2
XFILLER_2_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17988__A _18189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11855_ _12529_/A VGND VGND VPWR VPWR _13986_/A sky130_fd_sc_hd__buf_2
XFILLER_61_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17362_ _17361_/X VGND VGND VPWR VPWR _17382_/B sky130_fd_sc_hd__inv_2
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14574_ _15142_/A _14652_/B VGND VGND VPWR VPWR _14574_/X sky130_fd_sc_hd__or2_4
X_11786_ _11818_/A _21683_/A VGND VGND VPWR VPWR _11788_/B sky130_fd_sc_hd__or2_4
X_19101_ _20968_/A _18941_/X _11504_/Y _18946_/X VGND VGND VPWR VPWR _19101_/Y sky130_fd_sc_hd__a22oi_4
X_16313_ _13415_/A _16306_/X _16312_/X VGND VGND VPWR VPWR _16313_/X sky130_fd_sc_hd__or3_4
X_13525_ _12981_/A VGND VGND VPWR VPWR _13562_/A sky130_fd_sc_hd__buf_2
X_17293_ _14565_/Y _17295_/B VGND VGND VPWR VPWR _18583_/B sky130_fd_sc_hd__or2_4
XANTENNA__12925__A _12958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19032_ _11518_/B VGND VGND VPWR VPWR _19032_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16244_ _16243_/X _16244_/B VGND VGND VPWR VPWR _16244_/X sky130_fd_sc_hd__or2_4
XANTENNA__15301__A _14737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13456_ _12868_/A _13456_/B VGND VGND VPWR VPWR _13458_/B sky130_fd_sc_hd__or2_4
XFILLER_16_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12407_ _13102_/A _12407_/B _12406_/X VGND VGND VPWR VPWR _12407_/X sky130_fd_sc_hd__and3_4
XANTENNA__15020__B _15088_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16175_ _16223_/A _16175_/B VGND VGND VPWR VPWR _16178_/B sky130_fd_sc_hd__or2_4
XFILLER_51_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22273__A2 _22272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13387_ _13378_/X _23536_/Q VGND VGND VPWR VPWR _13387_/X sky130_fd_sc_hd__or2_4
X_15126_ _12209_/A _15126_/B VGND VGND VPWR VPWR _15127_/C sky130_fd_sc_hd__or2_4
X_12338_ _12338_/A VGND VGND VPWR VPWR _12338_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22134__A _22134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15057_ _12583_/A _23711_/Q VGND VGND VPWR VPWR _15058_/C sky130_fd_sc_hd__or2_4
X_19934_ _20000_/A VGND VGND VPWR VPWR _19934_/X sky130_fd_sc_hd__buf_2
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12269_ _12269_/A VGND VGND VPWR VPWR _13026_/A sky130_fd_sc_hd__buf_2
XFILLER_64_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14008_ _14008_/A VGND VGND VPWR VPWR _14847_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_5_17_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21973__A _22002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19865_ _19531_/X _19864_/X _20194_/A _19531_/X VGND VGND VPWR VPWR _24164_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15971__A _11933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18816_ _18815_/X VGND VGND VPWR VPWR _18841_/A sky130_fd_sc_hd__buf_2
XFILLER_110_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19796_ _19706_/A _19786_/Y _19787_/Y _19795_/X VGND VGND VPWR VPWR _19796_/X sky130_fd_sc_hd__a211o_4
XANTENNA__14266__A2 _14263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15690__B _15690_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15959_ _15959_/A VGND VGND VPWR VPWR _16096_/A sky130_fd_sc_hd__buf_2
X_18747_ _17007_/X _17081_/A _17077_/A _18746_/Y VGND VGND VPWR VPWR _18747_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14587__A _14146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13491__A _13491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18678_ _18677_/X VGND VGND VPWR VPWR _18678_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12029__A1 _11844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17629_ _17629_/A VGND VGND VPWR VPWR _17629_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12029__B2 _12028_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20640_ _20492_/A VGND VGND VPWR VPWR _20640_/X sky130_fd_sc_hd__buf_2
XANTENNA__21839__A2 _21829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20571_ _20534_/A _20570_/X VGND VGND VPWR VPWR _20571_/X sky130_fd_sc_hd__or2_4
XANTENNA__16307__A _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22310_ _23316_/Q VGND VGND VPWR VPWR _23316_/D sky130_fd_sc_hd__buf_2
X_23290_ _23354_/CLK _23290_/D VGND VGND VPWR VPWR _16391_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16026__B _15952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22241_ _22131_/X _22236_/X _14311_/B _22240_/X VGND VGND VPWR VPWR _22241_/X sky130_fd_sc_hd__o22a_4
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18522__A _18216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20275__B2 _20484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22172_ _22172_/A VGND VGND VPWR VPWR _22172_/X sky130_fd_sc_hd__buf_2
XFILLER_106_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21123_ _21115_/X VGND VGND VPWR VPWR _21123_/X sky130_fd_sc_hd__buf_2
XANTENNA__13666__A _15411_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22570__A2_N _22569_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12570__A _15487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21224__B1 _23933_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21054_ _20937_/X _21051_/X _15352_/B _21048_/X VGND VGND VPWR VPWR _24034_/D sky130_fd_sc_hd__o22a_4
XFILLER_43_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16977__A _17680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20005_ _24468_/Q VGND VGND VPWR VPWR _20005_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21775__B2 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15881__A _13529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_HCLK clkbuf_4_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22724__B1 HREADY VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11914__A _11913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21956_ _21935_/A VGND VGND VPWR VPWR _21956_/X sky130_fd_sc_hd__buf_2
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _20759_/X _20906_/X _19112_/A _20769_/X VGND VGND VPWR VPWR _20908_/B sky130_fd_sc_hd__o22a_4
XANTENNA__15105__B _23679_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19800__B _19800_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ _21887_/A VGND VGND VPWR VPWR _21887_/X sky130_fd_sc_hd__buf_2
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _13688_/A VGND VGND VPWR VPWR _14177_/A sky130_fd_sc_hd__buf_2
X_23626_ _23819_/CLK _23626_/D VGND VGND VPWR VPWR _23626_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _20838_/A VGND VGND VPWR VPWR _20838_/X sky130_fd_sc_hd__buf_2
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14944__B _14938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22219__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21123__A _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _24443_/Q IRQ[28] VGND VGND VPWR VPWR _20166_/A sky130_fd_sc_hd__and2_4
X_23557_ _23557_/CLK _23557_/D VGND VGND VPWR VPWR _14516_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20769_ _20242_/X VGND VGND VPWR VPWR _20769_/X sky130_fd_sc_hd__buf_2
XFILLER_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12745__A _12745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _12255_/X _13308_/X _13309_/X VGND VGND VPWR VPWR _13310_/X sky130_fd_sc_hd__and3_4
XANTENNA__16880__A1_N _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22508_ _22451_/X _22507_/X _14627_/B _22504_/X VGND VGND VPWR VPWR _23204_/D sky130_fd_sc_hd__o22a_4
X_14290_ _11911_/A _14290_/B _14290_/C VGND VGND VPWR VPWR _14290_/X sky130_fd_sc_hd__and3_4
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23488_ _23391_/CLK _23488_/D VGND VGND VPWR VPWR _14857_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ _13260_/A _13174_/B VGND VGND VPWR VPWR _13243_/B sky130_fd_sc_hd__or2_4
X_22439_ _20778_/A VGND VGND VPWR VPWR _22439_/X sky130_fd_sc_hd__buf_2
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13172_ _12722_/A _23953_/Q VGND VGND VPWR VPWR _13173_/C sky130_fd_sc_hd__or2_4
XFILLER_87_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12123_ _12167_/A _12123_/B VGND VGND VPWR VPWR _12123_/X sky130_fd_sc_hd__or2_4
X_24109_ _24203_/CLK _24109_/D HRESETn VGND VGND VPWR VPWR _17736_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17048__A _17007_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13576__A _13575_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17980_ _17969_/X _17974_/X _17975_/X _17979_/X VGND VGND VPWR VPWR _17980_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22007__A2 _22002_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12480__A _12528_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12054_ _12044_/X _12054_/B _12054_/C VGND VGND VPWR VPWR _12061_/B sky130_fd_sc_hd__and3_4
X_16931_ _17062_/A VGND VGND VPWR VPWR _16931_/X sky130_fd_sc_hd__buf_2
XFILLER_2_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21793__A _21817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15791__A _12443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16862_ _16861_/X VGND VGND VPWR VPWR _16865_/C sky130_fd_sc_hd__inv_2
X_19650_ _19497_/X HRDATA[9] _20400_/B _19496_/X VGND VGND VPWR VPWR _19650_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_77_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15813_ _12682_/X _15790_/X _15797_/X _15804_/X _15812_/X VGND VGND VPWR VPWR _15813_/X
+ sky130_fd_sc_hd__a32o_4
X_18601_ _18554_/X _18600_/X _20079_/A _18554_/X VGND VGND VPWR VPWR _24454_/D sky130_fd_sc_hd__a2bb2o_4
X_19581_ _19580_/X VGND VGND VPWR VPWR _19581_/X sky130_fd_sc_hd__buf_2
X_16793_ _16747_/X _16791_/X _16793_/C VGND VGND VPWR VPWR _16793_/X sky130_fd_sc_hd__and3_4
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23810__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20202__A _20488_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21518__B2 _21515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18532_ _18512_/X _18531_/X _20058_/A _18512_/X VGND VGND VPWR VPWR _24457_/D sky130_fd_sc_hd__a2bb2o_4
X_15744_ _11680_/X _15744_/B _15743_/X VGND VGND VPWR VPWR _15744_/X sky130_fd_sc_hd__or3_4
X_12956_ _13118_/A _12948_/X _12956_/C VGND VGND VPWR VPWR _12957_/C sky130_fd_sc_hd__and3_4
XANTENNA__14200__A _14215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12639__B _12639_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22191__B2 _22190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11907_ _12250_/A VGND VGND VPWR VPWR _14998_/A sky130_fd_sc_hd__buf_2
X_18463_ _18463_/A VGND VGND VPWR VPWR _18463_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11543__B IRQ[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15675_ _12709_/A _15675_/B _15675_/C VGND VGND VPWR VPWR _15679_/B sky130_fd_sc_hd__and3_4
X_12887_ _12887_/A _12879_/X _12886_/X VGND VGND VPWR VPWR _12887_/X sky130_fd_sc_hd__and3_4
X_17414_ _17411_/Y _17340_/X _17021_/A _17413_/X VGND VGND VPWR VPWR _17414_/X sky130_fd_sc_hd__o22a_4
X_14626_ _12449_/A _14626_/B _14625_/X VGND VGND VPWR VPWR _14626_/X sky130_fd_sc_hd__and3_4
X_11838_ _11592_/A VGND VGND VPWR VPWR _11838_/Y sky130_fd_sc_hd__inv_2
X_18394_ _17622_/B _17602_/B VGND VGND VPWR VPWR _18395_/C sky130_fd_sc_hd__and2_4
XFILLER_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22129__A _22129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17345_ _16894_/A _17364_/A _17365_/A VGND VGND VPWR VPWR _17345_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14557_ _11648_/X _14479_/B VGND VGND VPWR VPWR _14557_/X sky130_fd_sc_hd__or2_4
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11769_ _13102_/A VGND VGND VPWR VPWR _12822_/A sky130_fd_sc_hd__buf_2
XANTENNA__12655__A _12655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22494__A2 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19895__B1 _19894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15031__A _14617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13508_ _15876_/A _13434_/B VGND VGND VPWR VPWR _13508_/X sky130_fd_sc_hd__or2_4
XANTENNA__18162__A3 _18148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17276_ _17275_/X VGND VGND VPWR VPWR _17278_/B sky130_fd_sc_hd__inv_2
X_14488_ _13796_/A _14488_/B _14487_/X VGND VGND VPWR VPWR _14489_/C sky130_fd_sc_hd__and3_4
XANTENNA__20872__A _20279_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21117__A2_N _21116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19015_ _18994_/X _19013_/Y _19014_/Y _18999_/X VGND VGND VPWR VPWR _19015_/X sky130_fd_sc_hd__o22a_4
X_16227_ _16227_/A _23639_/Q VGND VGND VPWR VPWR _16228_/C sky130_fd_sc_hd__or2_4
X_13439_ _13463_/A _23279_/Q VGND VGND VPWR VPWR _13440_/C sky130_fd_sc_hd__or2_4
XANTENNA__15966__A _15937_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22246__A2 _22243_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16158_ _16158_/A _16158_/B VGND VGND VPWR VPWR _16158_/X sky130_fd_sc_hd__or2_4
XANTENNA__15685__B _15685_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17122__A1 _11912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15109_ _15109_/A _15033_/B VGND VGND VPWR VPWR _15109_/X sky130_fd_sc_hd__or2_4
XANTENNA__13486__A _12466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16089_ _12546_/A VGND VGND VPWR VPWR _16090_/A sky130_fd_sc_hd__buf_2
XANTENNA__12390__A _13557_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19917_ _22723_/A VGND VGND VPWR VPWR _19917_/X sky130_fd_sc_hd__buf_2
XANTENNA__21757__A1 _21534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21757__B2 _21752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19848_ _19839_/X _19847_/X _19592_/A VGND VGND VPWR VPWR _19848_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19779_ _19661_/A _19778_/X _19592_/A _19789_/B VGND VGND VPWR VPWR _19779_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21509__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20980__A2 _20873_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21810_ _21809_/X _21805_/X _12289_/B _21800_/X VGND VGND VPWR VPWR _21810_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15206__A _14246_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19901__A _22968_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22790_ _17283_/Y _22781_/X VGND VGND VPWR VPWR HWDATA[7] sky130_fd_sc_hd__nor2_4
XANTENNA__14110__A _14994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22182__A1 _22117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22182__B2 _22176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21741_ _21755_/A VGND VGND VPWR VPWR _21741_/X sky130_fd_sc_hd__buf_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24460_ _24126_/CLK _18457_/X HRESETn VGND VGND VPWR VPWR _20043_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_75_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21672_ _21560_/X _21669_/X _13831_/B _21666_/X VGND VGND VPWR VPWR _21672_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_4_13_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_26_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23411_ _23311_/CLK _22173_/X VGND VGND VPWR VPWR _23411_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20623_ _18813_/X VGND VGND VPWR VPWR _20623_/X sky130_fd_sc_hd__buf_2
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24391_ _24365_/CLK _24391_/D HRESETn VGND VGND VPWR VPWR _24391_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22485__A2 _22479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20496__A1 _20448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20554_ _20511_/X _20553_/X _24082_/Q _20488_/X VGND VGND VPWR VPWR _20554_/X sky130_fd_sc_hd__o22a_4
X_23342_ _23342_/CLK _23342_/D VGND VGND VPWR VPWR _15655_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20782__A _20400_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15876__A _15876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20485_ _24213_/Q _20398_/X _20484_/X VGND VGND VPWR VPWR _20486_/A sky130_fd_sc_hd__o21a_4
X_23273_ _23561_/CLK _23273_/D VGND VGND VPWR VPWR _23273_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22237__A2 _22236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14780__A _12509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19102__A2 _18999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22224_ _22103_/X _22222_/X _23378_/Q _22219_/X VGND VGND VPWR VPWR _23378_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21996__B2 _21992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22155_ _22162_/A VGND VGND VPWR VPWR _22155_/X sky130_fd_sc_hd__buf_2
XANTENNA__11909__A _11909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18861__A1 _15249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21106_ _20937_/X _21103_/X _15262_/B _21100_/X VGND VGND VPWR VPWR _24002_/D sky130_fd_sc_hd__o22a_4
X_22086_ _20393_/A VGND VGND VPWR VPWR _22086_/X sky130_fd_sc_hd__buf_2
XFILLER_87_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21037_ _21030_/A VGND VGND VPWR VPWR _21037_/X sky130_fd_sc_hd__buf_2
XFILLER_74_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20420__B2 _20374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21118__A _21118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12810_ _13563_/A _12810_/B _12810_/C VGND VGND VPWR VPWR _12814_/B sky130_fd_sc_hd__and3_4
XANTENNA__15116__A _14071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13790_ _13813_/A _13786_/X _13790_/C VGND VGND VPWR VPWR _13790_/X sky130_fd_sc_hd__or3_4
XANTENNA__14020__A _14020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22988_ _18309_/X _23004_/B VGND VGND VPWR VPWR _22988_/X sky130_fd_sc_hd__or2_4
XANTENNA__22173__A1 _22100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20957__A _22458_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22173__B2 _22169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12741_ _15820_/A _12737_/X _12740_/X VGND VGND VPWR VPWR _12741_/X sky130_fd_sc_hd__or3_4
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_0_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21939_ _21816_/X _21938_/X _12953_/B _21935_/X VGND VGND VPWR VPWR _21939_/X sky130_fd_sc_hd__o22a_4
XFILLER_31_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15460_ _12638_/A _15458_/X _15459_/X VGND VGND VPWR VPWR _15460_/X sky130_fd_sc_hd__and3_4
X_12672_ _12672_/A _12656_/X _12671_/X VGND VGND VPWR VPWR _12673_/C sky130_fd_sc_hd__or3_4
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23052__B _23038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23213__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14499_/A _14411_/B _14411_/C VGND VGND VPWR VPWR _14412_/C sky130_fd_sc_hd__and3_4
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11622_/X VGND VGND VPWR VPWR _20076_/A sky130_fd_sc_hd__inv_2
X_23609_ _23514_/CLK _23609_/D VGND VGND VPWR VPWR _23609_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _13776_/X _16840_/B _14267_/X _16840_/C VGND VGND VPWR VPWR _15391_/X sky130_fd_sc_hd__or4_4
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12475__A _12475_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _17130_/A VGND VGND VPWR VPWR _17130_/X sky130_fd_sc_hd__buf_2
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _14218_/X VGND VGND VPWR VPWR _15584_/A sky130_fd_sc_hd__buf_2
XANTENNA__21788__A _21787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11554_ _24423_/Q IRQ[8] VGND VGND VPWR VPWR _11554_/X sky130_fd_sc_hd__and2_4
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16155__A2 _11619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20692__A _20288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24377__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17061_ _16929_/B _17059_/X _20194_/A _11634_/B VGND VGND VPWR VPWR _17061_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15786__A _12849_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14273_ _13670_/A _14271_/X _14272_/X VGND VGND VPWR VPWR _14273_/X sky130_fd_sc_hd__and3_4
XANTENNA__22228__A2 _22222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14690__A _14673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16012_ _16048_/A VGND VGND VPWR VPWR _16058_/A sky130_fd_sc_hd__buf_2
X_13224_ _13260_/A _13165_/B VGND VGND VPWR VPWR _13224_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_33_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_66_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_3_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21987__B2 _21985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13155_ _12740_/A _13153_/X _13154_/X VGND VGND VPWR VPWR _13155_/X sky130_fd_sc_hd__and3_4
XANTENNA__18852__A1 _17178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12106_ _11996_/A _23101_/Q VGND VGND VPWR VPWR _12108_/B sky130_fd_sc_hd__or2_4
X_13086_ _13128_/A _13084_/X _13085_/X VGND VGND VPWR VPWR _13086_/X sky130_fd_sc_hd__and3_4
X_17963_ _17864_/X _17929_/X _17866_/X VGND VGND VPWR VPWR _17963_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21739__B2 _21738_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19702_ _19706_/A VGND VGND VPWR VPWR _19703_/A sky130_fd_sc_hd__inv_2
X_12037_ _11924_/A VGND VGND VPWR VPWR _16689_/A sky130_fd_sc_hd__buf_2
X_16914_ _16907_/C _16916_/A _16913_/X _16905_/X VGND VGND VPWR VPWR _16914_/X sky130_fd_sc_hd__or4_4
XFILLER_61_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22400__A2 _22392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17894_ _17893_/X _16977_/B _16999_/C _17894_/D VGND VGND VPWR VPWR _17894_/X sky130_fd_sc_hd__or4_4
XANTENNA__16410__A _11933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19633_ _19578_/X _19628_/X _19629_/X _19633_/D VGND VGND VPWR VPWR _19633_/X sky130_fd_sc_hd__or4_4
XFILLER_38_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16845_ _16837_/X _16839_/X _16843_/X _16845_/D VGND VGND VPWR VPWR _16845_/X sky130_fd_sc_hd__and4_4
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15026__A _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16776_ _16800_/A _23547_/Q VGND VGND VPWR VPWR _16777_/C sky130_fd_sc_hd__or2_4
X_19564_ _19422_/X _19563_/X HRDATA[7] _19438_/X VGND VGND VPWR VPWR _19621_/A sky130_fd_sc_hd__o22a_4
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13988_ _11976_/A _13965_/X _13972_/X _13979_/X _13987_/X VGND VGND VPWR VPWR _13988_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_34_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12369__B _12271_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15727_ _13082_/A _15727_/B _15727_/C VGND VGND VPWR VPWR _15728_/C sky130_fd_sc_hd__or3_4
X_18515_ _16971_/B VGND VGND VPWR VPWR _18515_/Y sky130_fd_sc_hd__inv_2
X_12939_ _12951_/A _12939_/B _12939_/C VGND VGND VPWR VPWR _12940_/C sky130_fd_sc_hd__and3_4
XFILLER_59_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19495_ HRDATA[30] VGND VGND VPWR VPWR _20650_/A sky130_fd_sc_hd__buf_2
XANTENNA__20714__A2 _20713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21911__B2 _21905_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17241__A _18728_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15658_ _12556_/A _15658_/B _15657_/X VGND VGND VPWR VPWR _15658_/X sky130_fd_sc_hd__or3_4
X_18446_ _18327_/A _18446_/B VGND VGND VPWR VPWR _18446_/X sky130_fd_sc_hd__and2_4
XFILLER_18_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14609_ _14117_/A _14607_/X _14608_/X VGND VGND VPWR VPWR _14613_/B sky130_fd_sc_hd__and3_4
X_18377_ _18224_/A VGND VGND VPWR VPWR _18377_/X sky130_fd_sc_hd__buf_2
X_15589_ _15589_/A _15589_/B _15589_/C VGND VGND VPWR VPWR _15589_/X sky130_fd_sc_hd__or3_4
XFILLER_33_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17328_ _14988_/X _17160_/A VGND VGND VPWR VPWR _17330_/A sky130_fd_sc_hd__or2_4
XFILLER_119_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21675__B1 _14486_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_115_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR _23635_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21698__A _21705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17259_ _17259_/A _17258_/Y VGND VGND VPWR VPWR _17259_/X sky130_fd_sc_hd__and2_4
XANTENNA__15696__A _15696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21427__B1 _15690_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20270_ _20270_/A _20270_/B _20269_/X VGND VGND VPWR VPWR _20270_/X sky130_fd_sc_hd__and3_4
XFILLER_66_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23856__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16304__B _16240_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18843__A1 _13575_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19615__B HRDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23960_ _24084_/CLK _21177_/X VGND VGND VPWR VPWR _23960_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16320__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22911_ _19201_/X _22911_/B _22911_/C VGND VGND VPWR VPWR HADDR[5] sky130_fd_sc_hd__and3_4
XFILLER_79_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23891_ _23827_/CLK _21320_/X VGND VGND VPWR VPWR _23891_/Q sky130_fd_sc_hd__dfxtp_4
X_22842_ _17439_/Y _22825_/X _22831_/X _22841_/X VGND VGND VPWR VPWR _22843_/A sky130_fd_sc_hd__a211o_4
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23236__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22773_ _22773_/A _22773_/B VGND VGND VPWR VPWR _22773_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21639__A2_N _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14775__A _13647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11614__D _13651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21902__B2 _21898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21724_ _21562_/X _21719_/X _14283_/B _21723_/X VGND VGND VPWR VPWR _23654_/D sky130_fd_sc_hd__o22a_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24443_ _24277_/CLK _18772_/X HRESETn VGND VGND VPWR VPWR _24443_/Q sky130_fd_sc_hd__dfrtp_4
X_21655_ _21662_/A VGND VGND VPWR VPWR _21655_/X sky130_fd_sc_hd__buf_2
XFILLER_40_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12295__A _12695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16990__A _17769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20606_ _20212_/X _20594_/X _20515_/X _20605_/Y VGND VGND VPWR VPWR _20606_/X sky130_fd_sc_hd__a211o_4
XFILLER_36_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24374_ _24277_/CLK _18889_/X HRESETn VGND VGND VPWR VPWR _24374_/Q sky130_fd_sc_hd__dfstp_4
X_21586_ _21590_/A VGND VGND VPWR VPWR _21602_/A sky130_fd_sc_hd__inv_2
XANTENNA__17334__A1 _15381_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23325_ _23485_/CLK _23325_/D VGND VGND VPWR VPWR _12146_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21401__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20537_ _21246_/A VGND VGND VPWR VPWR _20537_/X sky130_fd_sc_hd__buf_2
X_20468_ _20468_/A VGND VGND VPWR VPWR _20468_/X sky130_fd_sc_hd__buf_2
X_23256_ _23354_/CLK _23256_/D VGND VGND VPWR VPWR _23256_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12742__B _12823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22207_ _22207_/A VGND VGND VPWR VPWR _22222_/A sky130_fd_sc_hd__buf_2
XANTENNA__11639__A _13686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17637__A2 _17004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20399_ _20399_/A VGND VGND VPWR VPWR _20588_/A sky130_fd_sc_hd__buf_2
X_23187_ _23986_/CLK _23187_/D VGND VGND VPWR VPWR _12857_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22630__A2 _22629_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22138_ _22136_/X _22137_/X _14676_/B _22132_/X VGND VGND VPWR VPWR _22138_/X sky130_fd_sc_hd__o22a_4
XFILLER_47_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14960_ _11642_/A _14960_/B _14959_/X VGND VGND VPWR VPWR _14960_/X sky130_fd_sc_hd__and3_4
XANTENNA__17326__A _15249_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22069_ _22068_/X VGND VGND VPWR VPWR _22125_/A sky130_fd_sc_hd__buf_2
XANTENNA__16230__A _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23047__B _23038_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13911_ _13911_/A _13911_/B _13911_/C VGND VGND VPWR VPWR _13915_/B sky130_fd_sc_hd__and3_4
XFILLER_87_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14891_ _14895_/A _23584_/Q VGND VGND VPWR VPWR _14891_/X sky130_fd_sc_hd__or2_4
X_16630_ _16629_/X VGND VGND VPWR VPWR _16630_/X sky130_fd_sc_hd__buf_2
X_13842_ _11707_/A VGND VGND VPWR VPWR _14218_/A sky130_fd_sc_hd__buf_2
XFILLER_63_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22146__B2 _22071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16561_ _11936_/X _16561_/B _16560_/X VGND VGND VPWR VPWR _16562_/B sky130_fd_sc_hd__or3_4
XANTENNA__23063__A _20206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13773_ _13685_/Y _13772_/X VGND VGND VPWR VPWR _13776_/A sky130_fd_sc_hd__and2_4
X_15512_ _15512_/A _15512_/B VGND VGND VPWR VPWR _15513_/C sky130_fd_sc_hd__or2_4
X_18300_ _17837_/X _18034_/X _17846_/X _18036_/X VGND VGND VPWR VPWR _18300_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12724_ _15688_/A _12724_/B _12723_/X VGND VGND VPWR VPWR _12724_/X sky130_fd_sc_hd__or3_4
X_19280_ _19213_/A _19213_/B _19279_/Y VGND VGND VPWR VPWR _24264_/D sky130_fd_sc_hd__o21a_4
XANTENNA__23729__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16492_ _16471_/X _16423_/B VGND VGND VPWR VPWR _16494_/B sky130_fd_sc_hd__or2_4
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18231_ _16978_/B VGND VGND VPWR VPWR _18231_/Y sky130_fd_sc_hd__inv_2
X_15443_ _15443_/A _23084_/Q VGND VGND VPWR VPWR _15443_/X sky130_fd_sc_hd__or2_4
X_12655_ _12655_/A _12649_/X _12654_/X VGND VGND VPWR VPWR _12655_/X sky130_fd_sc_hd__or3_4
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ _11606_/A VGND VGND VPWR VPWR _15015_/A sky130_fd_sc_hd__buf_2
X_18162_ _18134_/X _18140_/Y _18148_/X _18159_/X _18161_/Y VGND VGND VPWR VPWR _18162_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _12567_/A _15300_/B VGND VGND VPWR VPWR _15375_/C sky130_fd_sc_hd__or2_4
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _12981_/A _12586_/B VGND VGND VPWR VPWR _12587_/C sky130_fd_sc_hd__or2_4
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17113_ _17322_/B VGND VGND VPWR VPWR _17114_/A sky130_fd_sc_hd__inv_2
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _15571_/A _14323_/X _14325_/C VGND VGND VPWR VPWR _14325_/X sky130_fd_sc_hd__and3_4
XFILLER_102_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11537_ _24422_/Q IRQ[7] _11536_/X VGND VGND VPWR VPWR _11538_/B sky130_fd_sc_hd__a21o_4
X_18093_ _16984_/X VGND VGND VPWR VPWR _18093_/Y sky130_fd_sc_hd__inv_2
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12933__A _12926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16405__A _13477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17044_ _17028_/X _17039_/X _17043_/X VGND VGND VPWR VPWR _17044_/Y sky130_fd_sc_hd__o21ai_4
X_14256_ _14218_/X _23625_/Q VGND VGND VPWR VPWR _14257_/C sky130_fd_sc_hd__or2_4
X_13207_ _13228_/A _13140_/B VGND VGND VPWR VPWR _13210_/B sky130_fd_sc_hd__or2_4
XANTENNA__18825__A1 _17277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22082__B1 _16708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14187_ _14218_/A VGND VGND VPWR VPWR _14205_/A sky130_fd_sc_hd__buf_2
XFILLER_67_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13138_ _12691_/A _13138_/B VGND VGND VPWR VPWR _13139_/C sky130_fd_sc_hd__or2_4
X_18995_ _11524_/A VGND VGND VPWR VPWR _18995_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13764__A _12937_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13069_ _13104_/A _13069_/B VGND VGND VPWR VPWR _13071_/B sky130_fd_sc_hd__or2_4
X_17946_ _17946_/A _17946_/B VGND VGND VPWR VPWR _17946_/X sky130_fd_sc_hd__and2_4
XFILLER_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21188__A2 _21183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21981__A _21988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17877_ _18180_/A VGND VGND VPWR VPWR _18390_/A sky130_fd_sc_hd__buf_2
XFILLER_93_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20935__A2 _20873_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19616_ _19450_/A VGND VGND VPWR VPWR _19616_/X sky130_fd_sc_hd__buf_2
XANTENNA__14298__C _14298_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19451__A HRDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16828_ _12434_/X _16827_/X _12434_/X _16827_/X VGND VGND VPWR VPWR _16889_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19547_ _19534_/X _19537_/Y _19543_/X _19445_/X _19546_/Y VGND VGND VPWR VPWR _19547_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20988__A1_N _19769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16759_ _16773_/A _16759_/B VGND VGND VPWR VPWR _16760_/C sky130_fd_sc_hd__or2_4
XANTENNA__22688__A2 _22686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18067__A _18267_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19478_ _19598_/A _19541_/A VGND VGND VPWR VPWR _19481_/B sky130_fd_sc_hd__or2_4
XFILLER_34_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12827__B _12827_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18429_ _18428_/A _18427_/X _18048_/X VGND VGND VPWR VPWR _18429_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13004__A _13004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19404__A2_N _18598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21440_ _21400_/A VGND VGND VPWR VPWR _21440_/X sky130_fd_sc_hd__buf_2
XFILLER_30_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21221__A _21791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21371_ _21249_/X _21369_/X _13123_/B _21366_/X VGND VGND VPWR VPWR _23858_/D sky130_fd_sc_hd__o22a_4
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16315__A _16188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12843__A _12752_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24360__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20322_ _20494_/A VGND VGND VPWR VPWR _20322_/X sky130_fd_sc_hd__buf_2
X_23110_ _23494_/CLK _23110_/D VGND VGND VPWR VPWR _14308_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20871__A1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24090_ _23472_/CLK _20375_/X VGND VGND VPWR VPWR _24090_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20871__B2 _20839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16034__B _15969_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20253_ _20473_/A VGND VGND VPWR VPWR _20253_/X sky130_fd_sc_hd__buf_2
X_23041_ _23041_/A VGND VGND VPWR VPWR HADDR[27] sky130_fd_sc_hd__inv_2
XANTENNA__22612__A2 _22607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20184_ _24447_/Q VGND VGND VPWR VPWR _20184_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22052__A _22052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13674__A _15442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22376__B2 _22372_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21891__A _21884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23943_ _23591_/CLK _21200_/X VGND VGND VPWR VPWR _23943_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24184__CLK _24162_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16985__A _16985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23874_ _23812_/CLK _23874_/D VGND VGND VPWR VPWR _15282_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22128__B2 _22120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22825_ _22824_/X VGND VGND VPWR VPWR _22825_/X sky130_fd_sc_hd__buf_2
XFILLER_77_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11922__A _11921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22756_ _22756_/A _22755_/B VGND VGND VPWR VPWR _22756_/Y sky130_fd_sc_hd__nand2_4
X_21707_ _21534_/X _21705_/X _23666_/Q _21702_/X VGND VGND VPWR VPWR _21707_/X sky130_fd_sc_hd__o22a_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15113__B _23615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22687_ _21246_/A _22686_/X _23091_/Q _22683_/X VGND VGND VPWR VPWR _22687_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18705__A _17117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12440_ _15392_/A VGND VGND VPWR VPWR _12441_/A sky130_fd_sc_hd__buf_2
X_24426_ _24365_/CLK _18797_/X HRESETn VGND VGND VPWR VPWR _24426_/Q sky130_fd_sc_hd__dfrtp_4
X_21638_ _21637_/X VGND VGND VPWR VPWR _21638_/X sky130_fd_sc_hd__buf_2
XFILLER_90_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24109__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18504__B1 _17878_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12371_ _13256_/A VGND VGND VPWR VPWR _12418_/A sky130_fd_sc_hd__buf_2
X_24357_ _24320_/CLK _24357_/D HRESETn VGND VGND VPWR VPWR _19079_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__13592__A2 _13591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20311__B1 _20310_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21569_ _21567_/X _21568_/X _14662_/B _21563_/X VGND VGND VPWR VPWR _23748_/D sky130_fd_sc_hd__o22a_4
XFILLER_20_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12753__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14110_ _14994_/A VGND VGND VPWR VPWR _14117_/A sky130_fd_sc_hd__buf_2
XFILLER_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23308_ _23794_/CLK _22318_/X VGND VGND VPWR VPWR _23308_/Q sky130_fd_sc_hd__dfxtp_4
X_15090_ _15109_/A _23583_/Q VGND VGND VPWR VPWR _15090_/X sky130_fd_sc_hd__or2_4
XANTENNA__13568__B _13568_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24288_ _24290_/CLK _19200_/X HRESETn VGND VGND VPWR VPWR _24288_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14041_ _14813_/A _23882_/Q VGND VGND VPWR VPWR _14041_/X sky130_fd_sc_hd__or2_4
XFILLER_10_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22064__B1 _23456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23239_ _23079_/CLK _22445_/X VGND VGND VPWR VPWR _13841_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__18807__A1 _15379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19536__A _19536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22603__A2 _22600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18440__A _18204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23058__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17800_ _17800_/A VGND VGND VPWR VPWR _17800_/X sky130_fd_sc_hd__buf_2
X_15992_ _16096_/A _15992_/B VGND VGND VPWR VPWR _15992_/X sky130_fd_sc_hd__or2_4
X_18780_ _12674_/X _18774_/X _20470_/A _18775_/X VGND VGND VPWR VPWR _18780_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22367__B2 _22365_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14943_ _11642_/A _14943_/B _14942_/X VGND VGND VPWR VPWR _14943_/X sky130_fd_sc_hd__and3_4
X_17731_ _17744_/A VGND VGND VPWR VPWR _17731_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21009__C _21162_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14874_ _14991_/A _14872_/X _14873_/X VGND VGND VPWR VPWR _14874_/X sky130_fd_sc_hd__and3_4
X_17662_ _24131_/Q _17662_/B VGND VGND VPWR VPWR _17662_/X sky130_fd_sc_hd__or2_4
XFILLER_97_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19401_ _19399_/X _18536_/Y _19399_/X _24200_/Q VGND VGND VPWR VPWR _19401_/X sky130_fd_sc_hd__a2bb2o_4
X_13825_ _13636_/A _13825_/B VGND VGND VPWR VPWR _13826_/C sky130_fd_sc_hd__or2_4
X_16613_ _11746_/X VGND VGND VPWR VPWR _16622_/A sky130_fd_sc_hd__buf_2
X_17593_ _17377_/X _17592_/X _17371_/X _17380_/B VGND VGND VPWR VPWR _17594_/A sky130_fd_sc_hd__a211o_4
XFILLER_95_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12928__A _12591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11832__A _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16544_ _11886_/X VGND VGND VPWR VPWR _16586_/A sky130_fd_sc_hd__buf_2
X_19332_ _19328_/A VGND VGND VPWR VPWR _19332_/X sky130_fd_sc_hd__buf_2
XANTENNA__15304__A _15030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21878__B1 _16405_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13756_ _15493_/A _13756_/B VGND VGND VPWR VPWR _13756_/X sky130_fd_sc_hd__or2_4
XFILLER_91_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17546__A1 _17542_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17546__B2 _17646_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21342__A2 _21340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16119__B _16189_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12707_ _12235_/A _23924_/Q VGND VGND VPWR VPWR _12707_/X sky130_fd_sc_hd__or2_4
XANTENNA__11551__B IRQ[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16475_ _16499_/A _16475_/B _16475_/C VGND VGND VPWR VPWR _16475_/X sky130_fd_sc_hd__and3_4
X_19263_ _19263_/A VGND VGND VPWR VPWR _19263_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15023__B _15023_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13687_ _13884_/A VGND VGND VPWR VPWR _13754_/A sky130_fd_sc_hd__buf_2
X_15426_ _15430_/A _15490_/B VGND VGND VPWR VPWR _15427_/C sky130_fd_sc_hd__or2_4
X_18214_ _17871_/A _18213_/Y VGND VGND VPWR VPWR _18214_/X sky130_fd_sc_hd__and2_4
XFILLER_31_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12638_ _12638_/A VGND VGND VPWR VPWR _12982_/A sky130_fd_sc_hd__buf_2
X_19194_ _19112_/A _19112_/B _19193_/Y VGND VGND VPWR VPWR _19194_/X sky130_fd_sc_hd__o21a_4
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22137__A _22125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21041__A _21027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15357_ _15325_/X _15355_/X _15357_/C VGND VGND VPWR VPWR _15361_/B sky130_fd_sc_hd__and3_4
X_18145_ _17864_/X _18143_/X _17823_/X _18144_/X VGND VGND VPWR VPWR _18145_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17849__A2 _17847_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13759__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12569_ _13718_/A VGND VGND VPWR VPWR _15487_/A sky130_fd_sc_hd__buf_2
XANTENNA__12663__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16135__A _16139_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14308_ _15552_/A _14308_/B VGND VGND VPWR VPWR _14308_/X sky130_fd_sc_hd__or2_4
XFILLER_117_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18076_ _17933_/A VGND VGND VPWR VPWR _18076_/X sky130_fd_sc_hd__buf_2
X_15288_ _14146_/X _15288_/B _15287_/X VGND VGND VPWR VPWR _15288_/X sky130_fd_sc_hd__or3_4
X_17027_ _17457_/B VGND VGND VPWR VPWR _17561_/B sky130_fd_sc_hd__buf_2
X_14239_ _14251_/A _23369_/Q VGND VGND VPWR VPWR _14239_/X sky130_fd_sc_hd__or2_4
XANTENNA__15974__A _15939_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19446__A _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16789__B _23835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13494__A _12655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18978_ _11527_/A _11526_/X _18973_/Y VGND VGND VPWR VPWR _18978_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_67_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17929_ _17914_/X _17925_/X _17926_/X _17928_/Y VGND VGND VPWR VPWR _17929_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22600__A _22600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20940_ _20875_/A _20754_/A VGND VGND VPWR VPWR _20940_/X sky130_fd_sc_hd__or2_4
XFILLER_66_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20871_ _20750_/X _20870_/X _14477_/B _20839_/X VGND VGND VPWR VPWR _20871_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22610_ _22456_/X _22607_/X _15276_/B _22604_/X VGND VGND VPWR VPWR _23138_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11742__A _11741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23590_ _23781_/CLK _21849_/X VGND VGND VPWR VPWR _14304_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_74_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6_0_HCLK_A clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22541_ _22422_/X _22536_/X _13291_/B _22540_/X VGND VGND VPWR VPWR _22541_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20541__B1 _24434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18525__A _18137_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22472_ _22486_/A VGND VGND VPWR VPWR _22472_/X sky130_fd_sc_hd__buf_2
XANTENNA__15868__B _15799_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24211_ _23522_/CLK _24211_/D HRESETn VGND VGND VPWR VPWR _24211_/Q sky130_fd_sc_hd__dfrtp_4
X_21423_ _21416_/A VGND VGND VPWR VPWR _21423_/X sky130_fd_sc_hd__buf_2
XANTENNA__13669__A _13636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21097__B2 _21093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12573__A _13708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16045__A _16045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19358__A2_N _18723_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24142_ _24230_/CLK _24142_/D HRESETn VGND VGND VPWR VPWR _24142_/Q sky130_fd_sc_hd__dfrtp_4
X_21354_ _21383_/A VGND VGND VPWR VPWR _21369_/A sky130_fd_sc_hd__buf_2
XFILLER_108_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20305_ _20242_/X VGND VGND VPWR VPWR _20305_/X sky130_fd_sc_hd__buf_2
XANTENNA__15884__A _15884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22046__B1 _15769_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24073_ _23910_/CLK _24073_/D VGND VGND VPWR VPWR _24073_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21285_ _21855_/A VGND VGND VPWR VPWR _21285_/X sky130_fd_sc_hd__buf_2
XFILLER_104_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23024_ _23014_/X _16985_/A _22997_/X _23023_/X VGND VGND VPWR VPWR _23025_/A sky130_fd_sc_hd__a211o_4
XFILLER_104_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20236_ _20467_/A VGND VGND VPWR VPWR _20424_/A sky130_fd_sc_hd__buf_2
XFILLER_115_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20167_ _24444_/Q IRQ[29] _20166_/X VGND VGND VPWR VPWR _20168_/B sky130_fd_sc_hd__a21boi_4
XANTENNA__23574__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20098_ _20086_/A _20098_/B VGND VGND VPWR VPWR _20098_/X sky130_fd_sc_hd__or2_4
X_11940_ _11995_/A _11940_/B _11940_/C VGND VGND VPWR VPWR _11947_/B sky130_fd_sc_hd__and3_4
X_23926_ _23473_/CLK _23926_/D VGND VGND VPWR VPWR _12270_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21021__B2 _21020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_23_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR _24165_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14947__B _14873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21126__A _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_86_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR _23358_/CLK sky130_fd_sc_hd__clkbuf_1
X_11871_ _13014_/A VGND VGND VPWR VPWR _12493_/A sky130_fd_sc_hd__buf_2
X_23857_ _23342_/CLK _23857_/D VGND VGND VPWR VPWR _13257_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12748__A _13004_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13610_ _12216_/A VGND VGND VPWR VPWR _13611_/A sky130_fd_sc_hd__buf_2
XANTENNA__11652__A _15611_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22808_ _14074_/A _22794_/X _22796_/X _22807_/X VGND VGND VPWR VPWR _22809_/B sky130_fd_sc_hd__o22a_4
X_14590_ _14725_/A _14679_/B VGND VGND VPWR VPWR _14590_/X sky130_fd_sc_hd__or2_4
XFILLER_38_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23788_ _23698_/CLK _21480_/X VGND VGND VPWR VPWR _23788_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21324__A2 _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13541_ _12413_/X _13539_/X _13540_/X VGND VGND VPWR VPWR _13541_/X sky130_fd_sc_hd__and3_4
X_22739_ _22738_/Y _24100_/Q _22738_/Y _24100_/Q VGND VGND VPWR VPWR _22746_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18435__A _18381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16260_ _15934_/X _16260_/B VGND VGND VPWR VPWR _16260_/X sky130_fd_sc_hd__or2_4
XFILLER_13_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13472_ _13448_/X _13552_/B VGND VGND VPWR VPWR _13474_/B sky130_fd_sc_hd__or2_4
XFILLER_90_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15211_ _14183_/A _15208_/X _15210_/X VGND VGND VPWR VPWR _15211_/X sky130_fd_sc_hd__and3_4
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12423_ _12384_/X _12323_/B VGND VGND VPWR VPWR _12423_/X sky130_fd_sc_hd__or2_4
X_24409_ _24435_/CLK _18829_/X HRESETn VGND VGND VPWR VPWR _24409_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13579__A _13350_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16191_ _16229_/A _16183_/X _16190_/X VGND VGND VPWR VPWR _16199_/B sky130_fd_sc_hd__or3_4
XANTENNA__21088__B2 _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15142_ _15142_/A _15212_/B VGND VGND VPWR VPWR _15144_/B sky130_fd_sc_hd__or2_4
X_12354_ _11680_/X _12354_/B _12353_/X VGND VGND VPWR VPWR _12354_/X sky130_fd_sc_hd__or3_4
XFILLER_86_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15073_ _15109_/A _23135_/Q VGND VGND VPWR VPWR _15076_/B sky130_fd_sc_hd__or2_4
X_19950_ _17989_/X _17047_/A _19949_/X _17874_/X _18747_/X VGND VGND VPWR VPWR _19950_/X
+ sky130_fd_sc_hd__a32o_4
X_12285_ _12284_/X _12285_/B VGND VGND VPWR VPWR _12288_/B sky130_fd_sc_hd__or2_4
XFILLER_101_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14024_ _12598_/A VGND VGND VPWR VPWR _14046_/A sky130_fd_sc_hd__buf_2
X_18901_ _15780_/B _18898_/X _24366_/Q _18899_/X VGND VGND VPWR VPWR _24366_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22588__B2 _22583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19881_ _19881_/A _19881_/B VGND VGND VPWR VPWR _19881_/X sky130_fd_sc_hd__or2_4
XFILLER_49_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19453__A1 _20224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19453__B2 HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18832_ _12430_/X _18827_/X _24406_/Q _18828_/X VGND VGND VPWR VPWR _18832_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21260__B2 _21254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14203__A _11738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18763_ _18762_/X VGND VGND VPWR VPWR _18788_/A sky130_fd_sc_hd__buf_2
XANTENNA__23001__A2 _17667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15975_ _15952_/A _23960_/Q VGND VGND VPWR VPWR _15976_/C sky130_fd_sc_hd__or2_4
XFILLER_48_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22420__A _20573_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17714_ _17712_/X _17713_/X VGND VGND VPWR VPWR _17714_/X sky130_fd_sc_hd__or2_4
XFILLER_48_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14926_ _13992_/A _14926_/B _14926_/C VGND VGND VPWR VPWR _14935_/B sky130_fd_sc_hd__or3_4
XFILLER_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18694_ _18327_/A _17853_/Y VGND VGND VPWR VPWR _18694_/X sky130_fd_sc_hd__and2_4
XFILLER_64_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14857__B _14857_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18329__B _18274_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17645_ _17645_/A _17535_/Y VGND VGND VPWR VPWR _17648_/A sky130_fd_sc_hd__and2_4
XFILLER_36_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14857_ _12472_/A _14857_/B VGND VGND VPWR VPWR _14857_/X sky130_fd_sc_hd__or2_4
XFILLER_21_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11562__A _20558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15034__A _13927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13808_ _13620_/A _23943_/Q VGND VGND VPWR VPWR _13808_/X sky130_fd_sc_hd__or2_4
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14788_ _13851_/A _14788_/B VGND VGND VPWR VPWR _14789_/C sky130_fd_sc_hd__or2_4
X_17576_ _17144_/Y _17570_/Y _17569_/A _17575_/X VGND VGND VPWR VPWR _17576_/X sky130_fd_sc_hd__o22a_4
XFILLER_63_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21315__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22512__B2 _22476_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19315_ _19313_/X _17884_/X _19313_/X _24252_/Q VGND VGND VPWR VPWR _24252_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13739_ _12612_/A _13731_/X _13739_/C VGND VGND VPWR VPWR _13740_/C sky130_fd_sc_hd__and3_4
X_16527_ _16538_/A _16602_/B VGND VGND VPWR VPWR _16527_/X sky130_fd_sc_hd__or2_4
XANTENNA__15969__A _15997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19246_ _19230_/A _19247_/A _19245_/Y VGND VGND VPWR VPWR _24281_/D sky130_fd_sc_hd__o21a_4
X_16458_ _12837_/A VGND VGND VPWR VPWR _16499_/A sky130_fd_sc_hd__buf_2
X_15409_ _15432_/A _23308_/Q VGND VGND VPWR VPWR _15409_/X sky130_fd_sc_hd__or2_4
X_16389_ _11915_/A _16387_/X _16389_/C VGND VGND VPWR VPWR _16389_/X sky130_fd_sc_hd__and3_4
X_19177_ _19177_/A VGND VGND VPWR VPWR _19177_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12393__A _12826_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18128_ _18056_/X _18127_/X _19990_/A _18056_/X VGND VGND VPWR VPWR _24471_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18059_ _18012_/X _16985_/X _18017_/Y VGND VGND VPWR VPWR _23027_/B sky130_fd_sc_hd__a21oi_4
X_21070_ _20339_/X _21068_/X _24028_/Q _21065_/X VGND VGND VPWR VPWR _24028_/D sky130_fd_sc_hd__o22a_4
XFILLER_63_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20021_ _18312_/X _20009_/X _20019_/Y _20020_/X VGND VGND VPWR VPWR _20021_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15209__A _11708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14113__A _14113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21003__A1 _20511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21003__B2 _20202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17424__A _13920_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21972_ _21966_/Y _21971_/X _21789_/X _21971_/X VGND VGND VPWR VPWR _23518_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13492__A1 _11980_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21554__A2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23711_ _23217_/CLK _23711_/D VGND VGND VPWR VPWR _23711_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20923_ _20922_/Y _20851_/X _20539_/B _20675_/X VGND VGND VPWR VPWR _20923_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12568__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24454__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ _23706_/CLK _23642_/D VGND VGND VPWR VPWR _16508_/B sky130_fd_sc_hd__dfxtp_4
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20854_ _20854_/A _20556_/A VGND VGND VPWR VPWR _20854_/Y sky130_fd_sc_hd__nand2_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21306__A2 _21305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12287__B _12287_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22503__B2 _22497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23573_ _23315_/CLK _21885_/X VGND VGND VPWR VPWR _12505_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20785_ _24392_/Q _20623_/X _24424_/Q _20682_/X VGND VGND VPWR VPWR _20785_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14783__A _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22524_ _22394_/X _22522_/X _16614_/B _22519_/X VGND VGND VPWR VPWR _22524_/X sky130_fd_sc_hd__o22a_4
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23059__A2 _19306_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15598__B _23915_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22267__B1 _16092_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22455_ _22454_/X _22452_/X _14787_/B _22447_/X VGND VGND VPWR VPWR _23235_/D sky130_fd_sc_hd__o22a_4
XFILLER_13_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20817__A1 _24199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21406_ _21221_/X _21405_/X _23837_/Q _21402_/X VGND VGND VPWR VPWR _21406_/X sky130_fd_sc_hd__o22a_4
XFILLER_41_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22386_ _22423_/A VGND VGND VPWR VPWR _22386_/X sky130_fd_sc_hd__buf_2
XFILLER_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24125_ _24126_/CLK _20032_/Y HRESETn VGND VGND VPWR VPWR _16951_/A sky130_fd_sc_hd__dfrtp_4
X_21337_ _21316_/A VGND VGND VPWR VPWR _21337_/X sky130_fd_sc_hd__buf_2
XANTENNA__21490__B2 _21488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12070_ _11971_/A VGND VGND VPWR VPWR _12098_/A sky130_fd_sc_hd__buf_2
X_24056_ _23316_/CLK _21024_/X VGND VGND VPWR VPWR _24056_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_46_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21268_ _20748_/A VGND VGND VPWR VPWR _21268_/X sky130_fd_sc_hd__buf_2
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23007_ _23006_/X VGND VGND VPWR VPWR HADDR[21] sky130_fd_sc_hd__inv_2
XANTENNA__11647__A _11647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20219_ _24158_/Q VGND VGND VPWR VPWR _20846_/B sky130_fd_sc_hd__buf_2
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21199_ _20797_/X _21197_/X _13652_/B _21194_/X VGND VGND VPWR VPWR _21199_/X sky130_fd_sc_hd__o22a_4
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14023__A _14815_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22240__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13862__A _13862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19865__A2_N _19864_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15760_ _11680_/X _15760_/B _15759_/X VGND VGND VPWR VPWR _15760_/X sky130_fd_sc_hd__or3_4
XFILLER_111_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12972_ _13118_/A _12972_/B _12971_/X VGND VGND VPWR VPWR _12988_/B sky130_fd_sc_hd__and3_4
XFILLER_18_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21545__A2 _21544_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22742__A1 SYSTICKCLKDIV[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11923_ _11995_/A _11923_/B _11923_/C VGND VGND VPWR VPWR _11923_/X sky130_fd_sc_hd__and3_4
X_14711_ _14714_/A _24068_/Q VGND VGND VPWR VPWR _14712_/C sky130_fd_sc_hd__or2_4
XFILLER_46_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15691_ _15664_/A _15691_/B _15691_/C VGND VGND VPWR VPWR _15695_/B sky130_fd_sc_hd__and3_4
X_23909_ _23973_/CLK _21281_/X VGND VGND VPWR VPWR _14453_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12478__A _12477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14642_ _14642_/A VGND VGND VPWR VPWR _15108_/A sky130_fd_sc_hd__buf_2
X_17430_ _17382_/X _17429_/X VGND VGND VPWR VPWR _17430_/Y sky130_fd_sc_hd__nor2_4
X_11854_ _11853_/X VGND VGND VPWR VPWR _16741_/A sky130_fd_sc_hd__buf_2
XANTENNA__24124__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14573_ _15019_/A VGND VGND VPWR VPWR _15142_/A sky130_fd_sc_hd__buf_2
X_17361_ _17361_/A _17360_/Y VGND VGND VPWR VPWR _17361_/X sky130_fd_sc_hd__or2_4
XANTENNA__15789__A _12859_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11785_ _11691_/X VGND VGND VPWR VPWR _12169_/A sky130_fd_sc_hd__buf_2
XFILLER_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20505__B1 _20504_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19100_ _19087_/X _19099_/X _18971_/A _11503_/A VGND VGND VPWR VPWR _24321_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13524_ _13561_/A _13456_/B VGND VGND VPWR VPWR _13527_/B sky130_fd_sc_hd__or2_4
X_16312_ _16366_/A _16309_/X _16311_/X VGND VGND VPWR VPWR _16312_/X sky130_fd_sc_hd__and3_4
XFILLER_53_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17292_ _17294_/B VGND VGND VPWR VPWR _17295_/B sky130_fd_sc_hd__inv_2
X_16243_ _16090_/A VGND VGND VPWR VPWR _16243_/X sky130_fd_sc_hd__buf_2
X_19031_ _24333_/Q VGND VGND VPWR VPWR _19031_/Y sky130_fd_sc_hd__inv_2
X_13455_ _12464_/A _13453_/X _13454_/X VGND VGND VPWR VPWR _13455_/X sky130_fd_sc_hd__and3_4
XFILLER_31_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12406_ _15889_/A _12406_/B _12405_/X VGND VGND VPWR VPWR _12406_/X sky130_fd_sc_hd__or3_4
XANTENNA__13102__A _13102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16174_ _13376_/X VGND VGND VPWR VPWR _16223_/A sky130_fd_sc_hd__buf_2
X_13386_ _13376_/X _13304_/B VGND VGND VPWR VPWR _13388_/B sky130_fd_sc_hd__or2_4
XANTENNA__22415__A _22100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15125_ _12202_/A _15125_/B VGND VGND VPWR VPWR _15125_/X sky130_fd_sc_hd__or2_4
X_12337_ _12189_/X _11618_/A _12280_/X _12281_/X _12336_/X VGND VGND VPWR VPWR _12338_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16413__A _15999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12941__A _13083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15056_ _15069_/A _15056_/B VGND VGND VPWR VPWR _15058_/B sky130_fd_sc_hd__or2_4
X_19933_ _19933_/A VGND VGND VPWR VPWR _20000_/A sky130_fd_sc_hd__buf_2
X_12268_ _12267_/X VGND VGND VPWR VPWR _12269_/A sky130_fd_sc_hd__buf_2
XANTENNA__19426__A1 HRDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19426__B2 _19416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12660__B _12660_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14007_ _11738_/A VGND VGND VPWR VPWR _14008_/A sky130_fd_sc_hd__buf_2
XANTENNA__15029__A _15006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21233__B2 _21230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19864_ _19445_/X _19863_/X _19494_/X _19775_/Y VGND VGND VPWR VPWR _19864_/X sky130_fd_sc_hd__o22a_4
XFILLER_96_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12199_ _12198_/X VGND VGND VPWR VPWR _15654_/A sky130_fd_sc_hd__buf_2
X_18815_ _18762_/A _18814_/X VGND VGND VPWR VPWR _18815_/X sky130_fd_sc_hd__or2_4
XFILLER_116_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19795_ _19524_/B _19794_/X _19872_/C VGND VGND VPWR VPWR _19795_/X sky130_fd_sc_hd__o21a_4
XFILLER_7_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22150__A _21583_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13772__A _11656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18746_ _18746_/A VGND VGND VPWR VPWR _18746_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24245__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15958_ _15994_/A _15958_/B _15958_/C VGND VGND VPWR VPWR _15963_/B sky130_fd_sc_hd__and3_4
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19375__A1_N _19374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14909_ _14912_/A _14909_/B VGND VGND VPWR VPWR _14909_/X sky130_fd_sc_hd__or2_4
X_18677_ _17323_/X _18675_/X _17779_/X _18676_/X VGND VGND VPWR VPWR _18677_/X sky130_fd_sc_hd__a211o_4
X_15889_ _15889_/A _15889_/B _15889_/C VGND VGND VPWR VPWR _15889_/X sky130_fd_sc_hd__or3_4
XANTENNA__16412__A1 _11852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17628_ _17628_/A _17582_/X _17628_/C VGND VGND VPWR VPWR _17629_/A sky130_fd_sc_hd__and3_4
XFILLER_24_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12029__A2 _11619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15699__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17559_ _17559_/A VGND VGND VPWR VPWR _18085_/A sky130_fd_sc_hd__inv_2
XFILLER_20_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20570_ _24241_/Q _20421_/X _20569_/X VGND VGND VPWR VPWR _20570_/X sky130_fd_sc_hd__o21a_4
XFILLER_108_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19229_ _24280_/Q _19249_/A VGND VGND VPWR VPWR _19247_/A sky130_fd_sc_hd__and2_4
XANTENNA__13012__A _13031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22240_ _22219_/A VGND VGND VPWR VPWR _22240_/X sky130_fd_sc_hd__buf_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13947__A _12217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22171_ _22098_/X _22165_/X _12819_/B _22169_/X VGND VGND VPWR VPWR _23412_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21472__B2 _21467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21122_ _20356_/X _21119_/X _23995_/Q _21116_/X VGND VGND VPWR VPWR _23995_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20027__A2 _17681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21224__A1 _21221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21053_ _20916_/X _21051_/X _14759_/B _21048_/X VGND VGND VPWR VPWR _21053_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19968__A2 _17769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21224__B2 _21218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21775__A2 _21769_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20004_ _20003_/X VGND VGND VPWR VPWR _20004_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16977__B _16977_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14778__A _14778_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20983__B1 _14903_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13682__A _13682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22724__A1 _19497_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21955_ _21845_/X _21952_/X _23527_/Q _21949_/X VGND VGND VPWR VPWR _21955_/X sky130_fd_sc_hd__o22a_4
XFILLER_41_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12298__A _15667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _20760_/X _20905_/X _24323_/Q _20767_/X VGND VGND VPWR VPWR _20906_/X sky130_fd_sc_hd__o22a_4
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21886_ _21814_/X _21880_/X _23572_/Q _21884_/X VGND VGND VPWR VPWR _21886_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23625_ _23336_/CLK _21770_/X VGND VGND VPWR VPWR _23625_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _22446_/A VGND VGND VPWR VPWR _20838_/A sky130_fd_sc_hd__buf_2
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11930__A _13813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23762__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15402__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _20297_/A IRQ[30] VGND VGND VPWR VPWR _11570_/X sky130_fd_sc_hd__and2_4
X_23556_ _23433_/CLK _23556_/D VGND VGND VPWR VPWR _23556_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20768_ _20760_/X _20766_/X _24329_/Q _20767_/X VGND VGND VPWR VPWR _20768_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21160__B1 _15079_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12745__B _12827_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22507_ _22471_/A VGND VGND VPWR VPWR _22507_/X sky130_fd_sc_hd__buf_2
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23487_ _23487_/CLK _23487_/D VGND VGND VPWR VPWR _23487_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20699_ HRDATA[12] _20699_/B VGND VGND VPWR VPWR _20699_/X sky130_fd_sc_hd__or2_4
XFILLER_52_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18713__A _18713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14018__A _14847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ _13214_/A _13240_/B _13240_/C VGND VGND VPWR VPWR _13240_/X sky130_fd_sc_hd__and3_4
XFILLER_108_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22438_ _22437_/X _22428_/X _13995_/B _22435_/X VGND VGND VPWR VPWR _23242_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24118__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13171_ _15689_/A _13171_/B VGND VGND VPWR VPWR _13171_/X sky130_fd_sc_hd__or2_4
XANTENNA__17329__A _15121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22369_ _22124_/X _22368_/X _23273_/Q _22365_/X VGND VGND VPWR VPWR _23273_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12761__A _13130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12122_ _16071_/A VGND VGND VPWR VPWR _12167_/A sky130_fd_sc_hd__buf_2
X_24108_ _24293_/CLK _24108_/D HRESETn VGND VGND VPWR VPWR _19108_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12053_ _16698_/A _23773_/Q VGND VGND VPWR VPWR _12054_/C sky130_fd_sc_hd__or2_4
X_16930_ _17024_/C _16929_/X VGND VGND VPWR VPWR _17062_/A sky130_fd_sc_hd__or2_4
X_24039_ _23591_/CLK _21047_/X VGND VGND VPWR VPWR _24039_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19959__A2 _19306_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19544__A HRDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16861_ _14724_/X _16860_/X _14724_/X _16860_/X VGND VGND VPWR VPWR _16861_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15791__B _15852_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14688__A _15105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18600_ _17639_/A _18576_/X _16927_/A _18599_/X VGND VGND VPWR VPWR _18600_/X sky130_fd_sc_hd__o22a_4
X_15812_ _15812_/A _15812_/B VGND VGND VPWR VPWR _15812_/X sky130_fd_sc_hd__and2_4
XANTENNA__24337__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19580_ _19839_/A VGND VGND VPWR VPWR _19580_/X sky130_fd_sc_hd__buf_2
XFILLER_115_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16792_ _16768_/X _16792_/B VGND VGND VPWR VPWR _16793_/C sky130_fd_sc_hd__or2_4
XFILLER_111_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24305__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21518__A2 _21508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18531_ _18480_/X _18529_/X _18508_/X _18530_/X VGND VGND VPWR VPWR _18531_/X sky130_fd_sc_hd__o22a_4
XFILLER_98_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12955_ _12955_/A _12951_/X _12954_/X VGND VGND VPWR VPWR _12956_/C sky130_fd_sc_hd__or3_4
X_15743_ _15743_/A _15741_/X _15743_/C VGND VGND VPWR VPWR _15743_/X sky130_fd_sc_hd__and3_4
XFILLER_34_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22191__A2 _22186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11906_ _11905_/Y VGND VGND VPWR VPWR _12250_/A sky130_fd_sc_hd__buf_2
XFILLER_94_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18462_ _18097_/A _18351_/B _18459_/Y _18016_/A _22949_/B VGND VGND VPWR VPWR _18463_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_34_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12886_ _12886_/A _12943_/B VGND VGND VPWR VPWR _12886_/X sky130_fd_sc_hd__or2_4
X_15674_ _12240_/A _15674_/B VGND VGND VPWR VPWR _15675_/C sky130_fd_sc_hd__or2_4
XANTENNA__12001__A _11997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_56_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17413_ _17413_/A _17413_/B VGND VGND VPWR VPWR _17413_/X sky130_fd_sc_hd__or2_4
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11837_ _16077_/A _11837_/B _11837_/C VGND VGND VPWR VPWR _11837_/X sky130_fd_sc_hd__and3_4
X_14625_ _14763_/A _24068_/Q VGND VGND VPWR VPWR _14625_/X sky130_fd_sc_hd__or2_4
XFILLER_92_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18393_ _17968_/X _18367_/Y _17933_/X _18392_/Y VGND VGND VPWR VPWR _18393_/X sky130_fd_sc_hd__a211o_4
XFILLER_18_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14556_ _14556_/A _14554_/X _14555_/X VGND VGND VPWR VPWR _14556_/X sky130_fd_sc_hd__and3_4
X_17344_ _17125_/Y _17344_/B VGND VGND VPWR VPWR _17365_/A sky130_fd_sc_hd__nor2_4
X_11768_ _15484_/A VGND VGND VPWR VPWR _13102_/A sky130_fd_sc_hd__buf_2
XANTENNA__19895__A1 _19884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ _12964_/A VGND VGND VPWR VPWR _13507_/X sky130_fd_sc_hd__buf_2
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14487_ _13623_/A _14487_/B VGND VGND VPWR VPWR _14487_/X sky130_fd_sc_hd__or2_4
X_17275_ _17272_/Y _17016_/X _17023_/X _17274_/Y VGND VGND VPWR VPWR _17275_/X sky130_fd_sc_hd__o22a_4
X_11699_ _13256_/A VGND VGND VPWR VPWR _12360_/A sky130_fd_sc_hd__buf_2
X_19014_ _24368_/Q VGND VGND VPWR VPWR _19014_/Y sky130_fd_sc_hd__inv_2
X_13438_ _13437_/X _13513_/B VGND VGND VPWR VPWR _13440_/B sky130_fd_sc_hd__or2_4
X_16226_ _16219_/A _16226_/B VGND VGND VPWR VPWR _16226_/X sky130_fd_sc_hd__or2_4
XANTENNA__22145__A _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16157_ _13395_/X VGND VGND VPWR VPWR _16158_/A sky130_fd_sc_hd__buf_2
XFILLER_31_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13767__A _12652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13369_ _13351_/X _13369_/B _13369_/C VGND VGND VPWR VPWR _13370_/C sky130_fd_sc_hd__and3_4
XANTENNA__21454__B2 _21453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17122__A2 _17105_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12671__A _13083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16143__A _16143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15108_ _15108_/A _15108_/B _15108_/C VGND VGND VPWR VPWR _15108_/X sky130_fd_sc_hd__or3_4
X_16088_ _16087_/X VGND VGND VPWR VPWR _16140_/A sky130_fd_sc_hd__buf_2
XFILLER_64_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15039_ _14752_/A _15039_/B _15039_/C VGND VGND VPWR VPWR _15039_/X sky130_fd_sc_hd__or3_4
X_19916_ _19909_/A VGND VGND VPWR VPWR _19916_/X sky130_fd_sc_hd__buf_2
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21206__B2 _21201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21757__A2 _21755_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16797__B _23803_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19847_ _19672_/C _19846_/X _19643_/A VGND VGND VPWR VPWR _19847_/X sky130_fd_sc_hd__o21a_4
XFILLER_60_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14598__A _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19778_ _19573_/A _19776_/X _19813_/A VGND VGND VPWR VPWR _19778_/X sky130_fd_sc_hd__o21a_4
XFILLER_42_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21509__A2 _21508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22706__B2 _22704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18729_ _17808_/X _18727_/X _18728_/X _17802_/X _17139_/X VGND VGND VPWR VPWR _18729_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_64_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22182__A2 _22179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21740_ _21740_/A VGND VGND VPWR VPWR _21755_/A sky130_fd_sc_hd__buf_2
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21671_ _21558_/X _21669_/X _13759_/B _21666_/X VGND VGND VPWR VPWR _23688_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12846__A _12435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23410_ _23314_/CLK _22174_/X VGND VGND VPWR VPWR _13039_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11750__A _11717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20622_ _20622_/A VGND VGND VPWR VPWR _20622_/X sky130_fd_sc_hd__buf_2
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24390_ _24365_/CLK _24390_/D HRESETn VGND VGND VPWR VPWR _24390_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21142__B1 _15799_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23341_ _23122_/CLK _22281_/X VGND VGND VPWR VPWR _15848_/B sky130_fd_sc_hd__dfxtp_4
X_20553_ _21249_/A VGND VGND VPWR VPWR _20553_/X sky130_fd_sc_hd__buf_2
XANTENNA__21693__B2 _21688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23272_ _23368_/CLK _23272_/D VGND VGND VPWR VPWR _23272_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15876__B _23885_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20484_ _20484_/A _20483_/X VGND VGND VPWR VPWR _20484_/X sky130_fd_sc_hd__or2_4
XANTENNA__14780__B _14780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22223_ _22100_/X _22222_/X _23379_/Q _22219_/X VGND VGND VPWR VPWR _22223_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21445__B2 _21401_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23165__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12581__A _14002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18310__B2 _18309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15124__A1 _14918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21996__A2 _21995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22154_ _22169_/A VGND VGND VPWR VPWR _22162_/A sky130_fd_sc_hd__buf_2
XFILLER_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21894__A _21887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21105_ _20916_/X _21103_/X _14797_/B _21100_/X VGND VGND VPWR VPWR _24003_/D sky130_fd_sc_hd__o22a_4
XFILLER_86_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15892__A _15892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22085_ _22083_/X _22077_/X _16408_/B _22084_/X VGND VGND VPWR VPWR _22085_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21036_ _20611_/X _21030_/X _13466_/B _21034_/X VGND VGND VPWR VPWR _24047_/D sky130_fd_sc_hd__o22a_4
XFILLER_47_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14301__A _12257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22987_ _22998_/A _22987_/B VGND VGND VPWR VPWR _22989_/B sky130_fd_sc_hd__or2_4
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22173__A2 _22172_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12740_ _12740_/A _12740_/B _12740_/C VGND VGND VPWR VPWR _12740_/X sky130_fd_sc_hd__and3_4
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21938_ _21938_/A VGND VGND VPWR VPWR _21938_/X sky130_fd_sc_hd__buf_2
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21381__B1 _15577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14955__B _23872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12671_ _13083_/A _12663_/X _12671_/C VGND VGND VPWR VPWR _12671_/X sky130_fd_sc_hd__and3_4
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ _21884_/A VGND VGND VPWR VPWR _21869_/X sky130_fd_sc_hd__buf_2
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _15633_/A _14410_/B VGND VGND VPWR VPWR _14411_/C sky130_fd_sc_hd__or2_4
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11622_/A _11621_/X VGND VGND VPWR VPWR _11622_/X sky130_fd_sc_hd__or2_4
X_23608_ _23539_/CLK _23608_/D VGND VGND VPWR VPWR _23608_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _14430_/X _14568_/Y _15388_/X _14430_/B _15389_/X VGND VGND VPWR VPWR _16840_/C
+ sky130_fd_sc_hd__o32a_4
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _14341_/A _14268_/B VGND VGND VPWR VPWR _14341_/X sky130_fd_sc_hd__or2_4
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _11550_/X _11552_/X VGND VGND VPWR VPWR _11553_/X sky130_fd_sc_hd__or2_4
X_23539_ _23539_/CLK _21939_/X VGND VGND VPWR VPWR _12953_/B sky130_fd_sc_hd__dfxtp_4
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18443__A _18443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17060_ _17024_/A VGND VGND VPWR VPWR _20194_/A sky130_fd_sc_hd__buf_2
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _12260_/X _14272_/B VGND VGND VPWR VPWR _14272_/X sky130_fd_sc_hd__or2_4
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16011_ _16039_/A _16009_/X _16011_/C VGND VGND VPWR VPWR _16011_/X sky130_fd_sc_hd__and3_4
X_13223_ _12383_/A VGND VGND VPWR VPWR _13260_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21436__B2 _21430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12491__A _13009_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13154_ _12730_/A _23985_/Q VGND VGND VPWR VPWR _13154_/X sky130_fd_sc_hd__or2_4
XFILLER_97_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12105_ _12051_/X _12105_/B _12104_/X VGND VGND VPWR VPWR _12105_/X sky130_fd_sc_hd__or3_4
XFILLER_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13085_ _13080_/A _13085_/B VGND VGND VPWR VPWR _13085_/X sky130_fd_sc_hd__or2_4
X_17962_ _17962_/A VGND VGND VPWR VPWR _17962_/X sky130_fd_sc_hd__buf_2
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19701_ _19674_/X _19699_/Y _20844_/B _19551_/A VGND VGND VPWR VPWR _19701_/X sky130_fd_sc_hd__a2bb2o_4
X_12036_ _16741_/A VGND VGND VPWR VPWR _12036_/X sky130_fd_sc_hd__buf_2
X_16913_ _16909_/B VGND VGND VPWR VPWR _16913_/X sky130_fd_sc_hd__buf_2
XFILLER_61_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21309__A _21301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17893_ _17680_/A VGND VGND VPWR VPWR _17893_/X sky130_fd_sc_hd__buf_2
XANTENNA__20213__A _20212_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19632_ _19629_/B _19631_/Y _19866_/B VGND VGND VPWR VPWR _19633_/D sky130_fd_sc_hd__o21a_4
XANTENNA__15307__A _13927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11835__A _11675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20411__A2 _20410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16844_ _13277_/X _16833_/Y VGND VGND VPWR VPWR _16845_/D sky130_fd_sc_hd__nand2_4
XFILLER_4_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19563_ _24149_/Q _19435_/A HRDATA[23] _19431_/X VGND VGND VPWR VPWR _19563_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11554__B IRQ[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16775_ _16799_/A _16775_/B VGND VGND VPWR VPWR _16775_/X sky130_fd_sc_hd__or2_4
X_13987_ _13987_/A _13987_/B VGND VGND VPWR VPWR _13987_/X sky130_fd_sc_hd__and2_4
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18618__A _18216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18514_ _18348_/A _18348_/B VGND VGND VPWR VPWR _18514_/Y sky130_fd_sc_hd__nand2_4
X_15726_ _12777_/X _15726_/B _15726_/C VGND VGND VPWR VPWR _15727_/C sky130_fd_sc_hd__and3_4
X_12938_ _12974_/A _23283_/Q VGND VGND VPWR VPWR _12939_/C sky130_fd_sc_hd__or2_4
X_19494_ _19454_/A VGND VGND VPWR VPWR _19494_/X sky130_fd_sc_hd__buf_2
XFILLER_34_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21911__A2 _21908_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21044__A _21015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18445_ _18445_/A VGND VGND VPWR VPWR _18445_/Y sky130_fd_sc_hd__inv_2
X_15657_ _12720_/A _15657_/B _15657_/C VGND VGND VPWR VPWR _15657_/X sky130_fd_sc_hd__and3_4
X_12869_ _12477_/X _23987_/Q VGND VGND VPWR VPWR _12869_/X sky130_fd_sc_hd__or2_4
XANTENNA__12666__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14608_ _14143_/A _14689_/B VGND VGND VPWR VPWR _14608_/X sky130_fd_sc_hd__or2_4
X_18376_ _18314_/X _18356_/X _18357_/X _18375_/X VGND VGND VPWR VPWR _18376_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21124__B1 _16398_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15588_ _15616_/A _15588_/B _15588_/C VGND VGND VPWR VPWR _15589_/C sky130_fd_sc_hd__and3_4
XFILLER_33_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17327_ _17325_/X _17326_/X VGND VGND VPWR VPWR _17327_/X sky130_fd_sc_hd__and2_4
XANTENNA__17879__B1 _17878_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20478__A2 _20477_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14539_ _14500_/X _14539_/B VGND VGND VPWR VPWR _14541_/B sky130_fd_sc_hd__or2_4
XFILLER_72_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21675__B2 _21673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19449__A _19449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17258_ _17860_/A _17255_/X _17868_/A VGND VGND VPWR VPWR _17258_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__15696__B _15769_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16209_ _16202_/A _16132_/B VGND VGND VPWR VPWR _16209_/X sky130_fd_sc_hd__or2_4
XANTENNA__13497__A _12926_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21427__B2 _21423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17189_ _17152_/X _17187_/X _17154_/X _17188_/X VGND VGND VPWR VPWR _17189_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16854__A1 _16840_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20123__A _20122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22910_ _18640_/X _22908_/Y _22924_/A _22909_/X VGND VGND VPWR VPWR _22911_/C sky130_fd_sc_hd__a211o_4
XANTENNA__11745__A _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15217__A _11661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23890_ _23826_/CLK _21321_/X VGND VGND VPWR VPWR _13104_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_68_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14121__A _14121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22841_ _14786_/Y _22826_/X _22794_/A VGND VGND VPWR VPWR _22841_/X sky130_fd_sc_hd__o21a_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24320__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13960__A _13960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22772_ _22772_/A VGND VGND VPWR VPWR _22773_/A sky130_fd_sc_hd__inv_2
XFILLER_77_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21902__A2 _21901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21723_ _21702_/A VGND VGND VPWR VPWR _21723_/X sky130_fd_sc_hd__buf_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12576__A _13700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24442_ _24277_/CLK _18773_/X HRESETn VGND VGND VPWR VPWR _24442_/Q sky130_fd_sc_hd__dfrtp_4
X_21654_ _21529_/X _21648_/X _12827_/B _21652_/X VGND VGND VPWR VPWR _23700_/D sky130_fd_sc_hd__o22a_4
X_20605_ _20605_/A VGND VGND VPWR VPWR _20605_/Y sky130_fd_sc_hd__inv_2
X_24373_ _24277_/CLK _18890_/X HRESETn VGND VGND VPWR VPWR _24373_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__15887__A _15892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19359__A _19370_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21585_ _21584_/X VGND VGND VPWR VPWR _21590_/A sky130_fd_sc_hd__buf_2
XFILLER_90_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14791__A _13862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18263__A _18204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23324_ _23324_/CLK _22302_/X VGND VGND VPWR VPWR _16550_/B sky130_fd_sc_hd__dfxtp_4
X_20536_ _22100_/A VGND VGND VPWR VPWR _21246_/A sky130_fd_sc_hd__buf_2
XFILLER_119_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23255_ _23313_/CLK _22407_/X VGND VGND VPWR VPWR _16158_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21418__B2 _21416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20467_ _20467_/A VGND VGND VPWR VPWR _20603_/A sky130_fd_sc_hd__buf_2
XFILLER_106_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22206_ _22200_/Y _22205_/X _22073_/X _22205_/X VGND VGND VPWR VPWR _22206_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23186_ _23122_/CLK _22538_/X VGND VGND VPWR VPWR _13005_/B sky130_fd_sc_hd__dfxtp_4
X_20398_ _20512_/A VGND VGND VPWR VPWR _20398_/X sky130_fd_sc_hd__buf_2
X_22137_ _22125_/A VGND VGND VPWR VPWR _22137_/X sky130_fd_sc_hd__buf_2
XANTENNA__22918__A1 _22886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22068_ _22068_/A _21917_/B _21784_/C _21008_/A VGND VGND VPWR VPWR _22068_/X sky130_fd_sc_hd__or4_4
XFILLER_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20033__A _19985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11655__A _13918_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19795__B1 _19872_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13910_ _13910_/A _24071_/Q VGND VGND VPWR VPWR _13911_/C sky130_fd_sc_hd__or2_4
X_21019_ _20356_/X _21016_/X _24059_/Q _21013_/X VGND VGND VPWR VPWR _21019_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15127__A _12196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14890_ _13985_/A _14890_/B _14889_/X VGND VGND VPWR VPWR _14894_/B sky130_fd_sc_hd__and3_4
XFILLER_74_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13841_ _13887_/A _13841_/B VGND VGND VPWR VPWR _13846_/B sky130_fd_sc_hd__or2_4
XFILLER_1_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_121_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR _23983_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14966__A _15074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22146__A2 _22137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13772_ _11656_/A _13772_/B _13772_/C VGND VGND VPWR VPWR _13772_/X sky130_fd_sc_hd__and3_4
X_16560_ _12020_/A _16558_/X _16560_/C VGND VGND VPWR VPWR _16560_/X sky130_fd_sc_hd__and3_4
XANTENNA__23063__B _23062_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20157__A1 _24434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15511_ _15480_/A _15511_/B VGND VGND VPWR VPWR _15511_/X sky130_fd_sc_hd__or2_4
X_12723_ _15664_/A _12721_/X _12723_/C VGND VGND VPWR VPWR _12723_/X sky130_fd_sc_hd__and3_4
X_16491_ _16499_/A _16489_/X _16490_/X VGND VGND VPWR VPWR _16491_/X sky130_fd_sc_hd__and3_4
XANTENNA__12486__A _13622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18770__A1 _12184_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18230_ _17667_/A _16981_/B _18174_/B VGND VGND VPWR VPWR _22998_/B sky130_fd_sc_hd__a21o_4
X_12654_ _12970_/A _12654_/B _12654_/C VGND VGND VPWR VPWR _12654_/X sky130_fd_sc_hd__and3_4
X_15442_ _15442_/A _15442_/B _15442_/C VGND VGND VPWR VPWR _15442_/X sky130_fd_sc_hd__or3_4
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24456__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21799__A _21799_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21106__B1 _15262_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _11905_/A VGND VGND VPWR VPWR _11606_/A sky130_fd_sc_hd__buf_2
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21657__A1 _21534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18161_ _17476_/C _18158_/X _18160_/X VGND VGND VPWR VPWR _18161_/Y sky130_fd_sc_hd__a21oi_4
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15797__A _15820_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12585_/A VGND VGND VPWR VPWR _12981_/A sky130_fd_sc_hd__buf_2
X_15373_ _14000_/A _15299_/B VGND VGND VPWR VPWR _15373_/X sky130_fd_sc_hd__or2_4
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21657__B2 _21652_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17112_ _17109_/Y _17010_/X _17018_/X _17111_/X VGND VGND VPWR VPWR _17322_/B sky130_fd_sc_hd__o22a_4
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11536_ _20855_/A IRQ[6] VGND VGND VPWR VPWR _11536_/X sky130_fd_sc_hd__and2_4
X_14324_ _14432_/A _14324_/B VGND VGND VPWR VPWR _14325_/C sky130_fd_sc_hd__or2_4
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18092_ _18056_/X _18091_/X _19986_/A _18056_/X VGND VGND VPWR VPWR _24472_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23480__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20208__A _20421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16405__B _16405_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14255_ _14359_/A _23209_/Q VGND VGND VPWR VPWR _14257_/B sky130_fd_sc_hd__or2_4
X_17043_ _17043_/A VGND VGND VPWR VPWR _17043_/X sky130_fd_sc_hd__buf_2
XFILLER_7_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13206_ _12383_/A VGND VGND VPWR VPWR _13228_/A sky130_fd_sc_hd__buf_2
X_14186_ _14186_/A _23337_/Q VGND VGND VPWR VPWR _14189_/B sky130_fd_sc_hd__or2_4
XANTENNA__22082__B2 _22072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11549__B IRQ[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24391__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22423__A _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13137_ _12221_/X _13137_/B VGND VGND VPWR VPWR _13137_/X sky130_fd_sc_hd__or2_4
X_18994_ _18994_/A VGND VGND VPWR VPWR _18994_/X sky130_fd_sc_hd__buf_2
XANTENNA__16421__A _16002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13068_ _13097_/A VGND VGND VPWR VPWR _13128_/A sky130_fd_sc_hd__buf_2
X_17945_ _16935_/X _17898_/X _17006_/X _17944_/X VGND VGND VPWR VPWR _17945_/X sky130_fd_sc_hd__o22a_4
XFILLER_117_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12019_ _11962_/X _23806_/Q VGND VGND VPWR VPWR _12020_/C sky130_fd_sc_hd__or2_4
XFILLER_117_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15037__A _15037_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19732__A _19784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17876_ _17270_/X _17875_/X VGND VGND VPWR VPWR _17876_/Y sky130_fd_sc_hd__nand2_4
XFILLER_94_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20878__A HRDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19615_ _19553_/A HRDATA[10] VGND VGND VPWR VPWR _19615_/X sky130_fd_sc_hd__and2_4
X_16827_ _12680_/B _16826_/X _12677_/X VGND VGND VPWR VPWR _16827_/X sky130_fd_sc_hd__o21a_4
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14876__A _14906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19546_ _20317_/B _19551_/A _19497_/X HRDATA[13] VGND VGND VPWR VPWR _19546_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16758_ _16772_/A _24027_/Q VGND VGND VPWR VPWR _16760_/B sky130_fd_sc_hd__or2_4
XFILLER_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21345__B1 _23872_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20148__B2 IRQ[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15709_ _13004_/A _15705_/X _15708_/X VGND VGND VPWR VPWR _15709_/X sky130_fd_sc_hd__or3_4
X_19477_ _19477_/A VGND VGND VPWR VPWR _19541_/A sky130_fd_sc_hd__buf_2
XANTENNA__21896__B2 _21891_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16689_ _16689_/A _16685_/X _16688_/X VGND VGND VPWR VPWR _16689_/X sky130_fd_sc_hd__or3_4
XFILLER_62_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_26_0_HCLK clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18428_ _18428_/A _18427_/X VGND VGND VPWR VPWR _18428_/X sky130_fd_sc_hd__or2_4
XFILLER_22_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21502__A _21527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18359_ _18295_/A _17480_/X VGND VGND VPWR VPWR _18362_/B sky130_fd_sc_hd__nor2_4
XFILLER_33_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15500__A _12612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21370_ _21246_/X _21369_/X _23859_/Q _21366_/X VGND VGND VPWR VPWR _21370_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12843__B _12841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20321_ _20493_/A VGND VGND VPWR VPWR _20321_/X sky130_fd_sc_hd__buf_2
XANTENNA__18306__A1_N _18189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14116__A _14143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18811__A _12100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13020__A _13020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23040_ _23014_/X _17951_/A _23026_/X _23039_/X VGND VGND VPWR VPWR _23041_/A sky130_fd_sc_hd__a211o_4
XFILLER_31_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20252_ _18867_/X VGND VGND VPWR VPWR _20473_/A sky130_fd_sc_hd__inv_2
XFILLER_115_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17427__A _14263_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20183_ _20183_/A VGND VGND VPWR VPWR _24110_/D sky130_fd_sc_hd__inv_2
XANTENNA__21820__B2 _21812_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23203__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22376__A2 _22375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23942_ _23845_/CLK _21202_/X VGND VGND VPWR VPWR _14302_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_69_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20387__A1 _18050_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23873_ _23487_/CLK _21344_/X VGND VGND VPWR VPWR _23873_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19792__A3 _19791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22128__A2 _22125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13690__A _13690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22824_ _18759_/A _22824_/B VGND VGND VPWR VPWR _22824_/X sky130_fd_sc_hd__or2_4
XFILLER_25_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22755_ _22751_/X _22755_/B _22754_/X VGND VGND VPWR VPWR _24097_/D sky130_fd_sc_hd__and3_4
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21706_ _21531_/X _21705_/X _23667_/Q _21702_/X VGND VGND VPWR VPWR _21706_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22686_ _22686_/A VGND VGND VPWR VPWR _22686_/X sky130_fd_sc_hd__buf_2
XFILLER_52_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24425_ _24425_/CLK _18798_/X HRESETn VGND VGND VPWR VPWR _20762_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21412__A _21419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21637_ _21659_/A VGND VGND VPWR VPWR _21637_/X sky130_fd_sc_hd__buf_2
XANTENNA__21639__B2 _21638_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19701__B1 _20844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15410__A _12211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12370_ _12388_/A _12368_/X _12370_/C VGND VGND VPWR VPWR _12370_/X sky130_fd_sc_hd__and3_4
X_24356_ _24321_/CLK _24356_/D HRESETn VGND VGND VPWR VPWR _19083_/A sky130_fd_sc_hd__dfstp_4
X_21568_ _21556_/A VGND VGND VPWR VPWR _21568_/X sky130_fd_sc_hd__buf_2
XFILLER_103_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23307_ _23557_/CLK _23307_/D VGND VGND VPWR VPWR _15539_/B sky130_fd_sc_hd__dfxtp_4
X_20519_ _20519_/A _20519_/B VGND VGND VPWR VPWR _20519_/Y sky130_fd_sc_hd__nand2_4
X_24287_ _24290_/CLK _24287_/D HRESETn VGND VGND VPWR VPWR _19108_/B sky130_fd_sc_hd__dfrtp_4
X_21499_ _21112_/A _21348_/B _21784_/C _20199_/B VGND VGND VPWR VPWR _21500_/A sky130_fd_sc_hd__or4_4
XANTENNA__24149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_46_0_HCLK clkbuf_7_46_0_HCLK/A VGND VGND VPWR VPWR _23847_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18721__A _18720_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14040_ _11798_/A VGND VGND VPWR VPWR _14040_/X sky130_fd_sc_hd__buf_2
X_23238_ _23494_/CLK _23238_/D VGND VGND VPWR VPWR _14268_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_5_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22064__B2 _22020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22243__A _22207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23169_ _23233_/CLK _23169_/D VGND VGND VPWR VPWR _15132_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_84_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18283__A3 _18273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15991_ _15986_/A _15988_/X _15991_/C VGND VGND VPWR VPWR _15995_/B sky130_fd_sc_hd__and3_4
XFILLER_62_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19768__B1 _16599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22367__A2 _22361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17730_ _17732_/B _17729_/X VGND VGND VPWR VPWR _17730_/X sky130_fd_sc_hd__or2_4
XANTENNA__19552__A _19416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14942_ _15074_/A _14883_/B VGND VGND VPWR VPWR _14942_/X sky130_fd_sc_hd__or2_4
X_17661_ _17661_/A _17459_/Y VGND VGND VPWR VPWR _17755_/A sky130_fd_sc_hd__and2_4
X_14873_ _14867_/X _14873_/B VGND VGND VPWR VPWR _14873_/X sky130_fd_sc_hd__or2_4
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19400_ _19396_/X _18518_/Y _19399_/X _24201_/Q VGND VGND VPWR VPWR _19400_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16612_ _16599_/X _16612_/B _16612_/C VGND VGND VPWR VPWR _16612_/X sky130_fd_sc_hd__or3_4
X_13824_ _15436_/A _13824_/B VGND VGND VPWR VPWR _13826_/B sky130_fd_sc_hd__or2_4
X_17592_ _17349_/A _17356_/X _17360_/Y VGND VGND VPWR VPWR _17592_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19331_ _19328_/X _18311_/X _19328_/X _24241_/Q VGND VGND VPWR VPWR _19331_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16543_ _12020_/A VGND VGND VPWR VPWR _16569_/A sky130_fd_sc_hd__buf_2
X_13755_ _12612_/A _13755_/B _13755_/C VGND VGND VPWR VPWR _13771_/B sky130_fd_sc_hd__and3_4
XFILLER_62_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21878__B2 _21877_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ _12706_/A _12706_/B _12705_/X VGND VGND VPWR VPWR _12706_/X sky130_fd_sc_hd__or3_4
X_19262_ _24273_/Q _19263_/A _19261_/Y VGND VGND VPWR VPWR _24273_/D sky130_fd_sc_hd__o21a_4
X_16474_ _16473_/X _16398_/B VGND VGND VPWR VPWR _16475_/C sky130_fd_sc_hd__or2_4
X_13686_ _13686_/A VGND VGND VPWR VPWR _13884_/A sky130_fd_sc_hd__buf_2
XANTENNA__22418__A _20552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18213_ _17862_/X _18037_/X _17869_/X VGND VGND VPWR VPWR _18213_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_73_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15425_ _15429_/A _23596_/Q VGND VGND VPWR VPWR _15425_/X sky130_fd_sc_hd__or2_4
X_12637_ _12957_/A _12610_/X _12636_/X VGND VGND VPWR VPWR _12673_/B sky130_fd_sc_hd__or3_4
X_19193_ _19112_/X VGND VGND VPWR VPWR _19193_/Y sky130_fd_sc_hd__inv_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12944__A _12982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18144_ _17921_/X _17981_/Y _17926_/X _17978_/Y VGND VGND VPWR VPWR _18144_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23996__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12568_ _12568_/A VGND VGND VPWR VPWR _13718_/A sky130_fd_sc_hd__buf_2
X_15356_ _15314_/A _15290_/B VGND VGND VPWR VPWR _15357_/C sky130_fd_sc_hd__or2_4
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16135__B _16135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11519_ _11519_/A _11519_/B VGND VGND VPWR VPWR _11520_/B sky130_fd_sc_hd__or2_4
X_14307_ _15558_/A _14303_/X _14306_/X VGND VGND VPWR VPWR _14307_/X sky130_fd_sc_hd__or3_4
XFILLER_116_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18075_ _18075_/A VGND VGND VPWR VPWR _18075_/Y sky130_fd_sc_hd__inv_2
X_12499_ _12211_/X VGND VGND VPWR VPWR _13016_/A sky130_fd_sc_hd__buf_2
X_15287_ _12860_/A _15285_/X _15286_/X VGND VGND VPWR VPWR _15287_/X sky130_fd_sc_hd__and3_4
XFILLER_7_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17026_ _17467_/B VGND VGND VPWR VPWR _17457_/B sky130_fd_sc_hd__buf_2
X_14238_ _13839_/A VGND VGND VPWR VPWR _14251_/A sky130_fd_sc_hd__buf_2
XANTENNA__22055__B2 _22049_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22153__A _22153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14169_ _15023_/A _23849_/Q VGND VGND VPWR VPWR _14169_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_3_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_113_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21992__A _21985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18977_ _18971_/X _18976_/X _18971_/X _11528_/A VGND VGND VPWR VPWR _18977_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17928_ _17928_/A VGND VGND VPWR VPWR _17928_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17859_ _17858_/X VGND VGND VPWR VPWR _17871_/A sky130_fd_sc_hd__buf_2
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20870_ _20870_/A VGND VGND VPWR VPWR _20870_/X sky130_fd_sc_hd__buf_2
XANTENNA__21318__B1 _23892_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19529_ _19494_/X _19498_/Y _19499_/Y _19528_/X VGND VGND VPWR VPWR _19529_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22530__A2 _22529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22540_ _22533_/A VGND VGND VPWR VPWR _22540_/X sky130_fd_sc_hd__buf_2
XANTENNA__13015__A _13015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20541__B2 _20449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21232__A _21802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22471_ _22471_/A VGND VGND VPWR VPWR _22486_/A sky130_fd_sc_hd__buf_2
XFILLER_10_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12854__A _12464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16326__A _16364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24210_ _23812_/CLK _19387_/X HRESETn VGND VGND VPWR VPWR _24210_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24001__CLK _24065_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21422_ _21251_/X _21419_/X _13179_/B _21416_/X VGND VGND VPWR VPWR _23825_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15230__A _15203_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21097__A2 _21096_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22294__B2 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24141_ _24229_/CLK _24141_/D HRESETn VGND VGND VPWR VPWR _24141_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21353_ _21347_/Y _21352_/X _21219_/X _21352_/X VGND VGND VPWR VPWR _21353_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20304_ _20293_/X _20302_/X _11533_/D _20303_/X VGND VGND VPWR VPWR _20304_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24072_ _23368_/CLK _24072_/D VGND VGND VPWR VPWR _24072_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22046__B2 _22042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21284_ _21282_/X _21283_/X _23908_/Q _21278_/X VGND VGND VPWR VPWR _21284_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15884__B _23821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24151__CLK _24223_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23023_ _23018_/A _23023_/B _23023_/C VGND VGND VPWR VPWR _23023_/X sky130_fd_sc_hd__and3_4
XFILLER_2_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13685__A _13684_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20235_ _20235_/A VGND VGND VPWR VPWR _20467_/A sky130_fd_sc_hd__buf_2
XFILLER_103_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20166_ _20166_/A _20165_/Y VGND VGND VPWR VPWR _20166_/X sky130_fd_sc_hd__or2_4
XANTENNA__18670__B1 _18398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16996__A _16996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22349__A2 _22347_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20097_ _20090_/B VGND VGND VPWR VPWR _20097_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23925_ _23315_/CLK _23925_/D VGND VGND VPWR VPWR _12614_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_58_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11933__A _12914_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15405__A _13813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11870_ _12465_/A VGND VGND VPWR VPWR _13014_/A sky130_fd_sc_hd__buf_2
XFILLER_72_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23856_ _24047_/CLK _23856_/D VGND VGND VPWR VPWR _13344_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20780__A1 _20750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20780__B2 _20724_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22807_ _22807_/A _17109_/Y VGND VGND VPWR VPWR _22807_/X sky130_fd_sc_hd__or2_4
XANTENNA__11652__B _12421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20999_ _20282_/A _20998_/X VGND VGND VPWR VPWR _20999_/Y sky130_fd_sc_hd__nand2_4
X_23787_ _24044_/CLK _21482_/X VGND VGND VPWR VPWR _23787_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18716__A _18728_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13540_ _15884_/A _13540_/B VGND VGND VPWR VPWR _13540_/X sky130_fd_sc_hd__or2_4
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22738_ SYSTICKCLKDIV[4] VGND VGND VPWR VPWR _22738_/Y sky130_fd_sc_hd__inv_2
X_13471_ _13467_/A _13469_/X _13471_/C VGND VGND VPWR VPWR _13471_/X sky130_fd_sc_hd__and3_4
X_22669_ _22668_/X VGND VGND VPWR VPWR _22669_/X sky130_fd_sc_hd__buf_2
XANTENNA__16236__A _16155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12764__A _12412_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12422_ _12967_/A VGND VGND VPWR VPWR _13550_/A sky130_fd_sc_hd__buf_2
X_15210_ _15234_/A _15210_/B VGND VGND VPWR VPWR _15210_/X sky130_fd_sc_hd__or2_4
X_24408_ _24277_/CLK _24408_/D HRESETn VGND VGND VPWR VPWR _24408_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21088__A2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16190_ _16206_/A _16186_/X _16189_/X VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__and3_4
XFILLER_12_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13579__B _13425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22285__B2 _22283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20981__A _22460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12353_ _12388_/A _12351_/X _12352_/X VGND VGND VPWR VPWR _12353_/X sky130_fd_sc_hd__and3_4
X_15141_ _14108_/A _15139_/X _15140_/X VGND VGND VPWR VPWR _15141_/X sky130_fd_sc_hd__and3_4
X_24339_ _23358_/CLK _19001_/X HRESETn VGND VGND VPWR VPWR _11524_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__17700__A2 _17375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15072_ _15072_/A VGND VGND VPWR VPWR _15109_/A sky130_fd_sc_hd__buf_2
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12284_ _12496_/A VGND VGND VPWR VPWR _12284_/X sky130_fd_sc_hd__buf_2
XANTENNA__15711__A1 _12716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22037__B2 _22035_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15794__B _15855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23069__A _16893_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14023_ _14815_/A _14023_/B _14023_/C VGND VGND VPWR VPWR _14029_/B sky130_fd_sc_hd__and3_4
X_18900_ _13575_/X _18898_/X _24367_/Q _18899_/X VGND VGND VPWR VPWR _24367_/D sky130_fd_sc_hd__o22a_4
XFILLER_107_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22588__A2 _22586_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13595__A _13595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19880_ _19740_/A _19880_/B VGND VGND VPWR VPWR _19880_/X sky130_fd_sc_hd__or2_4
XFILLER_84_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18256__A3 _18252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19453__A2 _19545_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21796__B1 _23612_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18831_ _16233_/X _18827_/X _20426_/A _18828_/X VGND VGND VPWR VPWR _24407_/D sky130_fd_sc_hd__o22a_4
XFILLER_84_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18661__B1 _18107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21260__A2 _21259_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18762_ _18762_/A _18761_/X VGND VGND VPWR VPWR _18762_/X sky130_fd_sc_hd__or2_4
X_15974_ _15939_/A _23896_/Q VGND VGND VPWR VPWR _15974_/X sky130_fd_sc_hd__or2_4
X_17713_ _16969_/A _17385_/X VGND VGND VPWR VPWR _17713_/X sky130_fd_sc_hd__or2_4
X_14925_ _14925_/A _14923_/X _14925_/C VGND VGND VPWR VPWR _14926_/C sky130_fd_sc_hd__and3_4
XFILLER_76_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18693_ _17327_/X _18693_/B VGND VGND VPWR VPWR _18693_/Y sky130_fd_sc_hd__nand2_4
XFILLER_63_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12939__A _12951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11843__A _11842_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17644_ _17644_/A _17535_/A VGND VGND VPWR VPWR _17765_/A sky130_fd_sc_hd__and2_4
XANTENNA__15315__A _14207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14856_ _13953_/A _14856_/B VGND VGND VPWR VPWR _14856_/X sky130_fd_sc_hd__or2_4
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12658__B _12658_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13807_ _13614_/A _13807_/B VGND VGND VPWR VPWR _13807_/X sky130_fd_sc_hd__or2_4
XANTENNA__11562__B IRQ[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17575_ _18047_/A _17573_/X _17574_/Y VGND VGND VPWR VPWR _17575_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15034__B _24063_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14787_ _13872_/A _14787_/B VGND VGND VPWR VPWR _14787_/X sky130_fd_sc_hd__or2_4
X_11999_ _11999_/A _11995_/X _11999_/C VGND VGND VPWR VPWR _11999_/X sky130_fd_sc_hd__or3_4
XFILLER_1_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19314_ _19303_/X _17771_/X _19313_/X _24253_/Q VGND VGND VPWR VPWR _24253_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22512__A2 _22507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20875__B _20317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16526_ _12022_/A VGND VGND VPWR VPWR _16538_/A sky130_fd_sc_hd__buf_2
X_13738_ _13738_/A _13738_/B _13738_/C VGND VGND VPWR VPWR _13739_/C sky130_fd_sc_hd__or3_4
XANTENNA__15969__B _15969_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14873__B _14873_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19245_ _19245_/A VGND VGND VPWR VPWR _19245_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16457_ _11727_/X _16457_/B _16456_/X VGND VGND VPWR VPWR _16457_/X sky130_fd_sc_hd__and3_4
XFILLER_31_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13669_ _13636_/A _24072_/Q VGND VGND VPWR VPWR _13669_/X sky130_fd_sc_hd__or2_4
XFILLER_108_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12674__A _12673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15408_ _15431_/A _15406_/X _15407_/X VGND VGND VPWR VPWR _15408_/X sky130_fd_sc_hd__and3_4
X_19176_ _19121_/A _19177_/A _19175_/Y VGND VGND VPWR VPWR _24300_/D sky130_fd_sc_hd__o21a_4
XFILLER_34_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16388_ _15997_/A _16388_/B VGND VGND VPWR VPWR _16389_/C sky130_fd_sc_hd__or2_4
XANTENNA__24174__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11567__A2 IRQ[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18127_ _18009_/X _18125_/X _18053_/X _18126_/X VGND VGND VPWR VPWR _18127_/X sky130_fd_sc_hd__o22a_4
X_15339_ _15332_/A _15266_/B VGND VGND VPWR VPWR _15339_/X sky130_fd_sc_hd__or2_4
XFILLER_8_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18361__A _18297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18058_ _18012_/X _18013_/B VGND VGND VPWR VPWR _18058_/Y sky130_fd_sc_hd__nand2_4
X_17009_ _17009_/A _17072_/A VGND VGND VPWR VPWR _17010_/A sky130_fd_sc_hd__or2_4
XFILLER_113_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_92_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR _23774_/CLK sky130_fd_sc_hd__clkbuf_1
X_20020_ _19996_/A VGND VGND VPWR VPWR _20020_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18404__B1 _18398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21971_ _21970_/X VGND VGND VPWR VPWR _21971_/X sky130_fd_sc_hd__buf_2
XANTENNA__12849__A _12849_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20922_ HRDATA[3] VGND VGND VPWR VPWR _20922_/Y sky130_fd_sc_hd__inv_2
X_23710_ _23774_/CLK _23710_/D VGND VGND VPWR VPWR _23710_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20853_ _20841_/X _20848_/X _20852_/X VGND VGND VPWR VPWR _20853_/X sky130_fd_sc_hd__a21o_4
X_23641_ _23770_/CLK _23641_/D VGND VGND VPWR VPWR _16368_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22503__A2 _22500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19904__B1 _20224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17440__A _12101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23572_ _23539_/CLK _21886_/X VGND VGND VPWR VPWR _23572_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20784_ _20619_/X _20783_/X _20617_/X VGND VGND VPWR VPWR _20784_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22523_ _22390_/X _22522_/X _12128_/B _22519_/X VGND VGND VPWR VPWR _22523_/X sky130_fd_sc_hd__o22a_4
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12584__A _12605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22454_ _20915_/A VGND VGND VPWR VPWR _22454_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21405_ _21419_/A VGND VGND VPWR VPWR _21405_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15895__A _13554_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19367__A _19370_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22385_ _22384_/X VGND VGND VPWR VPWR _22423_/A sky130_fd_sc_hd__inv_2
XFILLER_108_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24124_ _24126_/CLK _20037_/Y HRESETn VGND VGND VPWR VPWR _16952_/A sky130_fd_sc_hd__dfrtp_4
X_21336_ _21275_/X _21333_/X _13807_/B _21330_/X VGND VGND VPWR VPWR _21336_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21490__A2 _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24055_ _23316_/CLK _24055_/D VGND VGND VPWR VPWR _24055_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11928__A _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21267_ _21265_/X _21259_/X _23915_/Q _21266_/X VGND VGND VPWR VPWR _21267_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14304__A _14283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21778__B1 _14773_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23006_ _22985_/X _16946_/Y _22997_/X _23005_/X VGND VGND VPWR VPWR _23006_/X sky130_fd_sc_hd__a211o_4
X_20218_ _20218_/A HRDATA[15] VGND VGND VPWR VPWR _20218_/X sky130_fd_sc_hd__or2_4
X_21198_ _20779_/X _21197_/X _23945_/Q _21194_/X VGND VGND VPWR VPWR _23945_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22521__A _22521_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22990__A2 _17674_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20149_ _24420_/Q IRQ[5] _20147_/Y _20148_/X VGND VGND VPWR VPWR _20149_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__14958__B _23584_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21137__A _21130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12971_ _12655_/A _12967_/X _12971_/C VGND VGND VPWR VPWR _12971_/X sky130_fd_sc_hd__or3_4
XFILLER_58_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12759__A _12605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14710_ _11697_/A _14624_/B VGND VGND VPWR VPWR _14712_/B sky130_fd_sc_hd__or2_4
XFILLER_111_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24047__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15135__A _11879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11663__A _13886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11922_ _11921_/X _23742_/Q VGND VGND VPWR VPWR _11923_/C sky130_fd_sc_hd__or2_4
X_23908_ _23107_/CLK _21284_/X VGND VGND VPWR VPWR _23908_/Q sky130_fd_sc_hd__dfxtp_4
X_15690_ _12722_/A _15690_/B VGND VGND VPWR VPWR _15691_/C sky130_fd_sc_hd__or2_4
XANTENNA__21950__B1 _23531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12478__B _12607_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14641_ _11638_/A VGND VGND VPWR VPWR _14642_/A sky130_fd_sc_hd__buf_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11853_ _11852_/X VGND VGND VPWR VPWR _11853_/X sky130_fd_sc_hd__buf_2
X_23839_ _23217_/CLK _21396_/X VGND VGND VPWR VPWR _23839_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__18446__A _18327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17360_ _17360_/A VGND VGND VPWR VPWR _17360_/Y sky130_fd_sc_hd__inv_2
X_11784_ _11685_/X VGND VGND VPWR VPWR _11824_/A sky130_fd_sc_hd__buf_2
X_14572_ _14994_/A VGND VGND VPWR VPWR _15144_/A sky130_fd_sc_hd__buf_2
XFILLER_60_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16311_ _16323_/A _16245_/B VGND VGND VPWR VPWR _16311_/X sky130_fd_sc_hd__or2_4
X_13523_ _12980_/A VGND VGND VPWR VPWR _13561_/A sky130_fd_sc_hd__buf_2
XFILLER_57_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17291_ _14493_/Y _17012_/A _17018_/X _17290_/X VGND VGND VPWR VPWR _17294_/B sky130_fd_sc_hd__o22a_4
XFILLER_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12494__A _12494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19030_ _19002_/A VGND VGND VPWR VPWR _19030_/X sky130_fd_sc_hd__buf_2
X_16242_ _16147_/A _16240_/X _16241_/X VGND VGND VPWR VPWR _16242_/X sky130_fd_sc_hd__and3_4
X_13454_ _12865_/A _13521_/B VGND VGND VPWR VPWR _13454_/X sky130_fd_sc_hd__or2_4
XFILLER_16_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20269__B1 _20493_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12405_ _12388_/A _12405_/B _12404_/X VGND VGND VPWR VPWR _12405_/X sky130_fd_sc_hd__and3_4
X_13385_ _12830_/A VGND VGND VPWR VPWR _13388_/A sky130_fd_sc_hd__buf_2
X_16173_ _13399_/A VGND VGND VPWR VPWR _16206_/A sky130_fd_sc_hd__buf_2
XANTENNA__17134__B1 _17132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15124_ _14918_/X _14988_/X _15123_/Y VGND VGND VPWR VPWR _15124_/X sky130_fd_sc_hd__o21a_4
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12336_ _12892_/A _12292_/X _12300_/X _12326_/X _12335_/X VGND VGND VPWR VPWR _12336_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_6_16_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_12267_ _14128_/A VGND VGND VPWR VPWR _12267_/X sky130_fd_sc_hd__buf_2
X_15055_ _15072_/A VGND VGND VPWR VPWR _15069_/A sky130_fd_sc_hd__buf_2
X_19932_ _11625_/A _19931_/X _23064_/B _11625_/X VGND VGND VPWR VPWR _24141_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19426__A2 _16996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14006_ _14037_/A _13997_/X _14005_/X VGND VGND VPWR VPWR _14019_/B sky130_fd_sc_hd__or3_4
X_19863_ _19846_/B _19881_/A _19740_/A _19862_/Y VGND VGND VPWR VPWR _19863_/X sky130_fd_sc_hd__o22a_4
X_12198_ _13631_/A VGND VGND VPWR VPWR _12198_/X sky130_fd_sc_hd__buf_2
XFILLER_64_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18814_ _18813_/X VGND VGND VPWR VPWR _18814_/X sky130_fd_sc_hd__buf_2
XANTENNA__17525__A _17182_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19794_ _19730_/A _19522_/X VGND VGND VPWR VPWR _19794_/X sky130_fd_sc_hd__and2_4
XFILLER_23_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20992__A1 _20403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20992__B2 _20497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14868__B _14868_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18745_ _18744_/X VGND VGND VPWR VPWR _18745_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15957_ _15957_/A _23992_/Q VGND VGND VPWR VPWR _15958_/C sky130_fd_sc_hd__or2_4
XANTENNA__12669__A _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14908_ _13956_/A _14904_/X _14907_/X VGND VGND VPWR VPWR _14908_/X sky130_fd_sc_hd__or3_4
X_18676_ _18066_/A _17609_/Y VGND VGND VPWR VPWR _18676_/X sky130_fd_sc_hd__and2_4
XFILLER_37_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19357__A2_N _19356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15888_ _13522_/A _15888_/B _15887_/X VGND VGND VPWR VPWR _15889_/C sky130_fd_sc_hd__and3_4
X_17627_ _17627_/A _18024_/B _17583_/X _18081_/B VGND VGND VPWR VPWR _17628_/C sky130_fd_sc_hd__or4_4
XANTENNA__23414__CLK _23155_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14839_ _14815_/A _14839_/B _14839_/C VGND VGND VPWR VPWR _14839_/X sky130_fd_sc_hd__and3_4
XANTENNA__12029__A3 _11991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17558_ _18066_/B _17558_/B VGND VGND VPWR VPWR _17559_/A sky130_fd_sc_hd__or2_4
XFILLER_75_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_26_0_HCLK_A clkbuf_5_26_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15699__B _15699_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19362__A1 _19306_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16509_ _16194_/A _16507_/X _16509_/C VGND VGND VPWR VPWR _16510_/C sky130_fd_sc_hd__and3_4
X_17489_ _17195_/Y _17488_/X VGND VGND VPWR VPWR _17489_/X sky130_fd_sc_hd__or2_4
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23564__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19228_ _24279_/Q _19251_/A VGND VGND VPWR VPWR _19249_/A sky130_fd_sc_hd__and2_4
XFILLER_20_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22249__B2 _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21510__A _21795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19159_ _19129_/X VGND VGND VPWR VPWR _19159_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16604__A _16800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22170_ _22095_/X _22165_/X _12653_/B _22169_/X VGND VGND VPWR VPWR _22170_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21472__A2 _21470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16323__B _23577_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21121_ _20339_/X _21119_/X _23996_/Q _21116_/X VGND VGND VPWR VPWR _21121_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14124__A _14992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21052_ _20893_/X _21051_/X _14692_/B _21048_/X VGND VGND VPWR VPWR _24036_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22421__B2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20003_ _19994_/X _16945_/Y _20000_/X _20002_/X VGND VGND VPWR VPWR _20003_/X sky130_fd_sc_hd__o22a_4
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20983__A1 _20872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20983__B2 _20202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21454__A2_N _21453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12579__A _12935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21954_ _21843_/X _21952_/X _13636_/B _21949_/X VGND VGND VPWR VPWR _21954_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20735__A1 _20681_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20796__A _22127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20735__B2 _20625_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20905_ _20704_/X _20904_/Y _24259_/Q _20325_/X VGND VGND VPWR VPWR _20905_/X sky130_fd_sc_hd__o22a_4
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _21811_/X _21880_/X _12505_/B _21884_/X VGND VGND VPWR VPWR _21885_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18266__A _18266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14794__A _13872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _24198_/Q _20751_/X _20835_/Y VGND VGND VPWR VPWR _22446_/A sky130_fd_sc_hd__o21a_4
X_23624_ _23304_/CLK _23624_/D VGND VGND VPWR VPWR _13767_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22488__B2 _22483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20767_ _20525_/A VGND VGND VPWR VPWR _20767_/X sky130_fd_sc_hd__buf_2
X_23555_ _23907_/CLK _23555_/D VGND VGND VPWR VPWR _14803_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15402__B _15465_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21160__B2 _21115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22506_ _22449_/X _22500_/X _14479_/B _22504_/X VGND VGND VPWR VPWR _22506_/X sky130_fd_sc_hd__o22a_4
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23486_ _23514_/CLK _22022_/X VGND VGND VPWR VPWR _23486_/Q sky130_fd_sc_hd__dfxtp_4
X_20698_ _20613_/X _20697_/X _15437_/B _20592_/X VGND VGND VPWR VPWR _20698_/X sky130_fd_sc_hd__o22a_4
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22437_ _20747_/A VGND VGND VPWR VPWR _22437_/X sky130_fd_sc_hd__buf_2
XANTENNA__16514__A _16513_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13170_ _12682_/X _13143_/X _13151_/X _13161_/X _13169_/X VGND VGND VPWR VPWR _13170_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_13_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22368_ _22368_/A VGND VGND VPWR VPWR _22368_/X sky130_fd_sc_hd__buf_2
XFILLER_87_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13857__B _23751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22660__B2 _22654_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12121_ _11692_/X _12118_/X _12120_/X VGND VGND VPWR VPWR _12121_/X sky130_fd_sc_hd__and3_4
X_21319_ _21319_/A VGND VGND VPWR VPWR _21319_/X sky130_fd_sc_hd__buf_2
X_24107_ _24230_/CLK _22722_/X HRESETn VGND VGND VPWR VPWR _20190_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11658__A _11657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22299_ _22147_/X _22272_/A _15056_/B _22262_/A VGND VGND VPWR VPWR _23327_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14034__A _11647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12052_ _12083_/A _12128_/B VGND VGND VPWR VPWR _12054_/B sky130_fd_sc_hd__or2_4
X_24038_ _23845_/CLK _24038_/D VGND VGND VPWR VPWR _14305_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22412__A1 _22410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22412__B2 _22411_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14969__A _14243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13873__A _13909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16860_ _15386_/X _14855_/Y _15387_/B VGND VGND VPWR VPWR _16860_/X sky130_fd_sc_hd__o21a_4
XFILLER_46_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15811_ _12891_/A _15807_/X _15811_/C VGND VGND VPWR VPWR _15812_/B sky130_fd_sc_hd__or3_4
XFILLER_19_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23437__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16791_ _16803_/A _16791_/B VGND VGND VPWR VPWR _16791_/X sky130_fd_sc_hd__or2_4
XANTENNA__12489__A _12872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18919__A1 _15121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18530_ _17748_/X _17710_/X _17748_/X _17710_/X VGND VGND VPWR VPWR _18530_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18919__B2 _18892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15742_ _12795_/A _15670_/B VGND VGND VPWR VPWR _15743_/C sky130_fd_sc_hd__or2_4
X_12954_ _12954_/A _12952_/X _12953_/X VGND VGND VPWR VPWR _12954_/X sky130_fd_sc_hd__and3_4
XFILLER_111_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11905_ _11905_/A VGND VGND VPWR VPWR _11905_/Y sky130_fd_sc_hd__inv_2
X_18461_ _24121_/Q _18460_/Y _16974_/B VGND VGND VPWR VPWR _22949_/B sky130_fd_sc_hd__o21a_4
X_15673_ _12235_/A _15729_/B VGND VGND VPWR VPWR _15675_/B sky130_fd_sc_hd__or2_4
XFILLER_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12885_ _12885_/A VGND VGND VPWR VPWR _12886_/A sky130_fd_sc_hd__buf_2
Xclkbuf_5_7_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17412_ _17412_/A VGND VGND VPWR VPWR _17413_/A sky130_fd_sc_hd__inv_2
X_14624_ _14758_/A _14624_/B VGND VGND VPWR VPWR _14626_/B sky130_fd_sc_hd__or2_4
X_11836_ _16677_/A _11836_/B _11836_/C VGND VGND VPWR VPWR _11837_/C sky130_fd_sc_hd__or3_4
X_18392_ _18392_/A _18392_/B VGND VGND VPWR VPWR _18392_/Y sky130_fd_sc_hd__nor2_4
XFILLER_92_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16408__B _16408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19344__B2 _24233_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17343_ _17343_/A _17036_/A VGND VGND VPWR VPWR _17344_/B sky130_fd_sc_hd__and2_4
X_14555_ _14519_/X _14477_/B VGND VGND VPWR VPWR _14555_/X sky130_fd_sc_hd__or2_4
XFILLER_53_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11767_ _13901_/A VGND VGND VPWR VPWR _15484_/A sky130_fd_sc_hd__buf_2
XFILLER_92_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _13494_/X _13499_/X _13505_/X VGND VGND VPWR VPWR _13506_/X sky130_fd_sc_hd__or3_4
XFILLER_119_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17274_ _17039_/X _17273_/X _17043_/X VGND VGND VPWR VPWR _17274_/Y sky130_fd_sc_hd__o21ai_4
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14486_ _13622_/A _14486_/B VGND VGND VPWR VPWR _14488_/B sky130_fd_sc_hd__or2_4
X_11698_ _12383_/A VGND VGND VPWR VPWR _13256_/A sky130_fd_sc_hd__buf_2
X_19013_ _24336_/Q _11521_/B _19008_/Y VGND VGND VPWR VPWR _19013_/Y sky130_fd_sc_hd__a21oi_4
X_16225_ _16162_/X _16225_/B _16225_/C VGND VGND VPWR VPWR _16229_/B sky130_fd_sc_hd__and3_4
XFILLER_35_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21330__A _21316_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13437_ _12518_/X VGND VGND VPWR VPWR _13437_/X sky130_fd_sc_hd__buf_2
X_16156_ _13399_/A VGND VGND VPWR VPWR _16194_/A sky130_fd_sc_hd__buf_2
X_13368_ _13383_/A _13296_/B VGND VGND VPWR VPWR _13369_/C sky130_fd_sc_hd__or2_4
XANTENNA__22651__B2 _22647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15107_ _15107_/A _15105_/X _15107_/C VGND VGND VPWR VPWR _15108_/C sky130_fd_sc_hd__and3_4
X_12319_ _14322_/A VGND VGND VPWR VPWR _12320_/A sky130_fd_sc_hd__buf_2
XANTENNA__19735__A HRDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16087_ _13447_/X VGND VGND VPWR VPWR _16087_/X sky130_fd_sc_hd__buf_2
X_13299_ _15696_/A VGND VGND VPWR VPWR _13300_/A sky130_fd_sc_hd__buf_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15038_ _14778_/A _15038_/B _15038_/C VGND VGND VPWR VPWR _15039_/C sky130_fd_sc_hd__and3_4
X_19915_ _19909_/X _24148_/Q _19910_/X _20844_/B VGND VGND VPWR VPWR _24148_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21206__A2 _21204_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13783__A _15398_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19846_ _19872_/C _19846_/B VGND VGND VPWR VPWR _19846_/X sky130_fd_sc_hd__and2_4
XFILLER_68_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16989_ _16989_/A _16988_/X VGND VGND VPWR VPWR _17000_/A sky130_fd_sc_hd__or2_4
X_19777_ _19719_/A _19718_/A VGND VGND VPWR VPWR _19813_/A sky130_fd_sc_hd__or2_4
XFILLER_83_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12399__A _15882_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22167__B1 _16135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22706__A2 _22700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18728_ _18728_/A _18728_/B VGND VGND VPWR VPWR _18728_/X sky130_fd_sc_hd__or2_4
XFILLER_77_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21914__B1 _23551_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18659_ _18713_/A _17985_/X VGND VGND VPWR VPWR _18659_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15503__A _15491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21670_ _21555_/X _21669_/X _23689_/Q _21666_/X VGND VGND VPWR VPWR _23689_/D sky130_fd_sc_hd__o22a_4
XFILLER_75_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16318__B _16253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20621_ _20617_/X _20620_/X VGND VGND VPWR VPWR _20621_/Y sky130_fd_sc_hd__nand2_4
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21142__B2 _21137_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23340_ _24044_/CLK _22282_/X VGND VGND VPWR VPWR _15458_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_36_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13023__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20552_ _20552_/A VGND VGND VPWR VPWR _21249_/A sky130_fd_sc_hd__buf_2
XANTENNA__21693__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22336__A _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18533__B _18174_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23271_ _23591_/CLK _22371_/X VGND VGND VPWR VPWR _13863_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20483_ _24245_/Q _20421_/X _20482_/X VGND VGND VPWR VPWR _20483_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16334__A _16364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12862__A _12862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22222_ _22222_/A VGND VGND VPWR VPWR _22222_/X sky130_fd_sc_hd__buf_2
XANTENNA__21445__A2 _21440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24343__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22642__B2 _22640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16053__B _15981_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22153_ _22153_/A VGND VGND VPWR VPWR _22169_/A sky130_fd_sc_hd__inv_2
XANTENNA__15124__A2 _14988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21104_ _20893_/X _21103_/X _24004_/Q _21100_/X VGND VGND VPWR VPWR _24004_/D sky130_fd_sc_hd__o22a_4
XFILLER_82_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22084_ _22071_/X VGND VGND VPWR VPWR _22084_/X sky130_fd_sc_hd__buf_2
XANTENNA__15892__B _15836_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22071__A _22108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14789__A _13690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_62_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21035_ _20591_/X _21030_/X _24048_/Q _21034_/X VGND VGND VPWR VPWR _24048_/D sky130_fd_sc_hd__o22a_4
XFILLER_47_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17165__A _17164_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13693__A _14010_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20956__A1 _24193_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14301__B _14301_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19380__A _19379_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12102__A _12101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22986_ _23015_/A VGND VGND VPWR VPWR _22989_/A sky130_fd_sc_hd__buf_2
XANTENNA__19574__A1 _19481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21937_ _21814_/X _21931_/X _12803_/B _21935_/X VGND VGND VPWR VPWR _21937_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16509__A _16194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21381__B2 _21380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11941__A _16143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15413__A _15413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12670_ _12948_/A _12670_/B _12669_/X VGND VGND VPWR VPWR _12671_/C sky130_fd_sc_hd__or3_4
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21868_ _21901_/A VGND VGND VPWR VPWR _21884_/A sky130_fd_sc_hd__inv_2
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19326__B2 _24245_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11602_/X _11620_/X VGND VGND VPWR VPWR _11621_/X sky130_fd_sc_hd__or2_4
X_23607_ _23635_/CLK _21808_/X VGND VGND VPWR VPWR _23607_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20819_ _20819_/A VGND VGND VPWR VPWR _20819_/X sky130_fd_sc_hd__buf_2
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21799_ _21799_/A VGND VGND VPWR VPWR _21799_/X sky130_fd_sc_hd__buf_2
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14029__A _14847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ _14359_/A VGND VGND VPWR VPWR _14341_/A sky130_fd_sc_hd__buf_2
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ _24430_/Q IRQ[15] _11551_/X VGND VGND VPWR VPWR _11552_/X sky130_fd_sc_hd__a21o_4
X_23538_ _23986_/CLK _21940_/X VGND VGND VPWR VPWR _23538_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13868__A _13895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14271_ _12257_/A _14271_/B VGND VGND VPWR VPWR _14271_/X sky130_fd_sc_hd__or2_4
X_23469_ _23826_/CLK _23469_/D VGND VGND VPWR VPWR _15828_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12772__A _12954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16010_ _16025_/A _23512_/Q VGND VGND VPWR VPWR _16011_/C sky130_fd_sc_hd__or2_4
XFILLER_13_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13222_ _13214_/A _13222_/B _13222_/C VGND VGND VPWR VPWR _13227_/B sky130_fd_sc_hd__and3_4
XANTENNA__21436__A2 _21433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13153_ _12728_/A _13153_/B VGND VGND VPWR VPWR _13153_/X sky130_fd_sc_hd__or2_4
XFILLER_3_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12104_ _12100_/X _12102_/X _12104_/C VGND VGND VPWR VPWR _12104_/X sky130_fd_sc_hd__and3_4
X_13084_ _13119_/A _23922_/Q VGND VGND VPWR VPWR _13084_/X sky130_fd_sc_hd__or2_4
X_17961_ _17871_/A VGND VGND VPWR VPWR _17961_/X sky130_fd_sc_hd__buf_2
XFILLER_3_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12035_ _12035_/A VGND VGND VPWR VPWR _16897_/A sky130_fd_sc_hd__buf_2
X_16912_ _16904_/Y _17088_/A _16907_/C _16911_/X VGND VGND VPWR VPWR _16915_/B sky130_fd_sc_hd__a211o_4
X_19700_ HRDATA[22] VGND VGND VPWR VPWR _20844_/B sky130_fd_sc_hd__buf_2
XFILLER_26_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17075__A _18498_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17892_ _17645_/A VGND VGND VPWR VPWR _17951_/A sky130_fd_sc_hd__buf_2
XANTENNA__20947__A1 _20255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16843_ _14077_/X _16842_/X _14077_/X _16842_/X VGND VGND VPWR VPWR _16843_/X sky130_fd_sc_hd__a2bb2o_4
X_19631_ _19867_/B VGND VGND VPWR VPWR _19631_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19562_ _19784_/B _19536_/B VGND VGND VPWR VPWR _19562_/X sky130_fd_sc_hd__and2_4
XFILLER_93_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16774_ _16757_/X _16774_/B _16774_/C VGND VGND VPWR VPWR _16778_/B sky130_fd_sc_hd__and3_4
XANTENNA__12012__A _16143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13986_ _13986_/A _13986_/B _13985_/X VGND VGND VPWR VPWR _13987_/B sky130_fd_sc_hd__or3_4
XFILLER_46_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18513_ _18435_/X _18511_/X _20053_/A _18512_/X VGND VGND VPWR VPWR _24458_/D sky130_fd_sc_hd__a2bb2o_4
X_15725_ _15725_/A _15725_/B VGND VGND VPWR VPWR _15726_/C sky130_fd_sc_hd__or2_4
X_12937_ _12937_/A VGND VGND VPWR VPWR _12974_/A sky130_fd_sc_hd__buf_2
X_19493_ _19419_/A VGND VGND VPWR VPWR _19493_/X sky130_fd_sc_hd__buf_2
XANTENNA__16379__A1 _16302_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12947__A _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16419__A _16121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21372__B2 _21366_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11851__A _13491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18444_ _18390_/A _18444_/B _18442_/X _18444_/D VGND VGND VPWR VPWR _18445_/A sky130_fd_sc_hd__or4_4
X_15656_ _12286_/X _15656_/B VGND VGND VPWR VPWR _15657_/C sky130_fd_sc_hd__or2_4
X_12868_ _12868_/A _23667_/Q VGND VGND VPWR VPWR _12870_/B sky130_fd_sc_hd__or2_4
X_14607_ _14113_/A _14688_/B VGND VGND VPWR VPWR _14607_/X sky130_fd_sc_hd__or2_4
XANTENNA__11570__B IRQ[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11819_ _11819_/A _23806_/Q VGND VGND VPWR VPWR _11820_/C sky130_fd_sc_hd__or2_4
X_18375_ _18358_/X _18363_/Y _18371_/X _18373_/Y _18374_/X VGND VGND VPWR VPWR _18375_/X
+ sky130_fd_sc_hd__a32o_4
X_15587_ _14379_/A _23723_/Q VGND VGND VPWR VPWR _15588_/C sky130_fd_sc_hd__or2_4
X_12799_ _12799_/A _12799_/B VGND VGND VPWR VPWR _12799_/X sky130_fd_sc_hd__or2_4
XFILLER_72_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18634__A _18418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21124__B2 _21123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17326_ _15249_/X _17120_/A VGND VGND VPWR VPWR _17326_/X sky130_fd_sc_hd__or2_4
X_14538_ _13747_/A _14534_/X _14537_/X VGND VGND VPWR VPWR _14538_/X sky130_fd_sc_hd__or3_4
XANTENNA__21675__A2 _21669_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_2_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17257_ _17256_/X VGND VGND VPWR VPWR _17868_/A sky130_fd_sc_hd__buf_2
XFILLER_31_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13778__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14469_ _12878_/A _14539_/B VGND VGND VPWR VPWR _14469_/X sky130_fd_sc_hd__or2_4
XANTENNA__12682__A _13056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16208_ _16201_/A _16131_/B VGND VGND VPWR VPWR _16208_/X sky130_fd_sc_hd__or2_4
XANTENNA__21995__A _21988_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21427__A2 _21426_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17188_ _13591_/X _17161_/X _15782_/B _17157_/X VGND VGND VPWR VPWR _17188_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22624__B2 _22619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16139_ _16139_/A _24087_/Q VGND VGND VPWR VPWR _16139_/X sky130_fd_sc_hd__or2_4
XFILLER_6_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20938__A1 _20872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23752__CLK _23304_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20938__B2 _20839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19829_ _19829_/A _19829_/B VGND VGND VPWR VPWR _19829_/X sky130_fd_sc_hd__or2_4
XFILLER_96_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13018__A _13041_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22840_ _22840_/A VGND VGND VPWR VPWR HWDATA[19] sky130_fd_sc_hd__inv_2
XFILLER_110_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24108__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21235__A _21247_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22771_ _22754_/X _22773_/B _22770_/Y VGND VGND VPWR VPWR _24102_/D sky130_fd_sc_hd__and3_4
XANTENNA__16329__A _16447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21363__B2 _21359_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21722_ _21560_/X _21719_/X _13791_/B _21716_/X VGND VGND VPWR VPWR _21722_/X sky130_fd_sc_hd__o22a_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21653_ _21526_/X _21648_/X _12660_/B _21652_/X VGND VGND VPWR VPWR _21653_/X sky130_fd_sc_hd__o22a_4
X_24441_ _24277_/CLK _24441_/D HRESETn VGND VGND VPWR VPWR _20379_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_90_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20604_ _18375_/X _20424_/X _20516_/X _20603_/Y VGND VGND VPWR VPWR _20605_/A sky130_fd_sc_hd__a211o_4
X_21584_ _21684_/A _21634_/B _21684_/C _20199_/B VGND VGND VPWR VPWR _21584_/X sky130_fd_sc_hd__or4_4
X_24372_ _23358_/CLK _18893_/X HRESETn VGND VGND VPWR VPWR _24372_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_103_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20535_ _24211_/Q _20512_/X _20534_/X VGND VGND VPWR VPWR _22100_/A sky130_fd_sc_hd__o21a_4
X_23323_ _24059_/CLK _23323_/D VGND VGND VPWR VPWR _16775_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_53_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12592__A _12591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21418__A2 _21412_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20466_ _20422_/X _20844_/B _20286_/X VGND VGND VPWR VPWR _20466_/X sky130_fd_sc_hd__a21o_4
X_23254_ _23313_/CLK _23254_/D VGND VGND VPWR VPWR _12206_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23282__CLK _23314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16999__A _17680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22205_ _22212_/A VGND VGND VPWR VPWR _22205_/X sky130_fd_sc_hd__buf_2
XFILLER_49_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13200__B _13200_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23185_ _23217_/CLK _22539_/X VGND VGND VPWR VPWR _13144_/B sky130_fd_sc_hd__dfxtp_4
X_20397_ _20399_/A VGND VGND VPWR VPWR _20512_/A sky130_fd_sc_hd__buf_2
X_22136_ _20892_/A VGND VGND VPWR VPWR _22136_/X sky130_fd_sc_hd__buf_2
XANTENNA__20314__A _20314_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22067_ _21581_/A VGND VGND VPWR VPWR _22068_/A sky130_fd_sc_hd__buf_2
XANTENNA__15408__A _15431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14312__A _15556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21018_ _20339_/X _21016_/X _24060_/Q _21013_/X VGND VGND VPWR VPWR _24060_/D sky130_fd_sc_hd__o22a_4
XFILLER_59_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13840_ _13847_/A VGND VGND VPWR VPWR _13887_/A sky130_fd_sc_hd__buf_2
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15281__A1 _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14966__B _14899_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13771_ _11799_/A _13771_/B _13771_/C VGND VGND VPWR VPWR _13772_/C sky130_fd_sc_hd__or3_4
X_22969_ _18407_/X _22950_/X VGND VGND VPWR VPWR _22970_/C sky130_fd_sc_hd__or2_4
XFILLER_95_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20157__A2 IRQ[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15510_ _13737_/A _15508_/X _15509_/X VGND VGND VPWR VPWR _15514_/B sky130_fd_sc_hd__and3_4
XANTENNA__15143__A _14143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11671__A _11671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_69_0_HCLK clkbuf_6_34_0_HCLK/X VGND VGND VPWR VPWR _24320_/CLK sky130_fd_sc_hd__clkbuf_1
X_12722_ _12722_/A _24052_/Q VGND VGND VPWR VPWR _12723_/C sky130_fd_sc_hd__or2_4
XFILLER_43_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16490_ _16465_/A _16421_/B VGND VGND VPWR VPWR _16490_/X sky130_fd_sc_hd__or2_4
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15441_ _13631_/A _15441_/B _15440_/X VGND VGND VPWR VPWR _15442_/C sky130_fd_sc_hd__and3_4
X_12653_ _12953_/A _12653_/B VGND VGND VPWR VPWR _12654_/C sky130_fd_sc_hd__or2_4
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21106__B2 _21100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ _12529_/A VGND VGND VPWR VPWR _14995_/A sky130_fd_sc_hd__buf_2
X_18160_ _18160_/A VGND VGND VPWR VPWR _18160_/X sky130_fd_sc_hd__buf_2
XFILLER_106_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ _15334_/A _15372_/B _15372_/C VGND VGND VPWR VPWR _15372_/X sky130_fd_sc_hd__and3_4
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21657__A2 _21655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12605_/A VGND VGND VPWR VPWR _12585_/A sky130_fd_sc_hd__buf_2
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17111_ _19830_/A _17032_/B _12892_/A _17105_/X VGND VGND VPWR VPWR _17111_/X sky130_fd_sc_hd__o22a_4
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _14431_/A _14417_/B VGND VGND VPWR VPWR _14323_/X sky130_fd_sc_hd__or2_4
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ _24420_/Q IRQ[5] _11534_/X VGND VGND VPWR VPWR _11538_/A sky130_fd_sc_hd__a21o_4
X_18091_ _18009_/X _18088_/X _18053_/X _18090_/X VGND VGND VPWR VPWR _18091_/X sky130_fd_sc_hd__o22a_4
XFILLER_32_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17042_ _17042_/A VGND VGND VPWR VPWR _17043_/A sky130_fd_sc_hd__buf_2
X_14254_ _13839_/A VGND VGND VPWR VPWR _14359_/A sky130_fd_sc_hd__buf_2
XANTENNA__22606__B2 _22604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22704__A _22683_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13205_ _13231_/A _13203_/X _13205_/C VGND VGND VPWR VPWR _13211_/B sky130_fd_sc_hd__and3_4
X_14185_ _14197_/A VGND VGND VPWR VPWR _14186_/A sky130_fd_sc_hd__buf_2
XFILLER_98_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21290__B1 _15146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13136_ _13059_/Y _13135_/X VGND VGND VPWR VPWR _13136_/X sky130_fd_sc_hd__or2_4
X_18993_ _18988_/X _18992_/X _18988_/X _24340_/Q VGND VGND VPWR VPWR _18993_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13067_ _13096_/A _13067_/B _13067_/C VGND VGND VPWR VPWR _13072_/B sky130_fd_sc_hd__and3_4
X_17944_ _17899_/X _17905_/Y _17939_/X _17942_/Y _17943_/X VGND VGND VPWR VPWR _17944_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_61_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14222__A _11766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21042__B1 _15556_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12018_ _12022_/A _23102_/Q VGND VGND VPWR VPWR _12020_/B sky130_fd_sc_hd__or2_4
X_17875_ _17874_/X _17630_/X _17871_/A _17578_/X VGND VGND VPWR VPWR _17875_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15037__B _23615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21593__B2 _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19614_ HRDATA[26] VGND VGND VPWR VPWR _20754_/A sky130_fd_sc_hd__buf_2
XFILLER_4_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16826_ _12996_/X _16899_/B _13585_/Y VGND VGND VPWR VPWR _16826_/X sky130_fd_sc_hd__o21a_4
XFILLER_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16757_ _11691_/X VGND VGND VPWR VPWR _16757_/X sky130_fd_sc_hd__buf_2
X_19545_ _19545_/A VGND VGND VPWR VPWR _19551_/A sky130_fd_sc_hd__buf_2
XFILLER_19_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13969_ _13643_/A _13969_/B VGND VGND VPWR VPWR _13971_/B sky130_fd_sc_hd__or2_4
XANTENNA__20148__A2 IRQ[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16149__A _16145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12677__A _12559_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21345__B2 _21301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23155__CLK _23155_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15708_ _12747_/A _15708_/B _15708_/C VGND VGND VPWR VPWR _15708_/X sky130_fd_sc_hd__and3_4
XFILLER_80_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16688_ _16715_/A _16688_/B _16688_/C VGND VGND VPWR VPWR _16688_/X sky130_fd_sc_hd__and3_4
X_19476_ _19422_/X _19475_/X HRDATA[14] _19438_/X VGND VGND VPWR VPWR _19477_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21896__A2 _21894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12396__B _12289_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15639_ _13887_/A _23211_/Q VGND VGND VPWR VPWR _15641_/B sky130_fd_sc_hd__or2_4
X_18427_ _17261_/X _18402_/X _17261_/X _18396_/X VGND VGND VPWR VPWR _18427_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18358_ _18418_/A _18274_/A VGND VGND VPWR VPWR _18358_/X sky130_fd_sc_hd__or2_4
XANTENNA__22845__A1 _12752_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17309_ _14723_/B _17309_/B VGND VGND VPWR VPWR _17309_/X sky130_fd_sc_hd__or2_4
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18289_ _18198_/X _18284_/X _18224_/X _18288_/X VGND VGND VPWR VPWR _18289_/X sky130_fd_sc_hd__o22a_4
XFILLER_11_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20320_ _20447_/A VGND VGND VPWR VPWR _20332_/A sky130_fd_sc_hd__buf_2
XANTENNA__18811__B _12101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20251_ _20622_/A VGND VGND VPWR VPWR _20251_/X sky130_fd_sc_hd__buf_2
XANTENNA__13020__B _13085_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19474__B1 HRDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16612__A _16599_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22722__A1_N _22898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20182_ _19379_/X _16997_/X _19313_/A _20181_/X VGND VGND VPWR VPWR _20183_/A sky130_fd_sc_hd__o22a_4
XANTENNA__21820__A2 _21817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16331__B _16256_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14132__A _11909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23941_ _23973_/CLK _23941_/D VGND VGND VPWR VPWR _14533_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13971__A _12217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23872_ _23840_/CLK _23872_/D VGND VGND VPWR VPWR _23872_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19529__B2 _19528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22823_ _22813_/X _22823_/B VGND VGND VPWR VPWR HWDATA[15] sky130_fd_sc_hd__nor2_4
XFILLER_77_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12587__A _12970_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21336__B2 _21330_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22754_ _22768_/C VGND VGND VPWR VPWR _22754_/X sky130_fd_sc_hd__buf_2
XFILLER_44_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21705_ _21705_/A VGND VGND VPWR VPWR _21705_/X sky130_fd_sc_hd__buf_2
XFILLER_38_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22685_ _20509_/A _22679_/X _12823_/B _22683_/X VGND VGND VPWR VPWR _23092_/D sky130_fd_sc_hd__o22a_4
XFILLER_13_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24424_ _24365_/CLK _18799_/X HRESETn VGND VGND VPWR VPWR _24424_/Q sky130_fd_sc_hd__dfrtp_4
X_21636_ _21636_/A VGND VGND VPWR VPWR _21659_/A sky130_fd_sc_hd__inv_2
XANTENNA__22836__A1 _17504_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24355_ _24321_/CLK _24355_/D HRESETn VGND VGND VPWR VPWR _19089_/A sky130_fd_sc_hd__dfstp_4
X_21567_ _21282_/A VGND VGND VPWR VPWR _21567_/X sky130_fd_sc_hd__buf_2
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13211__A _13211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23306_ _23564_/CLK _23306_/D VGND VGND VPWR VPWR _22320_/A sky130_fd_sc_hd__dfxtp_4
X_20518_ _20518_/A VGND VGND VPWR VPWR _20518_/X sky130_fd_sc_hd__buf_2
X_21498_ _21498_/A VGND VGND VPWR VPWR _21498_/Y sky130_fd_sc_hd__inv_2
X_24286_ _24435_/CLK _19237_/X HRESETn VGND VGND VPWR VPWR _19235_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20449_ _20449_/A VGND VGND VPWR VPWR _20449_/X sky130_fd_sc_hd__buf_2
X_23237_ _23557_/CLK _22450_/X VGND VGND VPWR VPWR _14431_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22064__A2 _22059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19465__B1 HRDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23168_ _23233_/CLK _23168_/D VGND VGND VPWR VPWR _14863_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20044__A _19996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16241__B _23513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11666__A _11665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22119_ _20722_/A VGND VGND VPWR VPWR _22119_/X sky130_fd_sc_hd__buf_2
XANTENNA__15138__A _14136_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15990_ _16097_/A _24088_/Q VGND VGND VPWR VPWR _15991_/C sky130_fd_sc_hd__or2_4
X_23099_ _23515_/CLK _23099_/D VGND VGND VPWR VPWR _23099_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_95_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14042__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14941_ _11708_/A VGND VGND VPWR VPWR _15074_/A sky130_fd_sc_hd__buf_2
XFILLER_88_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21575__B2 _21515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13881__A _13909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17660_ _16985_/A _17653_/B _17654_/Y VGND VGND VPWR VPWR _17660_/X sky130_fd_sc_hd__a21o_4
XFILLER_75_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14872_ _14895_/A _14872_/B VGND VGND VPWR VPWR _14872_/X sky130_fd_sc_hd__or2_4
XFILLER_114_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16611_ _16616_/A _16608_/X _16611_/C VGND VGND VPWR VPWR _16612_/C sky130_fd_sc_hd__and3_4
X_13823_ _15411_/A _13821_/X _13823_/C VGND VGND VPWR VPWR _13827_/B sky130_fd_sc_hd__and3_4
XFILLER_21_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17591_ _18274_/A _17495_/A _17502_/X _17512_/A VGND VGND VPWR VPWR _17591_/X sky130_fd_sc_hd__or4_4
XFILLER_5_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12497__A _13015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21327__B2 _21323_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16542_ _16542_/A _16542_/B _16542_/C VGND VGND VPWR VPWR _16542_/X sky130_fd_sc_hd__or3_4
X_19330_ _19328_/X _18288_/X _19328_/X _24242_/Q VGND VGND VPWR VPWR _19330_/X sky130_fd_sc_hd__a2bb2o_4
X_13754_ _13754_/A _13750_/X _13754_/C VGND VGND VPWR VPWR _13755_/C sky130_fd_sc_hd__or3_4
XFILLER_71_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12705_ _12705_/A _12703_/X _12704_/X VGND VGND VPWR VPWR _12705_/X sky130_fd_sc_hd__and3_4
X_19261_ _19261_/A VGND VGND VPWR VPWR _19261_/Y sky130_fd_sc_hd__inv_2
X_16473_ _13354_/X VGND VGND VPWR VPWR _16473_/X sky130_fd_sc_hd__buf_2
XANTENNA__13105__B _23954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13685_ _13684_/X VGND VGND VPWR VPWR _13685_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18212_ _18212_/A VGND VGND VPWR VPWR _18212_/Y sky130_fd_sc_hd__inv_2
X_15424_ _15424_/A _15424_/B _15423_/X VGND VGND VPWR VPWR _15424_/X sky130_fd_sc_hd__and3_4
XFILLER_19_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12636_ _13118_/A _12625_/X _12635_/X VGND VGND VPWR VPWR _12636_/X sky130_fd_sc_hd__and3_4
X_19192_ _19113_/A _19112_/X _19191_/Y VGND VGND VPWR VPWR _24292_/D sky130_fd_sc_hd__o21a_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16416__B _23610_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18143_ _17812_/X _17976_/Y _17800_/X _17971_/Y VGND VGND VPWR VPWR _18143_/X sky130_fd_sc_hd__o22a_4
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15355_ _13871_/A _15289_/B VGND VGND VPWR VPWR _15355_/X sky130_fd_sc_hd__or2_4
XFILLER_89_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12567_ _12567_/A VGND VGND VPWR VPWR _12568_/A sky130_fd_sc_hd__buf_2
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18912__A _18898_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14306_ _15534_/A _14304_/X _14305_/X VGND VGND VPWR VPWR _14306_/X sky130_fd_sc_hd__and3_4
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11518_ _24333_/Q _11518_/B VGND VGND VPWR VPWR _11519_/B sky130_fd_sc_hd__or2_4
X_18074_ _17962_/A _18071_/X _17836_/A _18073_/X VGND VGND VPWR VPWR _18075_/A sky130_fd_sc_hd__o22a_4
XFILLER_89_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15286_ _14152_/A _15352_/B VGND VGND VPWR VPWR _15286_/X sky130_fd_sc_hd__or2_4
X_12498_ _12497_/X _23317_/Q VGND VGND VPWR VPWR _12502_/B sky130_fd_sc_hd__or2_4
XANTENNA__22434__A _20722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17025_ _17025_/A VGND VGND VPWR VPWR _17467_/B sky130_fd_sc_hd__inv_2
X_14237_ _14183_/A _14237_/B _14236_/X VGND VGND VPWR VPWR _14237_/X sky130_fd_sc_hd__and3_4
XANTENNA__22055__A2 _22052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19456__B1 HRDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12960__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14168_ _15026_/A _23689_/Q VGND VGND VPWR VPWR _14170_/B sky130_fd_sc_hd__or2_4
X_13119_ _13119_/A _13119_/B VGND VGND VPWR VPWR _13119_/X sky130_fd_sc_hd__or2_4
XFILLER_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19743__A _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14099_ _14136_/A _14099_/B _14098_/X VGND VGND VPWR VPWR _14099_/X sky130_fd_sc_hd__or3_4
X_18976_ _18965_/X _18974_/X _18975_/Y _18968_/X VGND VGND VPWR VPWR _18976_/X sky130_fd_sc_hd__o22a_4
X_17927_ _17817_/X _17219_/X _17825_/X _17230_/X VGND VGND VPWR VPWR _17928_/A sky130_fd_sc_hd__o22a_4
XFILLER_85_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18359__A _18295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21566__B2 _21563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13791__A _15429_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17858_ _18189_/A VGND VGND VPWR VPWR _17858_/X sky130_fd_sc_hd__buf_2
XANTENNA__18431__B2 _18430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16809_ _16622_/A _16809_/B _16808_/X VGND VGND VPWR VPWR _16810_/C sky130_fd_sc_hd__or3_4
X_17789_ _17779_/X _17789_/B _17789_/C _17788_/X VGND VGND VPWR VPWR _17790_/A sky130_fd_sc_hd__or4_4
XANTENNA__21318__B2 _21316_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19528_ _19500_/X _19535_/A _19528_/C _19527_/X VGND VGND VPWR VPWR _19528_/X sky130_fd_sc_hd__and4_4
XFILLER_81_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_52_0_HCLK clkbuf_6_26_0_HCLK/X VGND VGND VPWR VPWR _23915_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19459_ _19433_/Y VGND VGND VPWR VPWR _19459_/X sky130_fd_sc_hd__buf_2
XANTENNA__20541__A2 _20405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16607__A _11821_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22470_ _22464_/Y _22469_/X _22388_/X _22469_/X VGND VGND VPWR VPWR _22470_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16326__B _16266_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21421_ _21249_/X _21419_/X _13112_/B _21416_/X VGND VGND VPWR VPWR _23826_/D sky130_fd_sc_hd__o22a_4
XFILLER_13_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22294__A2 _22293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14127__A _14119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13031__A _13031_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21352_ _21359_/A VGND VGND VPWR VPWR _21352_/X sky130_fd_sc_hd__buf_2
X_24140_ _24229_/CLK _19960_/Y HRESETn VGND VGND VPWR VPWR _24140_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22344__A _22344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20303_ _20525_/A VGND VGND VPWR VPWR _20303_/X sky130_fd_sc_hd__buf_2
XFILLER_30_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13966__A _13966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21283_ _21271_/A VGND VGND VPWR VPWR _21283_/X sky130_fd_sc_hd__buf_2
X_24071_ _23368_/CLK _20820_/X VGND VGND VPWR VPWR _24071_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22046__A2 _22045_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16342__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12870__A _12870_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20234_ _17083_/A _16910_/X _16913_/X _11591_/C VGND VGND VPWR VPWR _20235_/A sky130_fd_sc_hd__or4_4
X_23022_ _18124_/X _23017_/B VGND VGND VPWR VPWR _23023_/C sky130_fd_sc_hd__or2_4
XANTENNA__19998__A1 _19994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19998__B2 _19997_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20165_ _24442_/Q IRQ[27] _20164_/X VGND VGND VPWR VPWR _20165_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_118_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18670__A1 _18142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20799__A HRDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20096_ NMI VGND VGND VPWR VPWR _20105_/A sky130_fd_sc_hd__inv_2
XANTENNA__21557__B2 _21551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23924_ _23315_/CLK _23924_/D VGND VGND VPWR VPWR _23924_/Q sky130_fd_sc_hd__dfxtp_4
X_23855_ _23859_/CLK _23855_/D VGND VGND VPWR VPWR _23855_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22806_ _22792_/X _22806_/B VGND VGND VPWR VPWR HWDATA[10] sky130_fd_sc_hd__nor2_4
XANTENNA__13206__A _12383_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11652__C _12965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23786_ _23692_/CLK _21483_/X VGND VGND VPWR VPWR _23786_/Q sky130_fd_sc_hd__dfxtp_4
X_20998_ _20283_/X _20989_/Y _20996_/X _20997_/Y _20459_/A VGND VGND VPWR VPWR _20998_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22519__A _22518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21423__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19922__B2 _20576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22737_ _22736_/Y _24097_/Q _22736_/Y _24097_/Q VGND VGND VPWR VPWR _22737_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13470_ _13450_/A _23823_/Q VGND VGND VPWR VPWR _13471_/C sky130_fd_sc_hd__or2_4
X_22668_ _22683_/A VGND VGND VPWR VPWR _22668_/X sky130_fd_sc_hd__buf_2
XFILLER_16_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12421_ _12421_/A VGND VGND VPWR VPWR _12967_/A sky130_fd_sc_hd__buf_2
X_24407_ _24277_/CLK _24407_/D HRESETn VGND VGND VPWR VPWR _20426_/A sky130_fd_sc_hd__dfrtp_4
X_21619_ _21590_/A VGND VGND VPWR VPWR _21619_/X sky130_fd_sc_hd__buf_2
XFILLER_16_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22285__A2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22599_ _22437_/X _22593_/X _14025_/B _22597_/X VGND VGND VPWR VPWR _23146_/D sky130_fd_sc_hd__o22a_4
XFILLER_21_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15140_ _14096_/X _15210_/B VGND VGND VPWR VPWR _15140_/X sky130_fd_sc_hd__or2_4
X_12352_ _12381_/A _12224_/B VGND VGND VPWR VPWR _12352_/X sky130_fd_sc_hd__or2_4
X_24338_ _23358_/CLK _19006_/X HRESETn VGND VGND VPWR VPWR _24338_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22254__A _22269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15071_ _11723_/A _15069_/X _15071_/C VGND VGND VPWR VPWR _15077_/B sky130_fd_sc_hd__and3_4
X_12283_ _13025_/A VGND VGND VPWR VPWR _15688_/A sky130_fd_sc_hd__buf_2
X_24269_ _24365_/CLK _24269_/D HRESETn VGND VGND VPWR VPWR _19218_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12780__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14022_ _14045_/A _23562_/Q VGND VGND VPWR VPWR _14023_/C sky130_fd_sc_hd__or2_4
XANTENNA__21245__B1 _23924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21796__B2 _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18830_ _17164_/X _18827_/X _24408_/Q _18828_/X VGND VGND VPWR VPWR _24408_/D sky130_fd_sc_hd__o22a_4
XFILLER_27_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15973_ _11852_/X _15942_/X _15954_/X _15963_/X _15972_/X VGND VGND VPWR VPWR _15973_/X
+ sky130_fd_sc_hd__a32o_4
X_18761_ _11844_/X _18866_/B _11620_/X _18812_/C VGND VGND VPWR VPWR _18761_/X sky130_fd_sc_hd__or4_4
XFILLER_96_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18179__A _18297_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14924_ _12582_/A _14860_/B VGND VGND VPWR VPWR _14925_/C sky130_fd_sc_hd__or2_4
X_17712_ _16970_/A _17393_/X VGND VGND VPWR VPWR _17712_/X sky130_fd_sc_hd__and2_4
X_18692_ _17327_/X _18693_/B VGND VGND VPWR VPWR _18692_/X sky130_fd_sc_hd__or2_4
X_14855_ _14855_/A VGND VGND VPWR VPWR _14855_/Y sky130_fd_sc_hd__inv_2
X_17643_ _17766_/A _17274_/Y VGND VGND VPWR VPWR _17946_/B sky130_fd_sc_hd__nand2_4
XFILLER_64_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13806_ _13682_/A _13783_/X _13790_/X _13797_/X _13805_/X VGND VGND VPWR VPWR _13806_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17574_ _16374_/X _17549_/B VGND VGND VPWR VPWR _17574_/Y sky130_fd_sc_hd__nand2_4
X_14786_ _14785_/X VGND VGND VPWR VPWR _14786_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12020__A _12020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11998_ _11998_/A _11998_/B _11998_/C VGND VGND VPWR VPWR _11999_/C sky130_fd_sc_hd__and3_4
XFILLER_95_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16525_ _15928_/X _16520_/X _16524_/Y VGND VGND VPWR VPWR _16525_/X sky130_fd_sc_hd__o21a_4
X_19313_ _19313_/A VGND VGND VPWR VPWR _19313_/X sky130_fd_sc_hd__buf_2
X_13737_ _13737_/A _13737_/B _13737_/C VGND VGND VPWR VPWR _13738_/C sky130_fd_sc_hd__and3_4
XANTENNA__19913__B2 _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_39_0_HCLK clkbuf_6_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_78_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12955__A _12955_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21720__B2 _21716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15331__A _13991_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16456_ _11715_/A _16388_/B VGND VGND VPWR VPWR _16456_/X sky130_fd_sc_hd__or2_4
X_19244_ _19231_/A _19245_/A _19243_/Y VGND VGND VPWR VPWR _24282_/D sky130_fd_sc_hd__o21a_4
X_13668_ _15436_/A _23464_/Q VGND VGND VPWR VPWR _13670_/B sky130_fd_sc_hd__or2_4
XFILLER_38_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15407_ _13630_/A _15407_/B VGND VGND VPWR VPWR _15407_/X sky130_fd_sc_hd__or2_4
X_12619_ _12650_/A VGND VGND VPWR VPWR _12660_/A sky130_fd_sc_hd__buf_2
X_19175_ _19122_/B VGND VGND VPWR VPWR _19175_/Y sky130_fd_sc_hd__inv_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16387_ _15999_/X _16387_/B VGND VGND VPWR VPWR _16387_/X sky130_fd_sc_hd__or2_4
X_13599_ _14782_/A VGND VGND VPWR VPWR _13600_/A sky130_fd_sc_hd__buf_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20287__A1 _20285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18126_ _17762_/X _17660_/X _17762_/X _17660_/X VGND VGND VPWR VPWR _18126_/X sky130_fd_sc_hd__a2bb2o_4
X_15338_ _14008_/A _15338_/B _15338_/C VGND VGND VPWR VPWR _15346_/B sky130_fd_sc_hd__or3_4
XANTENNA__15985__B _23416_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18057_ _17888_/X _18055_/X _19981_/A _18056_/X VGND VGND VPWR VPWR _24473_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13786__A _12450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15269_ _14158_/A _15269_/B VGND VGND VPWR VPWR _15269_/X sky130_fd_sc_hd__or2_4
XANTENNA__12690__A _12221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17008_ _17024_/C _17030_/B _17024_/A _17024_/B VGND VGND VPWR VPWR _17072_/A sky130_fd_sc_hd__or4_4
XFILLER_28_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21508__A _21532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18959_ _18959_/A VGND VGND VPWR VPWR _18959_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17705__B _17404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18404__A1 _18216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15506__A _13097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21970_ _21985_/A VGND VGND VPWR VPWR _21970_/X sky130_fd_sc_hd__buf_2
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20921_ _20841_/X _20920_/X VGND VGND VPWR VPWR _20921_/X sky130_fd_sc_hd__and2_4
XFILLER_27_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13026__A _13026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23640_ _23316_/CLK _21749_/X VGND VGND VPWR VPWR _23640_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20852_ _19699_/Y _20851_/X _20844_/B _20821_/B VGND VGND VPWR VPWR _20852_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22339__A _22368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19904__A1 _24157_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23571_ _23859_/CLK _21888_/X VGND VGND VPWR VPWR _12943_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20783_ _20642_/X _20781_/X _20783_/C VGND VGND VPWR VPWR _20783_/X sky130_fd_sc_hd__and3_4
XFILLER_23_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12865__A _12865_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20514__A2 _20895_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16337__A _13415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21711__B2 _21709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22522_ _22536_/A VGND VGND VPWR VPWR _22522_/X sky130_fd_sc_hd__buf_2
XFILLER_23_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16056__B _15984_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22453_ _22451_/X _22452_/X _14569_/B _22447_/X VGND VGND VPWR VPWR _23236_/D sky130_fd_sc_hd__o22a_4
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22267__A2 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21404_ _21400_/A VGND VGND VPWR VPWR _21419_/A sky130_fd_sc_hd__buf_2
XANTENNA__15895__B _15839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22384_ _22384_/A VGND VGND VPWR VPWR _22384_/X sky130_fd_sc_hd__buf_2
XANTENNA__24463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24123_ _24126_/CLK _20041_/Y HRESETn VGND VGND VPWR VPWR _24123_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13696__A _13695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21335_ _21273_/X _21333_/X _13651_/B _21330_/X VGND VGND VPWR VPWR _23880_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16072__A _16072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24054_ _23316_/CLK _21026_/X VGND VGND VPWR VPWR _24054_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21266_ _21242_/A VGND VGND VPWR VPWR _21266_/X sky130_fd_sc_hd__buf_2
XFILLER_89_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23836__CLK _23840_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21778__B2 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14304__B _14304_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23005_ _22989_/A _23005_/B _23005_/C VGND VGND VPWR VPWR _23005_/X sky130_fd_sc_hd__and3_4
XFILLER_46_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20217_ _20218_/A HRDATA[31] VGND VGND VPWR VPWR _20217_/X sky130_fd_sc_hd__or2_4
X_21197_ _21168_/A VGND VGND VPWR VPWR _21197_/X sky130_fd_sc_hd__buf_2
XFILLER_46_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16800__A _16800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20148_ _20966_/A IRQ[1] _11541_/Y _24418_/Q IRQ[3] VGND VGND VPWR VPWR _20148_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20450__B2 _20449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20322__A _20494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15416__A _15443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12970_ _12970_/A _12970_/B _12969_/X VGND VGND VPWR VPWR _12971_/C sky130_fd_sc_hd__and3_4
X_20079_ _20079_/A VGND VGND VPWR VPWR _20079_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11921_ _11901_/X VGND VGND VPWR VPWR _11921_/X sky130_fd_sc_hd__buf_2
X_23907_ _23907_/CLK _23907_/D VGND VGND VPWR VPWR _14802_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_66_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21950__B2 _21949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14640_ _11841_/A _13595_/A _14606_/X _11594_/A _14639_/X VGND VGND VPWR VPWR _14640_/X
+ sky130_fd_sc_hd__a32o_4
X_11852_ _11851_/X VGND VGND VPWR VPWR _11852_/X sky130_fd_sc_hd__buf_2
X_23838_ _23320_/CLK _21403_/X VGND VGND VPWR VPWR _23838_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14974__B _23840_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14571_ _14108_/A _14569_/X _14571_/C VGND VGND VPWR VPWR _14578_/B sky130_fd_sc_hd__and3_4
X_11783_ _11747_/X _11776_/X _11782_/X VGND VGND VPWR VPWR _11783_/X sky130_fd_sc_hd__or3_4
X_23769_ _23770_/CLK _23769_/D VGND VGND VPWR VPWR _16249_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16310_ _11713_/X VGND VGND VPWR VPWR _16323_/A sky130_fd_sc_hd__buf_2
X_13522_ _13522_/A _13522_/B _13521_/X VGND VGND VPWR VPWR _13528_/B sky130_fd_sc_hd__and3_4
X_17290_ _17290_/A _17413_/B VGND VGND VPWR VPWR _17290_/X sky130_fd_sc_hd__or2_4
XFILLER_70_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16241_ _16150_/A _23513_/Q VGND VGND VPWR VPWR _16241_/X sky130_fd_sc_hd__or2_4
X_13453_ _12462_/A _13453_/B VGND VGND VPWR VPWR _13453_/X sky130_fd_sc_hd__or2_4
XANTENNA__14990__A _14990_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12404_ _12419_/A _12298_/B VGND VGND VPWR VPWR _12404_/X sky130_fd_sc_hd__or2_4
XFILLER_70_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16172_ _16203_/A _16170_/X _16171_/X VGND VGND VPWR VPWR _16172_/X sky130_fd_sc_hd__and3_4
X_13384_ _13351_/X _13384_/B _13384_/C VGND VGND VPWR VPWR _13389_/B sky130_fd_sc_hd__and3_4
XANTENNA__17134__A1 _15251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18331__B1 _18082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15123_ _15051_/X _15119_/X _15122_/X VGND VGND VPWR VPWR _15123_/Y sky130_fd_sc_hd__o21ai_4
X_12335_ _11850_/A _12334_/X VGND VGND VPWR VPWR _12335_/X sky130_fd_sc_hd__and2_4
XFILLER_115_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18882__A1 _17277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20216__B _20445_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15054_ _14046_/A _15054_/B _15053_/X VGND VGND VPWR VPWR _15054_/X sky130_fd_sc_hd__and3_4
X_19931_ _19925_/X _19931_/B VGND VGND VPWR VPWR _19931_/X sky130_fd_sc_hd__and2_4
X_12266_ _13957_/A VGND VGND VPWR VPWR _14128_/A sky130_fd_sc_hd__buf_2
X_14005_ _14065_/A _14001_/X _14005_/C VGND VGND VPWR VPWR _14005_/X sky130_fd_sc_hd__and3_4
XFILLER_68_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19862_ _19862_/A VGND VGND VPWR VPWR _19862_/Y sky130_fd_sc_hd__inv_2
X_12197_ _13677_/A VGND VGND VPWR VPWR _13631_/A sky130_fd_sc_hd__buf_2
XANTENNA__12015__A _16536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16710__A _11936_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18813_ _18813_/A VGND VGND VPWR VPWR _18813_/X sky130_fd_sc_hd__buf_2
X_19793_ _19793_/A _19793_/B VGND VGND VPWR VPWR _19793_/X sky130_fd_sc_hd__or2_4
XFILLER_1_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11854__A _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18744_ _19943_/B _18743_/X VGND VGND VPWR VPWR _18744_/X sky130_fd_sc_hd__or2_4
X_15956_ _15956_/A VGND VGND VPWR VPWR _15957_/A sky130_fd_sc_hd__buf_2
XANTENNA__22194__B2 _22190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14907_ _14991_/A _14905_/X _14907_/C VGND VGND VPWR VPWR _14907_/X sky130_fd_sc_hd__and3_4
X_15887_ _15892_/A _15825_/B VGND VGND VPWR VPWR _15887_/X sky130_fd_sc_hd__or2_4
X_18675_ _18499_/X _17322_/X _18206_/A VGND VGND VPWR VPWR _18675_/X sky130_fd_sc_hd__a21o_4
XFILLER_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20744__A2 _20730_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21941__B2 _21935_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17626_ _17461_/X _17626_/B _17626_/C _17626_/D VGND VGND VPWR VPWR _18081_/B sky130_fd_sc_hd__and4_4
XFILLER_36_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14838_ _14845_/A _14780_/B VGND VGND VPWR VPWR _14839_/C sky130_fd_sc_hd__or2_4
XFILLER_24_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21063__A _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14769_ _15413_/A _14769_/B VGND VGND VPWR VPWR _14769_/X sky130_fd_sc_hd__or2_4
X_17557_ _17556_/X VGND VGND VPWR VPWR _17558_/B sky130_fd_sc_hd__inv_2
XANTENNA__12685__A _15654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16508_ _16159_/X _16508_/B VGND VGND VPWR VPWR _16509_/C sky130_fd_sc_hd__or2_4
X_17488_ _13350_/Y _17013_/A _17021_/A _17487_/X VGND VGND VPWR VPWR _17488_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18570__B1 _18565_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19227_ _24278_/Q _19226_/X VGND VGND VPWR VPWR _19251_/A sky130_fd_sc_hd__and2_4
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15996__A _15959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16439_ _13447_/X _16437_/X _16439_/C VGND VGND VPWR VPWR _16440_/C sky130_fd_sc_hd__and3_4
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22249__A2 _22222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21457__B1 _23805_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19158_ _24309_/Q _19129_/X _19157_/Y VGND VGND VPWR VPWR _19158_/X sky130_fd_sc_hd__o21a_4
XANTENNA__20407__A _20407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18109_ _17914_/X _17919_/Y _17910_/X _17916_/Y VGND VGND VPWR VPWR _18109_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19089_ _19089_/A VGND VGND VPWR VPWR _19089_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20126__B _20125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21209__B1 _14889_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21120_ _20315_/X _21119_/X _23997_/Q _21116_/X VGND VGND VPWR VPWR _21120_/X sky130_fd_sc_hd__o22a_4
XFILLER_86_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22622__A _22636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21051_ _21015_/A VGND VGND VPWR VPWR _21051_/X sky130_fd_sc_hd__buf_2
XFILLER_113_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22421__A2 _22416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18625__B2 _18624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20002_ _18196_/X _19985_/X _20001_/Y _19996_/X VGND VGND VPWR VPWR _20002_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20432__A1 _20293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20142__A IRQ[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14140__A _14318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22185__B2 _22183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23239__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21953_ _21840_/X _21952_/X _23529_/Q _21949_/X VGND VGND VPWR VPWR _23529_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21932__B2 _21928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20904_ _20903_/X VGND VGND VPWR VPWR _20904_/Y sky130_fd_sc_hd__inv_2
X_21884_ _21884_/A VGND VGND VPWR VPWR _21884_/X sky130_fd_sc_hd__buf_2
XFILLER_55_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24366__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _23336_/CLK _21772_/X VGND VGND VPWR VPWR _13825_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_110_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ _20634_/A _20834_/X VGND VGND VPWR VPWR _20835_/Y sky130_fd_sc_hd__nand2_4
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12595__A _12640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22488__A2 _22486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19889__B1 _19888_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20499__A1 _20494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23554_ _23812_/CLK _23554_/D VGND VGND VPWR VPWR _15274_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_22_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_22_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20766_ _20704_/X _20765_/Y _24265_/Q _20562_/X VGND VGND VPWR VPWR _20766_/X sky130_fd_sc_hd__o22a_4
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21160__A2 _21133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22505_ _22446_/X _22500_/X _14417_/B _22504_/X VGND VGND VPWR VPWR _23206_/D sky130_fd_sc_hd__o22a_4
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23485_ _23485_/CLK _23485_/D VGND VGND VPWR VPWR _23485_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20697_ _21263_/A VGND VGND VPWR VPWR _20697_/X sky130_fd_sc_hd__buf_2
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22436_ _22434_/X _22428_/X _15522_/B _22435_/X VGND VGND VPWR VPWR _23243_/D sky130_fd_sc_hd__o22a_4
XFILLER_104_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20317__A _18759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11939__A _11921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22367_ _22122_/X _22361_/X _13939_/B _22365_/X VGND VGND VPWR VPWR _23274_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22660__A2 _22657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14315__A _14315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12120_ _12153_/A _23517_/Q VGND VGND VPWR VPWR _12120_/X sky130_fd_sc_hd__or2_4
X_24106_ _24230_/CLK _24106_/D HRESETn VGND VGND VPWR VPWR _19430_/B sky130_fd_sc_hd__dfrtp_4
X_21318_ _21244_/X _21312_/X _23892_/Q _21316_/X VGND VGND VPWR VPWR _21318_/X sky130_fd_sc_hd__o22a_4
X_22298_ _22145_/X _22293_/X _14859_/B _22262_/A VGND VGND VPWR VPWR _22298_/X sky130_fd_sc_hd__o22a_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12051_ _11999_/A VGND VGND VPWR VPWR _12051_/X sky130_fd_sc_hd__buf_2
X_24037_ _23365_/CLK _21050_/X VGND VGND VPWR VPWR _14536_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21249_ _21249_/A VGND VGND VPWR VPWR _21249_/X sky130_fd_sc_hd__buf_2
XFILLER_105_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22412__A2 _22404_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16887__D _16886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15810_ _12890_/A _15810_/B _15810_/C VGND VGND VPWR VPWR _15811_/C sky130_fd_sc_hd__and3_4
XFILLER_77_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15146__A _15146_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16790_ _11782_/A _16788_/X _16790_/C VGND VGND VPWR VPWR _16790_/X sky130_fd_sc_hd__and3_4
XANTENNA__14050__A _14050_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18919__A2 _18891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15741_ _12792_/A _15669_/B VGND VGND VPWR VPWR _15741_/X sky130_fd_sc_hd__or2_4
XFILLER_98_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12953_ _12953_/A _12953_/B VGND VGND VPWR VPWR _12953_/X sky130_fd_sc_hd__or2_4
XANTENNA__14985__A _11798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_104_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR _23122_/CLK sky130_fd_sc_hd__clkbuf_1
X_11904_ _11875_/X _11904_/B _11904_/C VGND VGND VPWR VPWR _11904_/X sky130_fd_sc_hd__and3_4
XFILLER_59_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15672_ _15695_/A _15668_/X _15671_/X VGND VGND VPWR VPWR _15672_/X sky130_fd_sc_hd__or3_4
X_18460_ _16973_/B VGND VGND VPWR VPWR _18460_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12884_ _13608_/A VGND VGND VPWR VPWR _12885_/A sky130_fd_sc_hd__buf_2
XFILLER_61_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14623_ _15036_/A VGND VGND VPWR VPWR _14758_/A sky130_fd_sc_hd__buf_2
X_17411_ _14174_/X VGND VGND VPWR VPWR _17411_/Y sky130_fd_sc_hd__inv_2
X_11835_ _11675_/X _11835_/B _11834_/X VGND VGND VPWR VPWR _11836_/C sky130_fd_sc_hd__and3_4
X_18391_ _18390_/X VGND VGND VPWR VPWR _18391_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17342_/A VGND VGND VPWR VPWR _17364_/A sky130_fd_sc_hd__inv_2
X_14554_ _14554_/A _14476_/B VGND VGND VPWR VPWR _14554_/X sky130_fd_sc_hd__or2_4
X_11766_ _11766_/A VGND VGND VPWR VPWR _13901_/A sky130_fd_sc_hd__buf_2
XANTENNA__17355__A1 _15453_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17355__B2 _17354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22707__A _22671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24385__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13500_/X _13502_/X _13505_/C VGND VGND VPWR VPWR _13505_/X sky130_fd_sc_hd__and3_4
XFILLER_105_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17273_ _17273_/A _17561_/B VGND VGND VPWR VPWR _17273_/X sky130_fd_sc_hd__and2_4
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _15404_/A _14483_/X _14484_/X VGND VGND VPWR VPWR _14485_/X sky130_fd_sc_hd__and3_4
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11697_ _11697_/A VGND VGND VPWR VPWR _12383_/A sky130_fd_sc_hd__buf_2
XFILLER_105_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16705__A _11903_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16224_ _16193_/A _24087_/Q VGND VGND VPWR VPWR _16225_/C sky130_fd_sc_hd__or2_4
X_19012_ _19002_/X _19011_/X _19002_/X _24337_/Q VGND VGND VPWR VPWR _19012_/X sky130_fd_sc_hd__a2bb2o_4
X_13436_ _11913_/X _13434_/X _13436_/C VGND VGND VPWR VPWR _13436_/X sky130_fd_sc_hd__and3_4
XANTENNA__17107__A1 _14786_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17107__B2 _17106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16424__B _16424_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16155_ _11843_/X _11619_/X _16123_/X _11597_/X _16154_/X VGND VGND VPWR VPWR _16155_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11849__A _13056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13367_ _13358_/X _24016_/Q VGND VGND VPWR VPWR _13369_/B sky130_fd_sc_hd__or2_4
XFILLER_6_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22651__A2 _22650_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15106_ _11710_/A _23839_/Q VGND VGND VPWR VPWR _15107_/C sky130_fd_sc_hd__or2_4
X_12318_ _12196_/A VGND VGND VPWR VPWR _14322_/A sky130_fd_sc_hd__buf_2
X_16086_ _16109_/A _16084_/X _16086_/C VGND VGND VPWR VPWR _16086_/X sky130_fd_sc_hd__and3_4
X_13298_ _12914_/A _13293_/X _13298_/C VGND VGND VPWR VPWR _13298_/X sky130_fd_sc_hd__or3_4
XANTENNA__22442__A _22127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15037_ _15037_/A _23615_/Q VGND VGND VPWR VPWR _15038_/C sky130_fd_sc_hd__or2_4
X_19914_ _19909_/X _24149_/Q _19910_/X _20445_/B VGND VGND VPWR VPWR _24149_/D sky130_fd_sc_hd__o22a_4
X_12249_ _12695_/A _12246_/X _12248_/X VGND VGND VPWR VPWR _12249_/X sky130_fd_sc_hd__and3_4
XFILLER_68_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16440__A _11861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14879__B _14879_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19845_ _19541_/B _19835_/X _19445_/A _19876_/B VGND VGND VPWR VPWR _19845_/X sky130_fd_sc_hd__a211o_4
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19751__A HRDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19776_ _19775_/Y _19629_/A VGND VGND VPWR VPWR _19776_/X sky130_fd_sc_hd__and2_4
XFILLER_68_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16988_ _17645_/A _17894_/D VGND VGND VPWR VPWR _16988_/X sky130_fd_sc_hd__or2_4
XFILLER_7_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18727_ _17221_/Y _17100_/X VGND VGND VPWR VPWR _18727_/X sky130_fd_sc_hd__or2_4
X_15939_ _15939_/A _23352_/Q VGND VGND VPWR VPWR _15941_/B sky130_fd_sc_hd__or2_4
XFILLER_114_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21914__B2 _21869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18658_ _18658_/A _18657_/X VGND VGND VPWR VPWR _18658_/X sky130_fd_sc_hd__or2_4
XFILLER_91_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17609_ _17322_/X VGND VGND VPWR VPWR _17609_/Y sky130_fd_sc_hd__inv_2
X_18589_ _18216_/A _18118_/X VGND VGND VPWR VPWR _18589_/Y sky130_fd_sc_hd__nor2_4
X_20620_ _20285_/X HRDATA[15] _20226_/B _20619_/X VGND VGND VPWR VPWR _20620_/X sky130_fd_sc_hd__a211o_4
XANTENNA__21678__B1 _14779_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22617__A _22621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21142__A2 _21140_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23681__CLK _23819_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20551_ _24210_/Q _20512_/X _20550_/Y VGND VGND VPWR VPWR _20552_/A sky130_fd_sc_hd__o21a_4
X_23270_ _23270_/CLK _23270_/D VGND VGND VPWR VPWR _14279_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_118_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19099__A1 _18965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20482_ _20376_/X _20466_/X _20288_/X _20481_/Y VGND VGND VPWR VPWR _20482_/X sky130_fd_sc_hd__a211o_4
XFILLER_118_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22221_ _22098_/X _22215_/X _23380_/Q _22219_/X VGND VGND VPWR VPWR _22221_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11759__A _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18846__A1 _17191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19926__A _12101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22642__A2 _22636_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22152_ _22151_/X VGND VGND VPWR VPWR _22153_/A sky130_fd_sc_hd__buf_2
XFILLER_82_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21103_ _21067_/A VGND VGND VPWR VPWR _21103_/X sky130_fd_sc_hd__buf_2
XANTENNA__13974__A _12209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17446__A _12992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22083_ _20372_/A VGND VGND VPWR VPWR _22083_/X sky130_fd_sc_hd__buf_2
XANTENNA__16350__A _16364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21034_ _21027_/A VGND VGND VPWR VPWR _21034_/X sky130_fd_sc_hd__buf_2
XANTENNA__24187__CLK _24187_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20956__A2 _20873_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22985_ _22985_/A VGND VGND VPWR VPWR _22985_/X sky130_fd_sc_hd__buf_2
XFILLER_83_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17181__A _12841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21936_ _21811_/X _21931_/X _12633_/B _21935_/X VGND VGND VPWR VPWR _23541_/D sky130_fd_sc_hd__o22a_4
XFILLER_3_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21381__A2 _21376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15413__B _23916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21867_ _21866_/X VGND VGND VPWR VPWR _21901_/A sky130_fd_sc_hd__buf_2
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11619_/X VGND VGND VPWR VPWR _11620_/X sky130_fd_sc_hd__buf_2
X_23606_ _24084_/CLK _21810_/X VGND VGND VPWR VPWR _12289_/B sky130_fd_sc_hd__dfxtp_4
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20818_ _22129_/A VGND VGND VPWR VPWR _20819_/A sky130_fd_sc_hd__buf_2
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21798_ _21797_/X _21793_/X _23611_/Q _21788_/X VGND VGND VPWR VPWR _23611_/D sky130_fd_sc_hd__o22a_4
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _20656_/A IRQ[14] VGND VGND VPWR VPWR _11551_/X sky130_fd_sc_hd__and2_4
X_23537_ _23155_/CLK _23537_/D VGND VGND VPWR VPWR _23537_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20749_ _20613_/X _20748_/X _24074_/Q _20724_/X VGND VGND VPWR VPWR _24074_/D sky130_fd_sc_hd__o22a_4
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _12320_/A _14268_/X _14270_/C VGND VGND VPWR VPWR _14270_/X sky130_fd_sc_hd__and3_4
XFILLER_17_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23468_ _23794_/CLK _22048_/X VGND VGND VPWR VPWR _23468_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16244__B _16244_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13221_ _13239_/A _23569_/Q VGND VGND VPWR VPWR _13222_/C sky130_fd_sc_hd__or2_4
X_22419_ _22418_/X _22416_/X _13064_/B _22411_/X VGND VGND VPWR VPWR _22419_/X sky130_fd_sc_hd__o22a_4
XFILLER_10_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18837__A1 _12990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11669__A _11669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23399_ _23591_/CLK _22189_/X VGND VGND VPWR VPWR _23399_/Q sky130_fd_sc_hd__dfxtp_4
X_13152_ _13055_/A VGND VGND VPWR VPWR _15695_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_29_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR _23584_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22262__A _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12103_ _12098_/A _23645_/Q VGND VGND VPWR VPWR _12104_/C sky130_fd_sc_hd__or2_4
X_13083_ _13083_/A _13072_/X _13083_/C VGND VGND VPWR VPWR _13103_/B sky130_fd_sc_hd__and3_4
X_17960_ _17960_/A VGND VGND VPWR VPWR _17960_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22397__B2 _22387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12034_ _12034_/A _12033_/X VGND VGND VPWR VPWR _12035_/A sky130_fd_sc_hd__or2_4
X_16911_ _16910_/X _16916_/B _16903_/X VGND VGND VPWR VPWR _16911_/X sky130_fd_sc_hd__o21a_4
X_17891_ _18342_/A _17891_/B VGND VGND VPWR VPWR _17896_/A sky130_fd_sc_hd__or2_4
XFILLER_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19630_ _19630_/A _19599_/B VGND VGND VPWR VPWR _19867_/B sky130_fd_sc_hd__or2_4
X_16842_ _14267_/B _16841_/X _14265_/A VGND VGND VPWR VPWR _16842_/X sky130_fd_sc_hd__o21a_4
XFILLER_78_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23554__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19561_ _19561_/A VGND VGND VPWR VPWR _19784_/B sky130_fd_sc_hd__buf_2
XFILLER_20_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13985_ _13985_/A _13985_/B _13985_/C VGND VGND VPWR VPWR _13985_/X sky130_fd_sc_hd__and3_4
X_16773_ _16773_/A _23995_/Q VGND VGND VPWR VPWR _16774_/C sky130_fd_sc_hd__or2_4
XFILLER_98_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18187__A _17259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18512_ _18381_/A VGND VGND VPWR VPWR _18512_/X sky130_fd_sc_hd__buf_2
X_12936_ _12949_/A _24019_/Q VGND VGND VPWR VPWR _12939_/B sky130_fd_sc_hd__or2_4
X_15724_ _15724_/A _15724_/B VGND VGND VPWR VPWR _15726_/B sky130_fd_sc_hd__or2_4
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19492_ _19491_/X VGND VGND VPWR VPWR _19492_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17576__A1 _17144_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16379__A2 _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21372__A2 _21369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18443_ _18443_/A _17361_/A VGND VGND VPWR VPWR _18444_/D sky130_fd_sc_hd__and2_4
XANTENNA__15323__B _15260_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12867_ _12528_/A _12859_/X _12867_/C VGND VGND VPWR VPWR _12867_/X sky130_fd_sc_hd__or3_4
X_15655_ _12284_/X _15655_/B VGND VGND VPWR VPWR _15657_/B sky130_fd_sc_hd__or2_4
XFILLER_34_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11818_ _11818_/A _23102_/Q VGND VGND VPWR VPWR _11820_/B sky130_fd_sc_hd__or2_4
X_14606_ _15450_/A _14578_/X _14587_/X _14597_/X _14605_/X VGND VGND VPWR VPWR _14606_/X
+ sky130_fd_sc_hd__a32o_4
X_15586_ _15586_/A _23339_/Q VGND VGND VPWR VPWR _15588_/B sky130_fd_sc_hd__or2_4
X_18374_ _17513_/A _18373_/B _17634_/X VGND VGND VPWR VPWR _18374_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12798_ _12771_/X _12798_/B _12797_/X VGND VGND VPWR VPWR _12806_/B sky130_fd_sc_hd__or3_4
XANTENNA__22437__A _20747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _13699_/A _14537_/B _14536_/X VGND VGND VPWR VPWR _14537_/X sky130_fd_sc_hd__and3_4
X_17325_ _15251_/X _17150_/A VGND VGND VPWR VPWR _17325_/X sky130_fd_sc_hd__or2_4
X_11749_ _11803_/A _11749_/B VGND VGND VPWR VPWR _11749_/X sky130_fd_sc_hd__or2_4
XFILLER_105_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12963__A _12963_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20883__A1 _20403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14468_ _12460_/A _14464_/X _14467_/X VGND VGND VPWR VPWR _14468_/X sky130_fd_sc_hd__or3_4
X_17256_ _17256_/A _17249_/A VGND VGND VPWR VPWR _17256_/X sky130_fd_sc_hd__or2_4
X_13419_ _13376_/X _13336_/B VGND VGND VPWR VPWR _13419_/X sky130_fd_sc_hd__or2_4
X_16207_ _16229_/A _16203_/X _16207_/C VGND VGND VPWR VPWR _16215_/B sky130_fd_sc_hd__or3_4
XANTENNA__22085__B1 _16408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17187_ _15782_/B _17155_/X _13591_/X _17186_/X VGND VGND VPWR VPWR _17187_/X sky130_fd_sc_hd__o22a_4
X_14399_ _15615_/A _14309_/B VGND VGND VPWR VPWR _14400_/C sky130_fd_sc_hd__or2_4
XANTENNA__22624__A2 _22622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18650__A _18381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20635__A1 _24206_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16138_ _16107_/A _23479_/Q VGND VGND VPWR VPWR _16140_/B sky130_fd_sc_hd__or2_4
XFILLER_6_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22172__A _22172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13794__A _13794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16069_ _16069_/A _24088_/Q VGND VGND VPWR VPWR _16070_/C sky130_fd_sc_hd__or2_4
XFILLER_83_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22900__A _22968_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19828_ _19429_/A _19689_/Y _19872_/B _19827_/X VGND VGND VPWR VPWR _19828_/X sky130_fd_sc_hd__a211o_4
XFILLER_97_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19481__A _19481_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19759_ _19612_/A _19759_/B _19758_/X VGND VGND VPWR VPWR _19759_/X sky130_fd_sc_hd__or3_4
XANTENNA__17713__B _17385_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15514__A _12613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21899__B1 _23563_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22770_ _22741_/Y _22768_/A VGND VGND VPWR VPWR _22770_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__21363__A2 _21362_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22560__B2 _22554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21721_ _21558_/X _21719_/X _13627_/B _21716_/X VGND VGND VPWR VPWR _21721_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15233__B _15176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24440_ _24277_/CLK _24440_/D HRESETn VGND VGND VPWR VPWR _24440_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13034__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21652_ _21659_/A VGND VGND VPWR VPWR _21652_/X sky130_fd_sc_hd__buf_2
XFILLER_36_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_10_0_HCLK_A clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22347__A _22354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20603_ _20603_/A _20603_/B VGND VGND VPWR VPWR _20603_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21251__A _20574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24371_ _23358_/CLK _24371_/D HRESETn VGND VGND VPWR VPWR _24371_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__13969__A _13643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21583_ _21583_/A VGND VGND VPWR VPWR _21684_/C sky130_fd_sc_hd__buf_2
XANTENNA__12873__A _13032_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16345__A _16447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23322_ _24047_/CLK _23322_/D VGND VGND VPWR VPWR _22304_/A sky130_fd_sc_hd__dfxtp_4
X_20534_ _20534_/A _20533_/X VGND VGND VPWR VPWR _20534_/X sky130_fd_sc_hd__or2_4
XFILLER_14_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16064__B _23704_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23253_ _23827_/CLK _23253_/D VGND VGND VPWR VPWR _12564_/B sky130_fd_sc_hd__dfxtp_4
X_20465_ _20396_/X _20464_/X _12316_/B _20374_/X VGND VGND VPWR VPWR _20465_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22204_ _22219_/A VGND VGND VPWR VPWR _22212_/A sky130_fd_sc_hd__buf_2
XANTENNA__16999__B _16977_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20626__A1 _20448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20626__B2 _20625_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23184_ _23920_/CLK _22541_/X VGND VGND VPWR VPWR _13291_/B sky130_fd_sc_hd__dfxtp_4
X_20396_ _20511_/A VGND VGND VPWR VPWR _20396_/X sky130_fd_sc_hd__buf_2
XANTENNA__19806__D _19805_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22135_ _22134_/X _22125_/X _14520_/B _22132_/X VGND VGND VPWR VPWR _23429_/D sky130_fd_sc_hd__o22a_4
XFILLER_106_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22379__B2 _22344_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22066_ _11781_/B VGND VGND VPWR VPWR _22066_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21017_ _20315_/X _21016_/X _24061_/Q _21013_/X VGND VGND VPWR VPWR _24061_/D sky130_fd_sc_hd__o22a_4
XFILLER_48_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17904__A _18390_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12113__A _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21426__A _21419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15424__A _15424_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22000__B1 _23499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13770_ _13770_/A _13762_/X _13769_/X VGND VGND VPWR VPWR _13771_/C sky130_fd_sc_hd__and3_4
X_22968_ _22968_/A _18341_/Y _18384_/X VGND VGND VPWR VPWR _22968_/X sky130_fd_sc_hd__or3_4
XFILLER_74_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12721_ _15689_/A _23604_/Q VGND VGND VPWR VPWR _12721_/X sky130_fd_sc_hd__or2_4
XFILLER_83_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22551__B2 _22547_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21919_ _21919_/A VGND VGND VPWR VPWR _21935_/A sky130_fd_sc_hd__inv_2
XFILLER_71_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15143__B _15213_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22899_ _23015_/A VGND VGND VPWR VPWR _22899_/X sky130_fd_sc_hd__buf_2
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20984__B HRDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15440_ _13636_/A _15512_/B VGND VGND VPWR VPWR _15440_/X sky130_fd_sc_hd__or2_4
XFILLER_70_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12652_ _12652_/A VGND VGND VPWR VPWR _12953_/A sky130_fd_sc_hd__buf_2
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24202__CLK _24202_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22257__A _22286_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21106__A2 _21103_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _11974_/A VGND VGND VPWR VPWR _15047_/A sky130_fd_sc_hd__buf_2
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _14810_/A _15297_/B VGND VGND VPWR VPWR _15372_/C sky130_fd_sc_hd__or2_4
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13879__A _13879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12583_ _12583_/A VGND VGND VPWR VPWR _12605_/A sky130_fd_sc_hd__buf_2
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16255__A _15980_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12783__A _15725_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14322_ _14322_/A VGND VGND VPWR VPWR _15571_/A sky130_fd_sc_hd__buf_2
X_17110_ _21296_/A VGND VGND VPWR VPWR _19830_/A sky130_fd_sc_hd__inv_2
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ _20901_/A IRQ[4] VGND VGND VPWR VPWR _11534_/X sky130_fd_sc_hd__and2_4
X_18090_ _17659_/X _18089_/X _17659_/X _18089_/X VGND VGND VPWR VPWR _18090_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17041_ _17040_/X VGND VGND VPWR VPWR _17042_/A sky130_fd_sc_hd__buf_2
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ _14206_/A _14251_/X _14253_/C VGND VGND VPWR VPWR _14253_/X sky130_fd_sc_hd__and3_4
XANTENNA__22606__A2 _22600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19566__A _19517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18470__A _17874_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13204_ _12794_/A _13138_/B VGND VGND VPWR VPWR _13205_/C sky130_fd_sc_hd__or2_4
XFILLER_99_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14184_ _13709_/A VGND VGND VPWR VPWR _14206_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13135_ _12989_/A _13135_/B _13134_/X VGND VGND VPWR VPWR _13135_/X sky130_fd_sc_hd__and3_4
XANTENNA__17086__A _18048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21290__B2 _21230_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18992_ _18965_/X _18990_/Y _18991_/Y _18968_/X VGND VGND VPWR VPWR _18992_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20224__B _20224_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13066_ _13112_/A _23506_/Q VGND VGND VPWR VPWR _13067_/C sky130_fd_sc_hd__or2_4
X_17943_ _17282_/A _17942_/B _17878_/X VGND VGND VPWR VPWR _17943_/X sky130_fd_sc_hd__o21a_4
XFILLER_117_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22720__A _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12017_ _11999_/A _12017_/B _12017_/C VGND VGND VPWR VPWR _12017_/X sky130_fd_sc_hd__or3_4
XANTENNA__21042__B2 _21041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17874_ _17874_/A VGND VGND VPWR VPWR _17874_/X sky130_fd_sc_hd__buf_2
XFILLER_113_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19613_ _19549_/X _19589_/X _19612_/X _17533_/A _19585_/X VGND VGND VPWR VPWR _19613_/X
+ sky130_fd_sc_hd__a32o_4
X_16825_ _13583_/Y _16824_/X VGND VGND VPWR VPWR _16899_/B sky130_fd_sc_hd__and2_4
XFILLER_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12958__A _12958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11862__A _11861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19544_ HRDATA[29] VGND VGND VPWR VPWR _20317_/B sky130_fd_sc_hd__buf_2
X_16756_ _11823_/A _16754_/X _16755_/X VGND VGND VPWR VPWR _16756_/X sky130_fd_sc_hd__and3_4
XFILLER_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13968_ _13968_/A _13966_/X _13968_/C VGND VGND VPWR VPWR _13968_/X sky130_fd_sc_hd__and3_4
XFILLER_34_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21345__A2 _21340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22542__B2 _22540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16149__B _16219_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15707_ _15707_/A _15766_/B VGND VGND VPWR VPWR _15708_/C sky130_fd_sc_hd__or2_4
XANTENNA__15053__B _23487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12919_ _13016_/A _23859_/Q VGND VGND VPWR VPWR _12920_/C sky130_fd_sc_hd__or2_4
X_19475_ _24156_/Q _19435_/A HRDATA[30] _19431_/X VGND VGND VPWR VPWR _19475_/X sky130_fd_sc_hd__o22a_4
XFILLER_59_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13899_ _13700_/A _13899_/B _13899_/C VGND VGND VPWR VPWR _13900_/C sky130_fd_sc_hd__and3_4
X_16687_ _16714_/A _23739_/Q VGND VGND VPWR VPWR _16688_/C sky130_fd_sc_hd__or2_4
X_18426_ _18424_/X _18326_/Y _18249_/X _18425_/X VGND VGND VPWR VPWR _18426_/X sky130_fd_sc_hd__a211o_4
XFILLER_61_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15638_ _15626_/A _15636_/X _15637_/X VGND VGND VPWR VPWR _15642_/B sky130_fd_sc_hd__and3_4
XFILLER_72_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14892__B _14892_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13789__A _15404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18357_ _18202_/A VGND VGND VPWR VPWR _18357_/X sky130_fd_sc_hd__buf_2
X_15569_ _12441_/A _23211_/Q VGND VGND VPWR VPWR _15571_/B sky130_fd_sc_hd__or2_4
XANTENNA__12693__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17308_ _17143_/X _17860_/A VGND VGND VPWR VPWR _17308_/X sky130_fd_sc_hd__or2_4
XFILLER_33_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18288_ _17677_/X _18287_/X _17677_/X _18287_/X VGND VGND VPWR VPWR _18288_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17239_ _18750_/A _17084_/A VGND VGND VPWR VPWR _18249_/A sky130_fd_sc_hd__nand2_4
XFILLER_50_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18811__C _12036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20250_ _20468_/A VGND VGND VPWR VPWR _20622_/A sky130_fd_sc_hd__buf_2
XANTENNA__17708__B _17413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20181_ _18724_/X _20057_/X _20180_/Y _19929_/X VGND VGND VPWR VPWR _20181_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15509__A _15497_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21281__B2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_12_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR _23812_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__19816__A2_N _19815_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_75_0_HCLK clkbuf_7_75_0_HCLK/A VGND VGND VPWR VPWR _23867_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23940_ _23363_/CLK _23940_/D VGND VGND VPWR VPWR _14689_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_9_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13029__A _13029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21033__B2 _21027_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23871_ _23487_/CLK _21346_/X VGND VGND VPWR VPWR _23871_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12868__A _12868_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11772__A _16215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22822_ _15713_/Y _22814_/X _22795_/X _22821_/X VGND VGND VPWR VPWR _22823_/B sky130_fd_sc_hd__o22a_4
XANTENNA__15244__A _14210_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18737__B1 _17090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21336__A2 _21333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_3_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22753_ _24095_/D VGND VGND VPWR VPWR _22768_/C sky130_fd_sc_hd__inv_2
XFILLER_92_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21704_ _21529_/X _21698_/X _12799_/B _21702_/X VGND VGND VPWR VPWR _21704_/X sky130_fd_sc_hd__o22a_4
X_22684_ _20487_/A _22679_/X _12657_/B _22683_/X VGND VGND VPWR VPWR _23093_/D sky130_fd_sc_hd__o22a_4
XFILLER_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15898__B _15828_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22077__A _22101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24423_ _24425_/CLK _18800_/X HRESETn VGND VGND VPWR VPWR _24423_/Q sky130_fd_sc_hd__dfrtp_4
X_21635_ _21634_/X VGND VGND VPWR VPWR _21636_/A sky130_fd_sc_hd__buf_2
XANTENNA__13699__A _13699_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16075__A _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24354_ _24321_/CLK _24354_/D HRESETn VGND VGND VPWR VPWR _19094_/A sky130_fd_sc_hd__dfstp_4
XFILLER_103_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21566_ _21565_/X _21556_/X _14506_/B _21563_/X VGND VGND VPWR VPWR _21566_/X sky130_fd_sc_hd__o22a_4
X_23305_ _23433_/CLK _23305_/D VGND VGND VPWR VPWR _14217_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20517_ _20517_/A VGND VGND VPWR VPWR _20517_/X sky130_fd_sc_hd__buf_2
X_24285_ _24435_/CLK _24285_/D HRESETn VGND VGND VPWR VPWR _24285_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21497_ _21293_/X _21470_/A _23775_/Q _21452_/X VGND VGND VPWR VPWR _23775_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12108__A _16541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23236_ _24065_/CLK _23236_/D VGND VGND VPWR VPWR _14569_/B sky130_fd_sc_hd__dfxtp_4
X_20448_ _20255_/A VGND VGND VPWR VPWR _20448_/X sky130_fd_sc_hd__buf_2
XFILLER_88_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20325__A _20301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15419__A _13647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23167_ _23889_/CLK _22563_/X VGND VGND VPWR VPWR _23167_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21272__B2 _21266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20379_ _20379_/A VGND VGND VPWR VPWR _20380_/A sky130_fd_sc_hd__inv_2
XFILLER_69_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22118_ _22117_/X _22113_/X _15474_/B _22108_/X VGND VGND VPWR VPWR _22118_/X sky130_fd_sc_hd__o22a_4
X_23098_ _23706_/CLK _23098_/D VGND VGND VPWR VPWR _16434_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_7_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22540__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17228__B1 _17143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21024__B2 _21020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14940_ _15072_/A _14882_/B VGND VGND VPWR VPWR _14943_/B sky130_fd_sc_hd__or2_4
X_22049_ _22035_/A VGND VGND VPWR VPWR _22049_/X sky130_fd_sc_hd__buf_2
XFILLER_88_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21575__A2 _21568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14977__B _23456_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13881__B _13794_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14871_ _14912_/A VGND VGND VPWR VPWR _14895_/A sky130_fd_sc_hd__buf_2
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12778__A _12777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16610_ _16610_/A _23740_/Q VGND VGND VPWR VPWR _16611_/C sky130_fd_sc_hd__or2_4
X_13822_ _12211_/A _24071_/Q VGND VGND VPWR VPWR _13823_/C sky130_fd_sc_hd__or2_4
X_17590_ _17590_/A _17589_/X VGND VGND VPWR VPWR _17626_/C sky130_fd_sc_hd__or2_4
XANTENNA__21327__A2 _21326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22524__B2 _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13753_ _12638_/A _13753_/B _13753_/C VGND VGND VPWR VPWR _13754_/C sky130_fd_sc_hd__and3_4
X_16541_ _16541_/A _16541_/B _16540_/X VGND VGND VPWR VPWR _16542_/C sky130_fd_sc_hd__and3_4
XFILLER_16_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14993__A _14997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18465__A _18295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12704_ _15693_/A _12803_/B VGND VGND VPWR VPWR _12704_/X sky130_fd_sc_hd__or2_4
X_19260_ _19223_/A _19261_/A _19259_/Y VGND VGND VPWR VPWR _24274_/D sky130_fd_sc_hd__o21a_4
X_13684_ _13594_/X _13595_/X _13649_/X _11595_/A _13683_/X VGND VGND VPWR VPWR _13684_/X
+ sky130_fd_sc_hd__a32o_4
X_16472_ _16471_/X _16472_/B VGND VGND VPWR VPWR _16475_/B sky130_fd_sc_hd__or2_4
XFILLER_108_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18211_ _17861_/A _18210_/X _17836_/A _18041_/X VGND VGND VPWR VPWR _18212_/A sky130_fd_sc_hd__o22a_4
X_12635_ _12955_/A _12629_/X _12634_/X VGND VGND VPWR VPWR _12635_/X sky130_fd_sc_hd__or3_4
X_15423_ _12475_/A _15487_/B VGND VGND VPWR VPWR _15423_/X sky130_fd_sc_hd__or2_4
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19191_ _19113_/X VGND VGND VPWR VPWR _19191_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15601__B _23147_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15354_ _14008_/A _15354_/B _15354_/C VGND VGND VPWR VPWR _15362_/B sky130_fd_sc_hd__or3_4
X_18142_ _18142_/A VGND VGND VPWR VPWR _18392_/A sky130_fd_sc_hd__buf_2
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ _14002_/A VGND VGND VPWR VPWR _12567_/A sky130_fd_sc_hd__buf_2
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17703__B2 _17346_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22715__A _19770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11517_ _24332_/Q _11517_/B VGND VGND VPWR VPWR _11518_/B sky130_fd_sc_hd__or2_4
X_14305_ _15533_/A _14305_/B VGND VGND VPWR VPWR _14305_/X sky130_fd_sc_hd__or2_4
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15285_ _14149_/A _15285_/B VGND VGND VPWR VPWR _15285_/X sky130_fd_sc_hd__or2_4
X_18073_ _17845_/X _17253_/X _17797_/X _18072_/X VGND VGND VPWR VPWR _18073_/X sky130_fd_sc_hd__o22a_4
X_12497_ _13015_/A VGND VGND VPWR VPWR _12497_/X sky130_fd_sc_hd__buf_2
XANTENNA__12018__A _12022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14236_ _15190_/A _23817_/Q VGND VGND VPWR VPWR _14236_/X sky130_fd_sc_hd__or2_4
X_17024_ _17024_/A _17024_/B _17024_/C _17079_/A VGND VGND VPWR VPWR _17025_/A sky130_fd_sc_hd__or4_4
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14167_ _15045_/A VGND VGND VPWR VPWR _14617_/A sky130_fd_sc_hd__buf_2
X_13118_ _13118_/A _13110_/X _13117_/X VGND VGND VPWR VPWR _13134_/B sky130_fd_sc_hd__and3_4
X_14098_ _14098_/A _14093_/X _14097_/X VGND VGND VPWR VPWR _14098_/X sky130_fd_sc_hd__and3_4
X_18975_ _18975_/A VGND VGND VPWR VPWR _18975_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13049_ _13022_/A _13119_/B VGND VGND VPWR VPWR _13051_/B sky130_fd_sc_hd__or2_4
X_17926_ _17824_/X VGND VGND VPWR VPWR _17926_/X sky130_fd_sc_hd__buf_2
XFILLER_117_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23122__CLK _23122_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21566__A2 _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17857_ _17242_/A VGND VGND VPWR VPWR _18189_/A sky130_fd_sc_hd__buf_2
XFILLER_38_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12688__A _12688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16442__A1 _11982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16808_ _16621_/A _16806_/X _16807_/X VGND VGND VPWR VPWR _16808_/X sky130_fd_sc_hd__and3_4
X_17788_ _18066_/A _17267_/X VGND VGND VPWR VPWR _17788_/X sky130_fd_sc_hd__and2_4
XFILLER_81_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21318__A2 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19527_ _19523_/A _19829_/A _19861_/A _19526_/X VGND VGND VPWR VPWR _19527_/X sky130_fd_sc_hd__a211o_4
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16739_ _11966_/X _16739_/B _16739_/C VGND VGND VPWR VPWR _16740_/C sky130_fd_sc_hd__and3_4
XFILLER_35_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15999__A _13448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19458_ _19458_/A VGND VGND VPWR VPWR _19458_/X sky130_fd_sc_hd__buf_2
XFILLER_74_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18409_ _17753_/C _17753_/B _17696_/B VGND VGND VPWR VPWR _18409_/X sky130_fd_sc_hd__o21a_4
X_19389_ _19385_/A VGND VGND VPWR VPWR _19389_/X sky130_fd_sc_hd__buf_2
X_21420_ _21246_/X _21419_/X _23827_/Q _21416_/X VGND VGND VPWR VPWR _23827_/D sky130_fd_sc_hd__o22a_4
XANTENNA__13312__A _15697_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20829__B2 _20686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21351_ _21373_/A VGND VGND VPWR VPWR _21359_/A sky130_fd_sc_hd__buf_2
XANTENNA__16623__A _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20302_ _20622_/A _20300_/Y _24285_/Q _20301_/X VGND VGND VPWR VPWR _20302_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24070_ _23845_/CLK _20840_/X VGND VGND VPWR VPWR _14320_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_50_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21282_ _21282_/A VGND VGND VPWR VPWR _21282_/X sky130_fd_sc_hd__buf_2
XFILLER_85_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23021_ _23003_/A _23021_/B VGND VGND VPWR VPWR _23023_/B sky130_fd_sc_hd__nand2_4
X_20233_ _20459_/A VGND VGND VPWR VPWR _20233_/X sky130_fd_sc_hd__buf_2
XANTENNA__19934__A _20000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14143__A _14143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20164_ _11566_/X _20163_/Y VGND VGND VPWR VPWR _20164_/X sky130_fd_sc_hd__or2_4
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20095_ _19411_/X _20094_/X _19377_/X _22907_/B VGND VGND VPWR VPWR _24114_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21557__A2 _21556_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23923_ _23859_/CLK _21248_/X VGND VGND VPWR VPWR _23923_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12598__A _12598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_5_0_HCLK clkbuf_6_2_0_HCLK/X VGND VGND VPWR VPWR _24229_/CLK sky130_fd_sc_hd__clkbuf_1
X_23854_ _23342_/CLK _21377_/X VGND VGND VPWR VPWR _15766_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22506__B2 _22504_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22805_ _17411_/Y _22794_/X _22796_/X _22804_/X VGND VGND VPWR VPWR _22806_/B sky130_fd_sc_hd__o22a_4
X_23785_ _23561_/CLK _21485_/X VGND VGND VPWR VPWR _23785_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20997_ _20997_/A VGND VGND VPWR VPWR _20997_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11652__D _11652_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12110__B _23869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19383__B1 _19380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22736_ SYSTICKCLKDIV[1] VGND VGND VPWR VPWR _22736_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15702__A _15820_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22667_ _22671_/A VGND VGND VPWR VPWR _22683_/A sky130_fd_sc_hd__inv_2
XFILLER_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14318__A _14318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12420_ _12388_/A _12420_/B _12420_/C VGND VGND VPWR VPWR _12420_/X sky130_fd_sc_hd__and3_4
X_24406_ _24277_/CLK _18832_/X HRESETn VGND VGND VPWR VPWR _24406_/Q sky130_fd_sc_hd__dfrtp_4
X_21618_ _21553_/X _21612_/X _23722_/Q _21616_/X VGND VGND VPWR VPWR _23722_/D sky130_fd_sc_hd__o22a_4
X_22598_ _22434_/X _22593_/X _23147_/Q _22597_/X VGND VGND VPWR VPWR _22598_/X sky130_fd_sc_hd__o22a_4
X_12351_ _12360_/A _12222_/B VGND VGND VPWR VPWR _12351_/X sky130_fd_sc_hd__or2_4
X_24337_ _23358_/CLK _19012_/X HRESETn VGND VGND VPWR VPWR _24337_/Q sky130_fd_sc_hd__dfstp_4
X_21549_ _21548_/X _21544_/X _15463_/B _21539_/X VGND VGND VPWR VPWR _23756_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21493__B2 _21488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16533__A _12112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15070_ _12583_/A _23551_/Q VGND VGND VPWR VPWR _15071_/C sky130_fd_sc_hd__or2_4
XFILLER_68_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12282_ _13026_/A VGND VGND VPWR VPWR _12892_/A sky130_fd_sc_hd__buf_2
X_24268_ _24365_/CLK _24268_/D HRESETn VGND VGND VPWR VPWR _19217_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_119_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14021_ _14021_/A _23914_/Q VGND VGND VPWR VPWR _14023_/B sky130_fd_sc_hd__or2_4
X_23219_ _23155_/CLK _23219_/D VGND VGND VPWR VPWR _12983_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15149__A _14121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11677__A _13992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21245__B2 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19844__A _19844_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24199_ _24199_/CLK _19402_/X HRESETn VGND VGND VPWR VPWR _24199_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21796__A2 _21793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18760_ _17040_/A _17028_/A _18760_/C _17384_/Y VGND VGND VPWR VPWR _18812_/C sky130_fd_sc_hd__or4_4
XFILLER_7_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15972_ _11980_/X _15972_/B VGND VGND VPWR VPWR _15972_/X sky130_fd_sc_hd__and2_4
XFILLER_103_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22745__A1 SYSTICKCLKDIV[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17711_ _16970_/A _17393_/X VGND VGND VPWR VPWR _17748_/A sky130_fd_sc_hd__or2_4
X_14923_ _12340_/A _14859_/B VGND VGND VPWR VPWR _14923_/X sky130_fd_sc_hd__or2_4
X_18691_ _17989_/X _17614_/X _17874_/X _17332_/X VGND VGND VPWR VPWR _18693_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__20220__A2 HRDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17642_ _16989_/A VGND VGND VPWR VPWR _17766_/A sky130_fd_sc_hd__buf_2
XFILLER_36_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14854_ _14786_/Y _14851_/X _15387_/B VGND VGND VPWR VPWR _14855_/A sky130_fd_sc_hd__o21a_4
XFILLER_75_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13805_ _15420_/A _13805_/B VGND VGND VPWR VPWR _13805_/X sky130_fd_sc_hd__and2_4
XFILLER_75_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17573_ _18085_/A _17571_/Y _17572_/X VGND VGND VPWR VPWR _17573_/X sky130_fd_sc_hd__o21a_4
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11997_ _11997_/A _24062_/Q VGND VGND VPWR VPWR _11998_/C sky130_fd_sc_hd__or2_4
X_14785_ _11841_/A _13595_/A _14754_/X _11594_/A _14784_/X VGND VGND VPWR VPWR _14785_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16708__A _11921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19312_ _19933_/A VGND VGND VPWR VPWR _19313_/A sky130_fd_sc_hd__buf_2
X_16524_ _16523_/X VGND VGND VPWR VPWR _16524_/Y sky130_fd_sc_hd__inv_2
X_13736_ _12652_/A _13636_/B VGND VGND VPWR VPWR _13737_/C sky130_fd_sc_hd__or2_4
XANTENNA__21181__B1 _12640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21720__A2 _21719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16427__B _16427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19243_ _19231_/X VGND VGND VPWR VPWR _19243_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16455_ _11702_/A _16387_/B VGND VGND VPWR VPWR _16457_/B sky130_fd_sc_hd__or2_4
X_13667_ _15412_/A _13663_/X _13667_/C VGND VGND VPWR VPWR _13667_/X sky130_fd_sc_hd__or3_4
XFILLER_32_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14228__A _14207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15406_ _13794_/A _15406_/B VGND VGND VPWR VPWR _15406_/X sky130_fd_sc_hd__or2_4
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12618_ _15491_/A VGND VGND VPWR VPWR _12947_/A sky130_fd_sc_hd__buf_2
X_19174_ _19122_/A _19122_/B _19173_/Y VGND VGND VPWR VPWR _19174_/X sky130_fd_sc_hd__o21a_4
XFILLER_73_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13598_ _13986_/A VGND VGND VPWR VPWR _14782_/A sky130_fd_sc_hd__buf_2
X_16386_ _15929_/X _16382_/X _16385_/X VGND VGND VPWR VPWR _16386_/X sky130_fd_sc_hd__or3_4
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18125_ _17950_/X _18098_/X _18022_/X _18124_/X VGND VGND VPWR VPWR _18125_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20287__A2 _20650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12549_ _12914_/A _12549_/B _12548_/X VGND VGND VPWR VPWR _12549_/X sky130_fd_sc_hd__or3_4
X_15337_ _12598_/A _15335_/X _15336_/X VGND VGND VPWR VPWR _15338_/C sky130_fd_sc_hd__and3_4
XFILLER_34_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17539__A _17144_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12971__A _12655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18056_ _18129_/A VGND VGND VPWR VPWR _18056_/X sky130_fd_sc_hd__buf_2
X_15268_ _14727_/A _15266_/X _15268_/C VGND VGND VPWR VPWR _15268_/X sky130_fd_sc_hd__and3_4
XFILLER_67_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17007_ _12186_/B VGND VGND VPWR VPWR _17007_/X sky130_fd_sc_hd__buf_2
X_14219_ _14218_/X _23529_/Q VGND VGND VPWR VPWR _14220_/C sky130_fd_sc_hd__or2_4
XANTENNA__21236__B2 _21230_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19754__A _19754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22433__B1 _15454_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15199_ _14201_/A _15199_/B _15198_/X VGND VGND VPWR VPWR _15199_/X sky130_fd_sc_hd__or3_4
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18958_ _11530_/A VGND VGND VPWR VPWR _18958_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17909_ _17800_/X _17906_/Y _17812_/X _17908_/Y VGND VGND VPWR VPWR _17909_/X sky130_fd_sc_hd__o22a_4
X_18889_ _12430_/X _18884_/X _24374_/Q _18885_/X VGND VGND VPWR VPWR _18889_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20920_ _20842_/X _20918_/X _20919_/X HRDATA[11] _20847_/X VGND VGND VPWR VPWR _20920_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13307__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12211__A _12211_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21524__A _20464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20851_ _20850_/Y VGND VGND VPWR VPWR _20851_/X sky130_fd_sc_hd__buf_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16618__A _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15522__A _12233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23570_ _23986_/CLK _21889_/X VGND VGND VPWR VPWR _13085_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20782_ _20400_/B _20822_/B VGND VGND VPWR VPWR _20783_/C sky130_fd_sc_hd__or2_4
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21711__A2 _21705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22521_ _22521_/A VGND VGND VPWR VPWR _22536_/A sky130_fd_sc_hd__buf_2
XANTENNA__18427__A1_N _17261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19929__A _19996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14138__A _14121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13042__A _13015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22452_ _22384_/X VGND VGND VPWR VPWR _22452_/X sky130_fd_sc_hd__buf_2
X_21403_ _21397_/Y _21402_/X _21219_/X _21402_/X VGND VGND VPWR VPWR _21403_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17449__A _16569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13977__A _12209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22383_ _22068_/A _21582_/A _22383_/C _21784_/D VGND VGND VPWR VPWR _22384_/A sky130_fd_sc_hd__or4_4
XANTENNA__21475__B2 _21474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16353__A _13415_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24122_ _24126_/CLK _20047_/Y HRESETn VGND VGND VPWR VPWR _24122_/Q sky130_fd_sc_hd__dfrtp_4
X_21334_ _21270_/X _21333_/X _23881_/Q _21330_/X VGND VGND VPWR VPWR _23881_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15154__A1 _11847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24053_ _24021_/CLK _24053_/D VGND VGND VPWR VPWR _12643_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22424__B1 _13282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24326__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21265_ _21265_/A VGND VGND VPWR VPWR _21265_/X sky130_fd_sc_hd__buf_2
XFILLER_85_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23004_ _18222_/X _23004_/B VGND VGND VPWR VPWR _23005_/C sky130_fd_sc_hd__or2_4
XANTENNA__21778__A2 _21776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20216_ _24158_/Q _20445_/B VGND VGND VPWR VPWR _20216_/X sky130_fd_sc_hd__or2_4
X_21196_ _20748_/X _21190_/X _23946_/Q _21194_/X VGND VGND VPWR VPWR _23946_/D sky130_fd_sc_hd__o22a_4
XFILLER_46_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20986__B1 HRDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16800__B _23867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20450__A2 _20405_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20147_ _11534_/X VGND VGND VPWR VPWR _20147_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14601__A _15006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_45_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20078_ _18604_/X _18600_/X _20077_/X VGND VGND VPWR VPWR _20078_/X sky130_fd_sc_hd__o21a_4
XFILLER_92_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11920_ _11993_/A _11732_/B VGND VGND VPWR VPWR _11923_/B sky130_fd_sc_hd__or2_4
X_23906_ _23812_/CLK _23906_/D VGND VGND VPWR VPWR _15273_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_111_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12121__A _11692_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22520__A2_N _22519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21950__A2 _21945_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11851_ _13491_/A VGND VGND VPWR VPWR _11851_/X sky130_fd_sc_hd__buf_2
XFILLER_73_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23837_ _23867_/CLK _21406_/X VGND VGND VPWR VPWR _23837_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16528__A _16536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15432__A _15432_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14570_ _14096_/X _14646_/B VGND VGND VPWR VPWR _14571_/C sky130_fd_sc_hd__or2_4
XFILLER_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11782_ _11782_/A _11779_/X _11782_/C VGND VGND VPWR VPWR _11782_/X sky130_fd_sc_hd__and3_4
X_23768_ _23316_/CLK _23768_/D VGND VGND VPWR VPWR _23768_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_HCLK clkbuf_4_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13521_ _13559_/A _13521_/B VGND VGND VPWR VPWR _13521_/X sky130_fd_sc_hd__or2_4
X_22719_ _22967_/A VGND VGND VPWR VPWR _22719_/X sky130_fd_sc_hd__buf_2
X_23699_ _23699_/CLK _23699_/D VGND VGND VPWR VPWR _12976_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14048__A _14813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18743__A _18728_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13452_ _11861_/X _13452_/B _13452_/C VGND VGND VPWR VPWR _13452_/X sky130_fd_sc_hd__or3_4
X_16240_ _16145_/A _16240_/B VGND VGND VPWR VPWR _16240_/X sky130_fd_sc_hd__or2_4
XANTENNA__22265__A _22272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14990__B _23487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ _12418_/A _12297_/B VGND VGND VPWR VPWR _12405_/B sky130_fd_sc_hd__or2_4
X_13383_ _13383_/A _23984_/Q VGND VGND VPWR VPWR _13384_/C sky130_fd_sc_hd__or2_4
X_16171_ _16202_/A _16171_/B VGND VGND VPWR VPWR _16171_/X sky130_fd_sc_hd__or2_4
XANTENNA__17359__A _17191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21466__B2 _21460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24093__CLK _23485_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18331__A1 _18216_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12334_ _13055_/A _12334_/B _12333_/X VGND VGND VPWR VPWR _12334_/X sky130_fd_sc_hd__or3_4
X_15122_ _14918_/X _14988_/A _15120_/Y _15121_/X VGND VGND VPWR VPWR _15122_/X sky130_fd_sc_hd__o22a_4
X_15053_ _14068_/A _23487_/Q VGND VGND VPWR VPWR _15053_/X sky130_fd_sc_hd__or2_4
X_19930_ _19929_/X VGND VGND VPWR VPWR _19931_/B sky130_fd_sc_hd__inv_2
Xclkbuf_7_127_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR _23987_/CLK sky130_fd_sc_hd__clkbuf_1
X_12265_ _12706_/A _12249_/X _12264_/X VGND VGND VPWR VPWR _12265_/X sky130_fd_sc_hd__or3_4
XFILLER_99_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14004_ _14845_/A _23722_/Q VGND VGND VPWR VPWR _14005_/C sky130_fd_sc_hd__or2_4
XFILLER_29_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_6_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19861_ _19861_/A _19624_/A VGND VGND VPWR VPWR _19881_/A sky130_fd_sc_hd__or2_4
XANTENNA__21609__A _21602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12196_ _12196_/A VGND VGND VPWR VPWR _13677_/A sky130_fd_sc_hd__buf_2
XANTENNA__20513__A _18577_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18812_ _11599_/X _18866_/B _18812_/C _18812_/D VGND VGND VPWR VPWR _18813_/A sky130_fd_sc_hd__or4_4
XFILLER_68_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19792_ _19710_/X _19784_/X _19791_/X _16630_/X _19697_/X VGND VGND VPWR VPWR _19792_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18743_ _18728_/A _19941_/B VGND VGND VPWR VPWR _18743_/X sky130_fd_sc_hd__and2_4
X_15955_ _15984_/A _23672_/Q VGND VGND VPWR VPWR _15958_/B sky130_fd_sc_hd__or2_4
XANTENNA__22194__A2 _22193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19595__B1 HRDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14906_ _14906_/A _23616_/Q VGND VGND VPWR VPWR _14907_/C sky130_fd_sc_hd__or2_4
X_18674_ _17968_/X _17932_/Y _17933_/X _18673_/Y VGND VGND VPWR VPWR _18674_/X sky130_fd_sc_hd__a211o_4
XFILLER_48_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12031__A _11837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15886_ _15879_/A _15824_/B VGND VGND VPWR VPWR _15888_/B sky130_fd_sc_hd__or2_4
XFILLER_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21941__A2 _21938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17625_ _17590_/A _17591_/X _18274_/C VGND VGND VPWR VPWR _17626_/D sky130_fd_sc_hd__or3_4
XFILLER_97_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14837_ _14021_/A _14779_/B VGND VGND VPWR VPWR _14839_/B sky130_fd_sc_hd__or2_4
XFILLER_64_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12966__A _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11870__A _12465_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15342__A _14000_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17556_ _16077_/X _17572_/B VGND VGND VPWR VPWR _17556_/X sky130_fd_sc_hd__or2_4
X_14768_ _13600_/A _14764_/X _14767_/X VGND VGND VPWR VPWR _14768_/X sky130_fd_sc_hd__or3_4
X_16507_ _16158_/A _16430_/B VGND VGND VPWR VPWR _16507_/X sky130_fd_sc_hd__or2_4
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13719_ _15494_/A _23272_/Q VGND VGND VPWR VPWR _13719_/X sky130_fd_sc_hd__or2_4
XANTENNA__15061__B _23743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17487_ _17506_/A _17487_/B VGND VGND VPWR VPWR _17487_/X sky130_fd_sc_hd__or2_4
X_14699_ _14666_/X _14620_/B VGND VGND VPWR VPWR _14699_/X sky130_fd_sc_hd__or2_4
XANTENNA__18653__A _19994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19226_ _24277_/Q _19225_/X VGND VGND VPWR VPWR _19226_/X sky130_fd_sc_hd__and2_4
X_16438_ _16100_/X _16438_/B VGND VGND VPWR VPWR _16439_/C sky130_fd_sc_hd__or2_4
XFILLER_73_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13797__A _15435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21457__A1 _21221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19157_ _19157_/A VGND VGND VPWR VPWR _19157_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21457__B2 _21453_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16369_ _16447_/A _16369_/B _16369_/C VGND VGND VPWR VPWR _16370_/C sky130_fd_sc_hd__and3_4
XFILLER_30_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18108_ _17914_/X _17913_/Y _17800_/A _17908_/Y VGND VGND VPWR VPWR _18108_/X sky130_fd_sc_hd__o22a_4
X_19088_ _24323_/Q _11508_/B _11508_/X VGND VGND VPWR VPWR _19088_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__22903__A _18664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18039_ _18038_/X VGND VGND VPWR VPWR _18039_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21209__B2 _21165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12206__A _12553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21050_ _20870_/X _21044_/X _14536_/B _21048_/X VGND VGND VPWR VPWR _21050_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18086__B1 _17998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18625__A2 _18613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20001_ _24469_/Q VGND VGND VPWR VPWR _20001_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15517__A _11656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14421__A _15643_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22709__B2 _22704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22185__A2 _22179_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18828__A _18835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13037__A _12917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21952_ _21919_/A VGND VGND VPWR VPWR _21952_/X sky130_fd_sc_hd__buf_2
XFILLER_55_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20903_ _20425_/A _20900_/Y _20902_/X _19089_/Y _20709_/X VGND VGND VPWR VPWR _20903_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21254__A _21242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21883_ _21809_/X _21880_/X _12271_/B _21877_/X VGND VGND VPWR VPWR _23574_/D sky130_fd_sc_hd__o22a_4
XFILLER_58_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16348__A _16188_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12876__A _12876_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11780__A _11758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23622_ _23845_/CLK _21774_/X VGND VGND VPWR VPWR _14324_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15252__A _11879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20834_ _20673_/X _20824_/Y _20832_/X _20833_/Y _20692_/X VGND VGND VPWR VPWR _20834_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_70_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19889__A1 _19884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21145__B1 _23979_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12595__B _12463_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23553_ _23391_/CLK _21912_/X VGND VGND VPWR VPWR _23553_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20765_ _20764_/X VGND VGND VPWR VPWR _20765_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21696__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18561__A1 _17792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22504_ _22483_/A VGND VGND VPWR VPWR _22504_/X sky130_fd_sc_hd__buf_2
XANTENNA__18561__B2 _17338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23484_ _24026_/CLK _22026_/X VGND VGND VPWR VPWR _23484_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20696_ _20696_/A VGND VGND VPWR VPWR _21263_/A sky130_fd_sc_hd__buf_2
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22435_ _22423_/A VGND VGND VPWR VPWR _22435_/X sky130_fd_sc_hd__buf_2
XANTENNA__17179__A _17178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22645__B1 _15821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13500__A _12982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20317__B _20317_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22366_ _22119_/X _22361_/X _23275_/Q _22365_/X VGND VGND VPWR VPWR _23275_/D sky130_fd_sc_hd__o22a_4
XFILLER_100_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24105_ _24199_/CLK _22725_/X HRESETn VGND VGND VPWR VPWR _18652_/A sky130_fd_sc_hd__dfrtp_4
X_21317_ _21241_/X _21312_/X _12639_/B _21316_/X VGND VGND VPWR VPWR _23893_/D sky130_fd_sc_hd__o22a_4
X_22297_ _22143_/X _22293_/X _15128_/B _22262_/A VGND VGND VPWR VPWR _23329_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16811__A _16677_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23953__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12050_ _16689_/A _12050_/B _12050_/C VGND VGND VPWR VPWR _12050_/X sky130_fd_sc_hd__or3_4
X_24036_ _23363_/CLK _24036_/D VGND VGND VPWR VPWR _14692_/B sky130_fd_sc_hd__dfxtp_4
X_21248_ _21246_/X _21247_/X _23923_/Q _21242_/X VGND VGND VPWR VPWR _21248_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20423__A2 _20800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15427__A _15431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21179_ _20464_/X _21176_/X _12287_/B _21173_/X VGND VGND VPWR VPWR _21179_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21620__B2 _21616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15146__B _15146_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15740_ _12777_/X _15737_/X _15739_/X VGND VGND VPWR VPWR _15744_/B sky130_fd_sc_hd__and3_4
X_12952_ _12976_/A _22311_/A VGND VGND VPWR VPWR _12952_/X sky130_fd_sc_hd__or2_4
XFILLER_24_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11903_ _11903_/A _23518_/Q VGND VGND VPWR VPWR _11904_/C sky130_fd_sc_hd__or2_4
XFILLER_94_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21164__A _21168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15671_ _12705_/A _15669_/X _15670_/X VGND VGND VPWR VPWR _15671_/X sky130_fd_sc_hd__and3_4
X_12883_ _12883_/A VGND VGND VPWR VPWR _13608_/A sky130_fd_sc_hd__buf_2
X_17410_ _17621_/A VGND VGND VPWR VPWR _17422_/C sky130_fd_sc_hd__inv_2
XANTENNA__11690__A _16447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14622_ _13600_/A _14616_/X _14621_/X VGND VGND VPWR VPWR _14622_/X sky130_fd_sc_hd__or3_4
X_11834_ _11834_/A _11834_/B _11833_/X VGND VGND VPWR VPWR _11834_/X sky130_fd_sc_hd__or3_4
X_18390_ _18390_/A _18390_/B _18390_/C _18389_/X VGND VGND VPWR VPWR _18390_/X sky130_fd_sc_hd__or4_4
XFILLER_14_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21136__B1 _23985_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17042_/A VGND VGND VPWR VPWR _17363_/A sky130_fd_sc_hd__inv_2
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11765_ _14020_/A VGND VGND VPWR VPWR _11766_/A sky130_fd_sc_hd__buf_2
X_14553_ _13754_/A _14549_/X _14552_/X VGND VGND VPWR VPWR _14553_/X sky130_fd_sc_hd__or3_4
XFILLER_109_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11624__B1 NMI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17355__A2 _17340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _15892_/A _13504_/B VGND VGND VPWR VPWR _13505_/C sky130_fd_sc_hd__or2_4
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17272_ _16743_/X VGND VGND VPWR VPWR _17272_/Y sky130_fd_sc_hd__inv_2
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _14247_/A VGND VGND VPWR VPWR _11697_/A sky130_fd_sc_hd__buf_2
X_14484_ _13620_/A _14484_/B VGND VGND VPWR VPWR _14484_/X sky130_fd_sc_hd__or2_4
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20508__A _22413_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19011_ _18994_/X _19009_/X _19010_/Y _18999_/X VGND VGND VPWR VPWR _19011_/X sky130_fd_sc_hd__o22a_4
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16223_ _16223_/A _23479_/Q VGND VGND VPWR VPWR _16225_/B sky130_fd_sc_hd__or2_4
X_13435_ _13463_/A _13435_/B VGND VGND VPWR VPWR _13436_/C sky130_fd_sc_hd__or2_4
XFILLER_35_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21439__B2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13366_ _13357_/X _13364_/X _13366_/C VGND VGND VPWR VPWR _13370_/B sky130_fd_sc_hd__and3_4
X_16154_ _11982_/X _16130_/X _16137_/X _16144_/X _16153_/X VGND VGND VPWR VPWR _16154_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22723__A _22723_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15105_ _15105_/A _23679_/Q VGND VGND VPWR VPWR _15105_/X sky130_fd_sc_hd__or2_4
X_12317_ _12705_/A _12312_/X _12316_/X VGND VGND VPWR VPWR _12317_/X sky130_fd_sc_hd__and3_4
X_13297_ _13281_/X _13294_/X _13296_/X VGND VGND VPWR VPWR _13298_/C sky130_fd_sc_hd__and3_4
X_16085_ _16097_/A _23511_/Q VGND VGND VPWR VPWR _16086_/C sky130_fd_sc_hd__or2_4
XANTENNA__12026__A _16113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12248_ _12726_/A _12248_/B VGND VGND VPWR VPWR _12248_/X sky130_fd_sc_hd__or2_4
X_15036_ _15036_/A _23199_/Q VGND VGND VPWR VPWR _15038_/B sky130_fd_sc_hd__or2_4
X_19913_ _19909_/X _24150_/Q _19910_/X _20800_/A VGND VGND VPWR VPWR _24150_/D sky130_fd_sc_hd__o22a_4
XFILLER_9_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24372__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19844_ _19844_/A VGND VGND VPWR VPWR _19844_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15337__A _12598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12179_ _11820_/A _12177_/X _12179_/C VGND VGND VPWR VPWR _12179_/X sky130_fd_sc_hd__and3_4
XANTENNA__21611__B2 _21609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17291__A1 _14493_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19775_ _19607_/X VGND VGND VPWR VPWR _19775_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17291__B2 _17290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15056__B _15056_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16987_ _17646_/A _16986_/X VGND VGND VPWR VPWR _17894_/D sky130_fd_sc_hd__or2_4
XFILLER_111_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22167__A2 _22165_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19568__B1 HRDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18726_ _17962_/X _18365_/X _17964_/X VGND VGND VPWR VPWR _18726_/Y sky130_fd_sc_hd__o21ai_4
X_15938_ _15937_/X VGND VGND VPWR VPWR _15976_/A sky130_fd_sc_hd__buf_2
XFILLER_42_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21914__A2 _21887_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14895__B _14962_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18657_ _17090_/X _18655_/X _18656_/X VGND VGND VPWR VPWR _18657_/X sky130_fd_sc_hd__and3_4
XFILLER_77_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15869_ _13529_/X _15867_/X _15869_/C VGND VGND VPWR VPWR _15869_/X sky130_fd_sc_hd__and3_4
XFILLER_64_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12696__A _15688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16168__A _16198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18791__A1 _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17608_ _17608_/A _17295_/X _17607_/X VGND VGND VPWR VPWR _17619_/B sky130_fd_sc_hd__and3_4
XANTENNA__15072__A _15072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18588_ _18500_/X _18587_/X _17608_/A VGND VGND VPWR VPWR _18588_/X sky130_fd_sc_hd__o21a_4
XANTENNA_clkbuf_4_10_0_HCLK_A clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17539_ _17144_/Y _17570_/A VGND VGND VPWR VPWR _17957_/B sky130_fd_sc_hd__and2_4
XANTENNA__21802__A _21802_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21678__B2 _21673_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15800__A _15823_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20550_ _20588_/A _20550_/B VGND VGND VPWR VPWR _20550_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__20350__A1 _17944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_9_0_HCLK clkbuf_6_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__20418__A _20418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19209_ _19209_/A _19209_/B VGND VGND VPWR VPWR _19209_/X sky130_fd_sc_hd__and2_4
XANTENNA__22627__B1 _16489_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20481_ _20481_/A VGND VGND VPWR VPWR _20481_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22220_ _22095_/X _22215_/X _12651_/B _22219_/X VGND VGND VPWR VPWR _23381_/D sky130_fd_sc_hd__o22a_4
XFILLER_49_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22633__A _22633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22151_ _21784_/A _21917_/B _22383_/C _21866_/D VGND VGND VPWR VPWR _22151_/X sky130_fd_sc_hd__or4_4
XANTENNA__16631__A _16630_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21102_ _20870_/X _21096_/X _14442_/B _21100_/X VGND VGND VPWR VPWR _21102_/X sky130_fd_sc_hd__o22a_4
X_22082_ _22081_/X _22077_/X _16708_/B _22072_/X VGND VGND VPWR VPWR _23451_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21249__A _21249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_110_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR _24082_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_99_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16350__B _16282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21033_ _20574_/X _21030_/X _24049_/Q _21027_/X VGND VGND VPWR VPWR _24049_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19942__A _18265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14151__A _14151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13990__A _13989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22984_ _22984_/A VGND VGND VPWR VPWR HADDR[17] sky130_fd_sc_hd__inv_2
XFILLER_60_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21935_ _21935_/A VGND VGND VPWR VPWR _21935_/X sky130_fd_sc_hd__buf_2
XFILLER_76_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16078__A _16008_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21866_ _21684_/A _21784_/B _21784_/C _21866_/D VGND VGND VPWR VPWR _21866_/X sky130_fd_sc_hd__or4_4
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _24199_/Q _20751_/X _20816_/X VGND VGND VPWR VPWR _22129_/A sky130_fd_sc_hd__o21a_4
X_23605_ _23315_/CLK _23605_/D VGND VGND VPWR VPWR _12525_/B sky130_fd_sc_hd__dfxtp_4
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21712__A _21705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21797_ _21797_/A VGND VGND VPWR VPWR _21797_/X sky130_fd_sc_hd__buf_2
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _24428_/Q IRQ[13] _11549_/X VGND VGND VPWR VPWR _11550_/X sky130_fd_sc_hd__a21o_4
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20748_ _20748_/A VGND VGND VPWR VPWR _20748_/X sky130_fd_sc_hd__buf_2
X_23536_ _23635_/CLK _23536_/D VGND VGND VPWR VPWR _23536_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23467_ _23404_/CLK _22050_/X VGND VGND VPWR VPWR _23467_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20679_ _20619_/X _20678_/X _20617_/X VGND VGND VPWR VPWR _20679_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_109_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14326__A _12460_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _13228_/A _13162_/B VGND VGND VPWR VPWR _13222_/B sky130_fd_sc_hd__or2_4
XFILLER_7_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13230__A _13242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22418_ _20552_/A VGND VGND VPWR VPWR _22418_/X sky130_fd_sc_hd__buf_2
X_23398_ _23781_/CLK _22191_/X VGND VGND VPWR VPWR _23398_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22543__A _22536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13151_ _13317_/A _13146_/X _13150_/X VGND VGND VPWR VPWR _13151_/X sky130_fd_sc_hd__or3_4
X_22349_ _22091_/X _22347_/X _16103_/B _22344_/X VGND VGND VPWR VPWR _23287_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16541__A _16541_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12102_ _12101_/X _12177_/B VGND VGND VPWR VPWR _12102_/X sky130_fd_sc_hd__or2_4
X_13082_ _13082_/A _13082_/B _13082_/C VGND VGND VPWR VPWR _13083_/C sky130_fd_sc_hd__or3_4
XFILLER_65_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23043__B1 _22899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12033_ _18728_/A _12029_/X VGND VGND VPWR VPWR _12033_/X sky130_fd_sc_hd__and2_4
X_16910_ _16910_/A VGND VGND VPWR VPWR _16910_/X sky130_fd_sc_hd__buf_2
X_24019_ _23311_/CLK _21083_/X VGND VGND VPWR VPWR _24019_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19798__B1 _16907_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22397__A2 _22392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15157__A _11909_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17890_ _16988_/X VGND VGND VPWR VPWR _17891_/B sky130_fd_sc_hd__inv_2
X_16841_ _16841_/A _16840_/X VGND VGND VPWR VPWR _16841_/X sky130_fd_sc_hd__and2_4
XFILLER_24_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14996__A _14121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18468__A _18244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_15_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19560_ _19556_/Y _19766_/A VGND VGND VPWR VPWR _19579_/A sky130_fd_sc_hd__and2_4
XFILLER_65_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16772_ _16772_/A _23675_/Q VGND VGND VPWR VPWR _16774_/B sky130_fd_sc_hd__or2_4
XFILLER_59_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13984_ _13984_/A _23850_/Q VGND VGND VPWR VPWR _13985_/C sky130_fd_sc_hd__or2_4
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18511_ _18480_/X _18507_/X _18508_/X _18510_/X VGND VGND VPWR VPWR _18511_/X sky130_fd_sc_hd__o22a_4
X_15723_ _13100_/A _15721_/X _15722_/X VGND VGND VPWR VPWR _15727_/B sky130_fd_sc_hd__and3_4
X_12935_ _12935_/A VGND VGND VPWR VPWR _12949_/A sky130_fd_sc_hd__buf_2
X_19491_ _19449_/X _19454_/X _19489_/Y _18864_/C _19490_/X VGND VGND VPWR VPWR _19491_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_98_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17091__B _17090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18773__A1 _16514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18442_ _18442_/A _17360_/A VGND VGND VPWR VPWR _18442_/X sky130_fd_sc_hd__and2_4
XFILLER_18_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15654_ _15654_/A _15652_/X _15653_/X VGND VGND VPWR VPWR _15658_/B sky130_fd_sc_hd__and3_4
X_12866_ _12870_/A _12866_/B _12865_/X VGND VGND VPWR VPWR _12867_/C sky130_fd_sc_hd__and3_4
XFILLER_2_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20580__A1 _20448_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21109__B1 _23999_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22718__A _19108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14605_ _11976_/A _14605_/B VGND VGND VPWR VPWR _14605_/X sky130_fd_sc_hd__and2_4
X_11817_ _11772_/X _11817_/B _11816_/X VGND VGND VPWR VPWR _11836_/B sky130_fd_sc_hd__and3_4
X_18373_ _17513_/A _18373_/B VGND VGND VPWR VPWR _18373_/Y sky130_fd_sc_hd__nand2_4
X_15585_ _15623_/A _15585_/B _15585_/C VGND VGND VPWR VPWR _15589_/B sky130_fd_sc_hd__and3_4
X_12797_ _12813_/A _12793_/X _12796_/X VGND VGND VPWR VPWR _12797_/X sky130_fd_sc_hd__and3_4
XFILLER_37_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17322_/X _17323_/X VGND VGND VPWR VPWR _17324_/X sky130_fd_sc_hd__and2_4
X_14536_ _14536_/A _14536_/B VGND VGND VPWR VPWR _14536_/X sky130_fd_sc_hd__or2_4
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11729_/X VGND VGND VPWR VPWR _11748_/X sky130_fd_sc_hd__buf_2
XFILLER_30_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20238__A _20447_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17255_ _17837_/A _17253_/X _17254_/X VGND VGND VPWR VPWR _17255_/X sky130_fd_sc_hd__o21a_4
XFILLER_70_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14467_ _12862_/A _14467_/B _14467_/C VGND VGND VPWR VPWR _14467_/X sky130_fd_sc_hd__and3_4
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11679_ _13908_/A VGND VGND VPWR VPWR _12626_/A sky130_fd_sc_hd__buf_2
XANTENNA__14236__A _15190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16206_ _16206_/A _16206_/B _16206_/C VGND VGND VPWR VPWR _16207_/C sky130_fd_sc_hd__and3_4
XANTENNA__13140__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13418_ _13357_/X _13416_/X _13417_/X VGND VGND VPWR VPWR _13422_/B sky130_fd_sc_hd__and3_4
X_17186_ _17145_/A VGND VGND VPWR VPWR _17186_/X sky130_fd_sc_hd__buf_2
XANTENNA__23229__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14398_ _15586_/A _14308_/B VGND VGND VPWR VPWR _14400_/B sky130_fd_sc_hd__or2_4
X_16137_ _16113_/A _16137_/B _16137_/C VGND VGND VPWR VPWR _16137_/X sky130_fd_sc_hd__or3_4
XANTENNA__17547__A _16376_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20635__A2 _20614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13349_ _11842_/X _11618_/X _13316_/X _11596_/X _13348_/X VGND VGND VPWR VPWR _13349_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21832__B2 _21824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16068_ _16064_/A _23480_/Q VGND VGND VPWR VPWR _16070_/B sky130_fd_sc_hd__or2_4
XFILLER_103_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13794__B _13794_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16170__B _16096_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15019_ _15019_/A _23871_/Q VGND VGND VPWR VPWR _15021_/B sky130_fd_sc_hd__or2_4
XFILLER_102_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15067__A _15115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17264__A1 _16596_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19827_ _19670_/X _19817_/C _19827_/C VGND VGND VPWR VPWR _19827_/X sky130_fd_sc_hd__and3_4
XANTENNA__17264__B2 _17263_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19481__B _19481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19758_ _19754_/X _19757_/X _19481_/B _19683_/X VGND VGND VPWR VPWR _19758_/X sky130_fd_sc_hd__o22a_4
XFILLER_42_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18097__B _18174_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18709_ _18605_/X _18708_/X _24449_/Q _18604_/X VGND VGND VPWR VPWR _24449_/D sky130_fd_sc_hd__o22a_4
X_19689_ _19689_/A VGND VGND VPWR VPWR _19689_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21899__B2 _21898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17405__A1_N _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21720_ _21555_/X _21719_/X _23657_/Q _21716_/X VGND VGND VPWR VPWR _23657_/D sky130_fd_sc_hd__o22a_4
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13315__A _12716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22560__A2 _22557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21651_ _21524_/X _21648_/X _12331_/B _21645_/X VGND VGND VPWR VPWR _23702_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21532__A _21532_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_35_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR _23781_/CLK sky130_fd_sc_hd__clkbuf_1
X_20602_ _20517_/X _20601_/X _24303_/Q _20527_/X VGND VGND VPWR VPWR _20603_/B sky130_fd_sc_hd__o22a_4
XFILLER_90_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15530__A _12260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24370_ _23326_/CLK _18895_/X HRESETn VGND VGND VPWR VPWR _24370_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA_clkbuf_4_9_0_HCLK_A clkbuf_4_9_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19002__A _19002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21582_ _21582_/A VGND VGND VPWR VPWR _21634_/B sky130_fd_sc_hd__buf_2
Xclkbuf_7_98_0_HCLK clkbuf_6_49_0_HCLK/X VGND VGND VPWR VPWR _23217_/CLK sky130_fd_sc_hd__clkbuf_1
X_23321_ _24026_/CLK _22305_/X VGND VGND VPWR VPWR _16259_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20533_ _24243_/Q _20421_/X _20532_/X VGND VGND VPWR VPWR _20533_/X sky130_fd_sc_hd__o21a_4
XFILLER_36_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14146__A _14119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13050__A _12512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23252_ _24047_/CLK _22414_/X VGND VGND VPWR VPWR _12758_/B sky130_fd_sc_hd__dfxtp_4
X_20464_ _20464_/A VGND VGND VPWR VPWR _20464_/X sky130_fd_sc_hd__buf_2
XANTENNA__24154__CLK _24293_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22203_ _22207_/A VGND VGND VPWR VPWR _22219_/A sky130_fd_sc_hd__inv_2
XFILLER_106_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16999__C _16999_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23183_ _23827_/CLK _22542_/X VGND VGND VPWR VPWR _13434_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17457__A _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20395_ _20280_/X _20394_/X _16365_/B _20374_/X VGND VGND VPWR VPWR _24089_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16361__A _11727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_HCLK clkbuf_2_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_118_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22134_ _22134_/A VGND VGND VPWR VPWR _22134_/X sky130_fd_sc_hd__buf_2
XANTENNA__22379__A2 _22375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22065_ _21863_/X _22031_/A _15033_/B _22020_/X VGND VGND VPWR VPWR _23455_/D sky130_fd_sc_hd__o22a_4
XFILLER_0_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22810__B _14786_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21016_ _21030_/A VGND VGND VPWR VPWR _21016_/X sky130_fd_sc_hd__buf_2
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17192__A _17191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15705__A _12744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22000__B2 _21999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22967_ _22967_/A VGND VGND VPWR VPWR _22967_/X sky130_fd_sc_hd__buf_2
XFILLER_5_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19952__B1 _17998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22551__A2 _22550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18755__B2 _18754_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12720_ _12720_/A _12720_/B _12720_/C VGND VGND VPWR VPWR _12724_/B sky130_fd_sc_hd__and3_4
XANTENNA__13225__A _13257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21918_ _21917_/X VGND VGND VPWR VPWR _21919_/A sky130_fd_sc_hd__buf_2
XFILLER_16_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22898_ _22898_/A _22897_/X VGND VGND VPWR VPWR HADDR[3] sky130_fd_sc_hd__nor2_4
XFILLER_71_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12651_ _12976_/A _12651_/B VGND VGND VPWR VPWR _12654_/B sky130_fd_sc_hd__or2_4
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21849_ _21847_/X _21841_/X _14304_/B _21848_/X VGND VGND VPWR VPWR _21849_/X sky130_fd_sc_hd__o22a_4
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16536__A _16536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18507__B2 _18506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19704__B1 _19877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _11599_/X _18866_/B VGND VGND VPWR VPWR _11602_/X sky130_fd_sc_hd__or2_4
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15440__A _13636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _12582_/A VGND VGND VPWR VPWR _12583_/A sky130_fd_sc_hd__buf_2
X_15370_ _14010_/A _15296_/B VGND VGND VPWR VPWR _15372_/B sky130_fd_sc_hd__or2_4
XANTENNA__24175__D _24175_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ _11911_/A _14317_/X _14321_/C VGND VGND VPWR VPWR _14321_/X sky130_fd_sc_hd__and3_4
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _24348_/Q _11532_/X _24350_/Q _11533_/D VGND VGND VPWR VPWR _11533_/X sky130_fd_sc_hd__or4_4
X_23519_ _23487_/CLK _23519_/D VGND VGND VPWR VPWR _23519_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ _17040_/A _17105_/B VGND VGND VPWR VPWR _17040_/X sky130_fd_sc_hd__or2_4
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14252_ _14252_/A _24073_/Q VGND VGND VPWR VPWR _14253_/C sky130_fd_sc_hd__or2_4
XFILLER_109_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13203_ _12791_/A _13137_/B VGND VGND VPWR VPWR _13203_/X sky130_fd_sc_hd__or2_4
XANTENNA__13895__A _13895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14183_ _14183_/A _14183_/B _14183_/C VGND VGND VPWR VPWR _14190_/B sky130_fd_sc_hd__and3_4
XFILLER_99_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13134_ _12672_/A _13134_/B _13133_/X VGND VGND VPWR VPWR _13134_/X sky130_fd_sc_hd__or3_4
XANTENNA__21290__A2 _21283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18991_ _24372_/Q VGND VGND VPWR VPWR _18991_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18691__B1 _17874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13065_ _13065_/A VGND VGND VPWR VPWR _13112_/A sky130_fd_sc_hd__buf_2
X_17942_ _17282_/A _17942_/B VGND VGND VPWR VPWR _17942_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__19582__A _19582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12016_ _16541_/A _12016_/B _12016_/C VGND VGND VPWR VPWR _12017_/C sky130_fd_sc_hd__and3_4
XFILLER_117_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21042__A2 _21037_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17873_ _17101_/X VGND VGND VPWR VPWR _17874_/A sky130_fd_sc_hd__buf_2
XFILLER_39_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18198__A _18198_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16824_ _13590_/X _13593_/B _13280_/X _16824_/D VGND VGND VPWR VPWR _16824_/X sky130_fd_sc_hd__or4_4
X_19612_ _19612_/A _19592_/X _19606_/Y _19611_/X VGND VGND VPWR VPWR _19612_/X sky130_fd_sc_hd__or4_4
XFILLER_24_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19543_ _19829_/A _19542_/X VGND VGND VPWR VPWR _19543_/X sky130_fd_sc_hd__or2_4
X_16755_ _16618_/X _23771_/Q VGND VGND VPWR VPWR _16755_/X sky130_fd_sc_hd__or2_4
X_13967_ _12472_/X _23818_/Q VGND VGND VPWR VPWR _13968_/C sky130_fd_sc_hd__or2_4
XANTENNA__22542__A2 _22536_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15706_ _15706_/A _15765_/B VGND VGND VPWR VPWR _15708_/B sky130_fd_sc_hd__or2_4
XFILLER_59_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13135__A _12989_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12918_ _13015_/A _12976_/B VGND VGND VPWR VPWR _12920_/B sky130_fd_sc_hd__or2_4
X_19474_ _19458_/X _19473_/X HRDATA[13] _19462_/X VGND VGND VPWR VPWR _19598_/A sky130_fd_sc_hd__o22a_4
X_16686_ _16686_/A _16749_/B VGND VGND VPWR VPWR _16688_/B sky130_fd_sc_hd__or2_4
XFILLER_46_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13898_ _13910_/A _23399_/Q VGND VGND VPWR VPWR _13899_/C sky130_fd_sc_hd__or2_4
XFILLER_62_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18425_ _18425_/A _18425_/B VGND VGND VPWR VPWR _18425_/X sky130_fd_sc_hd__and2_4
XFILLER_62_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21352__A _21359_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15637_ _15637_/A _24075_/Q VGND VGND VPWR VPWR _15637_/X sky130_fd_sc_hd__or2_4
X_12849_ _12849_/A _12849_/B _12849_/C VGND VGND VPWR VPWR _12849_/X sky130_fd_sc_hd__and3_4
XANTENNA__16446__A _11715_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_2_0_HCLK_A clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18356_ _17893_/X _18354_/X _16951_/A _18355_/Y VGND VGND VPWR VPWR _18356_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15568_ _14464_/A _15566_/X _15567_/X VGND VGND VPWR VPWR _15568_/X sky130_fd_sc_hd__and3_4
XANTENNA__12693__B _24020_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17307_ _17306_/X VGND VGND VPWR VPWR _17307_/Y sky130_fd_sc_hd__inv_2
X_14519_ _13879_/A VGND VGND VPWR VPWR _14519_/X sky130_fd_sc_hd__buf_2
X_18287_ _17678_/X _18286_/X _17675_/B VGND VGND VPWR VPWR _18287_/X sky130_fd_sc_hd__o21a_4
X_15499_ _13738_/A _15499_/B _15499_/C VGND VGND VPWR VPWR _15500_/C sky130_fd_sc_hd__or3_4
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17238_ _17238_/A VGND VGND VPWR VPWR _18716_/B sky130_fd_sc_hd__inv_2
XANTENNA__22058__B2 _22056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22183__A _22169_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17169_ _17227_/A _17149_/X _17251_/A _17168_/Y VGND VGND VPWR VPWR _17169_/X sky130_fd_sc_hd__o22a_4
X_20180_ _20180_/A VGND VGND VPWR VPWR _20180_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21281__A2 _21271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22911__A _19201_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12214__A _15654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21569__B1 _14662_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21033__A2 _21030_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21527__A _21527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13029__B _23954_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22230__B2 _22226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15525__A _15552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23870_ _23320_/CLK _21353_/X VGND VGND VPWR VPWR _23870_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22821_ _22821_/A _17283_/Y VGND VGND VPWR VPWR _22821_/X sky130_fd_sc_hd__or2_4
XANTENNA__15244__B _23617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18737__A1 _18656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13045__A _12553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22752_ _22727_/A _24097_/Q VGND VGND VPWR VPWR _22755_/B sky130_fd_sc_hd__nand2_4
XFILLER_25_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20544__A1 _20494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22358__A _22351_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21703_ _21526_/X _21698_/X _12627_/B _21702_/X VGND VGND VPWR VPWR _21703_/X sky130_fd_sc_hd__o22a_4
X_22683_ _22683_/A VGND VGND VPWR VPWR _22683_/X sky130_fd_sc_hd__buf_2
XFILLER_55_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15260__A _14318_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21634_ _21784_/A _21634_/B _21684_/C _21634_/D VGND VGND VPWR VPWR _21634_/X sky130_fd_sc_hd__or4_4
X_24422_ _24425_/CLK _24422_/D HRESETn VGND VGND VPWR VPWR _24422_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18274__C _18274_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22297__B2 _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21565_ _20870_/A VGND VGND VPWR VPWR _21565_/X sky130_fd_sc_hd__buf_2
X_24353_ _24320_/CLK _24353_/D HRESETn VGND VGND VPWR VPWR _19098_/A sky130_fd_sc_hd__dfstp_4
XFILLER_103_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23544__CLK _23539_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20516_ _20516_/A VGND VGND VPWR VPWR _20516_/X sky130_fd_sc_hd__buf_2
X_23304_ _23304_/CLK _22322_/X VGND VGND VPWR VPWR _23304_/Q sky130_fd_sc_hd__dfxtp_4
X_24284_ _24435_/CLK _24284_/D HRESETn VGND VGND VPWR VPWR _24284_/Q sky130_fd_sc_hd__dfrtp_4
X_21496_ _21291_/X _21491_/X _23776_/Q _21452_/X VGND VGND VPWR VPWR _23776_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22093__A _20463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23235_ _23107_/CLK _23235_/D VGND VGND VPWR VPWR _14787_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20447_ _20447_/A VGND VGND VPWR VPWR _20447_/X sky130_fd_sc_hd__buf_2
XFILLER_118_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14604__A _14752_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23166_ _23358_/CLK _22570_/X VGND VGND VPWR VPWR _11779_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21272__A2 _21271_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20378_ _24409_/Q _20519_/B VGND VGND VPWR VPWR _20378_/Y sky130_fd_sc_hd__nand2_4
XFILLER_49_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22117_ _20696_/A VGND VGND VPWR VPWR _22117_/X sky130_fd_sc_hd__buf_2
XFILLER_79_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23097_ _23770_/CLK _22678_/X VGND VGND VPWR VPWR _16293_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_66_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12124__A _16072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17228__A1 _17144_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22048_ _21833_/X _22045_/X _23468_/Q _22042_/X VGND VGND VPWR VPWR _22048_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21437__A _21416_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22221__B2 _22219_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15435__A _15435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14870_ _13956_/A _14865_/X _14869_/X VGND VGND VPWR VPWR _14870_/X sky130_fd_sc_hd__or3_4
XFILLER_48_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21980__B1 _23513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13821_ _15432_/A _23463_/Q VGND VGND VPWR VPWR _13821_/X sky130_fd_sc_hd__or2_4
XFILLER_63_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23999_ _23130_/CLK _23999_/D VGND VGND VPWR VPWR _23999_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22524__A2 _22522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16540_ _16565_/A _16620_/B VGND VGND VPWR VPWR _16540_/X sky130_fd_sc_hd__or2_4
XFILLER_21_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13752_ _12937_/A _23400_/Q VGND VGND VPWR VPWR _13753_/C sky130_fd_sc_hd__or2_4
XFILLER_90_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14993__B _23711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24198__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12703_ _12735_/A _23316_/Q VGND VGND VPWR VPWR _12703_/X sky130_fd_sc_hd__or2_4
X_16471_ _13352_/X VGND VGND VPWR VPWR _16471_/X sky130_fd_sc_hd__buf_2
X_13683_ _11977_/X _13658_/X _13667_/X _13674_/X _13682_/X VGND VGND VPWR VPWR _13683_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12794__A _12794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18210_ _17864_/A _17833_/X _17975_/A _17844_/X VGND VGND VPWR VPWR _18210_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24127__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15422_ _13651_/A _23884_/Q VGND VGND VPWR VPWR _15424_/B sky130_fd_sc_hd__or2_4
XANTENNA__15170__A _14152_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12634_ _12954_/A _12632_/X _12634_/C VGND VGND VPWR VPWR _12634_/X sky130_fd_sc_hd__and3_4
X_19190_ _19114_/A _19113_/X _19189_/Y VGND VGND VPWR VPWR _24293_/D sky130_fd_sc_hd__o21a_4
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22288__B2 _22283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18141_ _17962_/X _18113_/X _17869_/X VGND VGND VPWR VPWR _18141_/Y sky130_fd_sc_hd__o21ai_4
X_15353_ _15325_/X _15351_/X _15353_/C VGND VGND VPWR VPWR _15354_/C sky130_fd_sc_hd__and3_4
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _11707_/A VGND VGND VPWR VPWR _14002_/A sky130_fd_sc_hd__buf_2
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_81_0_HCLK clkbuf_6_40_0_HCLK/X VGND VGND VPWR VPWR _24344_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18900__A1 _13575_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14304_ _14283_/A _14304_/B VGND VGND VPWR VPWR _14304_/X sky130_fd_sc_hd__or2_4
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22715__B _16996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11516_ _24331_/Q _11516_/B VGND VGND VPWR VPWR _11517_/B sky130_fd_sc_hd__or2_4
X_18072_ _17824_/X _17843_/Y _17921_/A _17849_/Y VGND VGND VPWR VPWR _18072_/X sky130_fd_sc_hd__o22a_4
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15284_ _15144_/A _15282_/X _15283_/X VGND VGND VPWR VPWR _15288_/B sky130_fd_sc_hd__and3_4
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12496_ _12496_/A VGND VGND VPWR VPWR _13015_/A sky130_fd_sc_hd__buf_2
XANTENNA__16911__B1 _16903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17023_ _17022_/X VGND VGND VPWR VPWR _17023_/X sky130_fd_sc_hd__buf_2
X_14235_ _11708_/A VGND VGND VPWR VPWR _15190_/A sky130_fd_sc_hd__buf_2
XANTENNA__14514__A _11670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14166_ _11608_/A _14166_/B _14165_/X VGND VGND VPWR VPWR _14171_/B sky130_fd_sc_hd__and3_4
XFILLER_67_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13117_ _13101_/A _13113_/X _13117_/C VGND VGND VPWR VPWR _13117_/X sky130_fd_sc_hd__or3_4
X_14097_ _14096_/X _23273_/Q VGND VGND VPWR VPWR _14097_/X sky130_fd_sc_hd__or2_4
X_18974_ _18972_/Y _18973_/Y _11528_/X VGND VGND VPWR VPWR _18974_/X sky130_fd_sc_hd__o21a_4
XANTENNA__18416__B1 _18016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13048_ _13048_/A _13048_/B _13047_/X VGND VGND VPWR VPWR _13048_/X sky130_fd_sc_hd__or3_4
X_17925_ _17249_/X _17925_/B VGND VGND VPWR VPWR _17925_/X sky130_fd_sc_hd__and2_4
XANTENNA__12969__A _12981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11873__A _11872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15345__A _13992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17856_ _17933_/A VGND VGND VPWR VPWR _17856_/X sky130_fd_sc_hd__buf_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20774__A1 _20640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16807_ _16800_/A _23643_/Q VGND VGND VPWR VPWR _16807_/X sky130_fd_sc_hd__or2_4
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15064__B _23999_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17787_ _18443_/A VGND VGND VPWR VPWR _18066_/A sky130_fd_sc_hd__buf_2
XFILLER_82_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14999_ _15019_/A _23999_/Q VGND VGND VPWR VPWR _15001_/B sky130_fd_sc_hd__or2_4
XANTENNA__18719__A1 _18443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18656__A _18656_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17560__A _16155_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16738_ _11997_/A _23867_/Q VGND VGND VPWR VPWR _16739_/C sky130_fd_sc_hd__or2_4
X_19526_ _19672_/D _19526_/B _19525_/X VGND VGND VPWR VPWR _19526_/X sky130_fd_sc_hd__and3_4
XANTENNA__20526__A1 _20518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20526__B2 _20525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21082__A _21075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19457_ _19572_/B VGND VGND VPWR VPWR _19561_/A sky130_fd_sc_hd__buf_2
X_16669_ _16662_/A _23484_/Q VGND VGND VPWR VPWR _16671_/B sky130_fd_sc_hd__or2_4
X_18408_ _18314_/X _18385_/X _18357_/X _18407_/X VGND VGND VPWR VPWR _18408_/X sky130_fd_sc_hd__o22a_4
X_19388_ _19385_/X _18293_/X _19385_/X _24209_/Q VGND VGND VPWR VPWR _24209_/D sky130_fd_sc_hd__a2bb2o_4
X_18339_ _18291_/X _18338_/X _20025_/A _18291_/X VGND VGND VPWR VPWR _18339_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18391__A _18390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12209__A _12209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16904__A _16903_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21350_ _21383_/A VGND VGND VPWR VPWR _21373_/A sky130_fd_sc_hd__inv_2
XFILLER_30_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17719__B _17287_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20301_ _20301_/A VGND VGND VPWR VPWR _20301_/X sky130_fd_sc_hd__buf_2
X_21281_ _21280_/X _21271_/X _14453_/B _21278_/X VGND VGND VPWR VPWR _21281_/X sky130_fd_sc_hd__o22a_4
XANTENNA__14424__A _14423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23020_ _23020_/A VGND VGND VPWR VPWR HADDR[23] sky130_fd_sc_hd__inv_2
X_20232_ _20515_/A VGND VGND VPWR VPWR _20459_/A sky130_fd_sc_hd__buf_2
XFILLER_89_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20163_ _24440_/Q IRQ[25] _20162_/X VGND VGND VPWR VPWR _20163_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_118_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20094_ _20176_/A _20092_/X _20093_/Y _19936_/X VGND VGND VPWR VPWR _20094_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12879__A _12879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23922_ _23922_/CLK _21250_/X VGND VGND VPWR VPWR _23922_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15255__A _14315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23853_ _23922_/CLK _21378_/X VGND VGND VPWR VPWR _15839_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22506__A2 _22500_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22804_ _22807_/A _17115_/Y VGND VGND VPWR VPWR _22804_/X sky130_fd_sc_hd__or2_4
XFILLER_26_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20996_ _18752_/X _20332_/A _20640_/X _20995_/Y VGND VGND VPWR VPWR _20996_/X sky130_fd_sc_hd__a211o_4
X_23784_ _23304_/CLK _21486_/X VGND VGND VPWR VPWR _13757_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22088__A _20418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19383__A1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19383__B2 _24212_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22735_ SYSTICKCLKDIV[0] _22750_/A _22734_/X VGND VGND VPWR VPWR _22735_/X sky130_fd_sc_hd__a21bo_4
XFILLER_13_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24349__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16086__A _16109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13503__A _12959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22666_ _22665_/X VGND VGND VPWR VPWR _22671_/A sky130_fd_sc_hd__buf_2
XFILLER_71_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24405_ _24277_/CLK _24405_/D HRESETn VGND VGND VPWR VPWR _20469_/A sky130_fd_sc_hd__dfrtp_4
X_21617_ _21550_/X _21612_/X _23723_/Q _21616_/X VGND VGND VPWR VPWR _23723_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17146__B1 _17144_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22597_ _22583_/A VGND VGND VPWR VPWR _22597_/X sky130_fd_sc_hd__buf_2
XANTENNA__12119__A _16072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12350_ _12350_/A VGND VGND VPWR VPWR _12388_/A sky130_fd_sc_hd__buf_2
X_24336_ _23358_/CLK _19017_/X HRESETn VGND VGND VPWR VPWR _24336_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21493__A2 _21491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21548_ _21263_/A VGND VGND VPWR VPWR _21548_/X sky130_fd_sc_hd__buf_2
XFILLER_5_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12281_ _11596_/A VGND VGND VPWR VPWR _12281_/X sky130_fd_sc_hd__buf_2
XANTENNA__11958__A _12739_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21479_ _21261_/X _21477_/X _15836_/B _21474_/X VGND VGND VPWR VPWR _23789_/D sky130_fd_sc_hd__o22a_4
X_24267_ _23260_/CLK _19274_/X HRESETn VGND VGND VPWR VPWR _19216_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14334__A _13682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14020_ _14020_/A VGND VGND VPWR VPWR _14055_/A sky130_fd_sc_hd__buf_2
XFILLER_107_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23218_ _23155_/CLK _22488_/X VGND VGND VPWR VPWR _13045_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21245__A2 _21235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24198_ _24473_/CLK _19404_/X HRESETn VGND VGND VPWR VPWR _24198_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23149_ _23698_/CLK _22595_/X VGND VGND VPWR VPWR _15863_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_0_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15971_ _11933_/X _15966_/X _15971_/C VGND VGND VPWR VPWR _15972_/B sky130_fd_sc_hd__or3_4
XFILLER_62_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17710_ _18348_/A _17413_/X _17749_/B VGND VGND VPWR VPWR _17710_/X sky130_fd_sc_hd__a21o_4
X_14922_ _15063_/A _14922_/B _14922_/C VGND VGND VPWR VPWR _14926_/B sky130_fd_sc_hd__and3_4
X_18690_ _18604_/X _18688_/X _18689_/Y _11629_/X VGND VGND VPWR VPWR _24450_/D sky130_fd_sc_hd__a22oi_4
XFILLER_76_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17641_ _17769_/A _17263_/Y VGND VGND VPWR VPWR _17641_/X sky130_fd_sc_hd__and2_4
XFILLER_110_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14853_ _14785_/X _14852_/Y VGND VGND VPWR VPWR _15387_/B sky130_fd_sc_hd__or2_4
XFILLER_36_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ _13647_/A _13800_/X _13803_/X VGND VGND VPWR VPWR _13805_/B sky130_fd_sc_hd__or3_4
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17572_ _17165_/Y _17572_/B VGND VGND VPWR VPWR _17572_/X sky130_fd_sc_hd__or2_4
X_14784_ _15420_/A _14761_/X _14768_/X _14775_/X _14783_/X VGND VGND VPWR VPWR _14784_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11996_ _11996_/A _23614_/Q VGND VGND VPWR VPWR _11998_/B sky130_fd_sc_hd__or2_4
X_19311_ _22888_/A VGND VGND VPWR VPWR _19933_/A sky130_fd_sc_hd__buf_2
XFILLER_90_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16523_ _16378_/Y _16516_/X _16515_/X _16522_/Y VGND VGND VPWR VPWR _16523_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16708__B _16708_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13735_ _13735_/A _23304_/Q VGND VGND VPWR VPWR _13737_/B sky130_fd_sc_hd__or2_4
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21181__B2 _21180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19242_ _19232_/A _19231_/X _19241_/Y VGND VGND VPWR VPWR _24283_/D sky130_fd_sc_hd__o21a_4
XFILLER_31_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16454_ _16355_/X _16447_/X _16453_/X VGND VGND VPWR VPWR _16454_/X sky130_fd_sc_hd__or3_4
X_13666_ _15411_/A _13666_/B _13665_/X VGND VGND VPWR VPWR _13667_/C sky130_fd_sc_hd__and3_4
X_15405_ _13813_/A _15401_/X _15405_/C VGND VGND VPWR VPWR _15405_/X sky130_fd_sc_hd__or3_4
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12617_ _12617_/A VGND VGND VPWR VPWR _15491_/A sky130_fd_sc_hd__buf_2
X_19173_ _19123_/B VGND VGND VPWR VPWR _19173_/Y sky130_fd_sc_hd__inv_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16385_ _11915_/A _16383_/X _16384_/X VGND VGND VPWR VPWR _16385_/X sky130_fd_sc_hd__and3_4
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ _15450_/A VGND VGND VPWR VPWR _13597_/X sky130_fd_sc_hd__buf_2
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18124_ _18099_/X _18106_/Y _18120_/X _18122_/Y _18123_/X VGND VGND VPWR VPWR _18124_/X
+ sky130_fd_sc_hd__a32o_4
X_15336_ _12567_/A _15277_/B VGND VGND VPWR VPWR _15336_/X sky130_fd_sc_hd__or2_4
X_12548_ _12493_/A _12546_/X _12548_/C VGND VGND VPWR VPWR _12548_/X sky130_fd_sc_hd__and3_4
XFILLER_12_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22681__A1 _20442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22681__B2 _22676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18055_ _18009_/X _18051_/X _18053_/X _18054_/X VGND VGND VPWR VPWR _18055_/X sky130_fd_sc_hd__o22a_4
XFILLER_8_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11868__A _13654_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15267_ _11894_/A _15267_/B VGND VGND VPWR VPWR _15268_/C sky130_fd_sc_hd__or2_4
X_12479_ _12466_/X _12479_/B _12478_/X VGND VGND VPWR VPWR _12480_/C sky130_fd_sc_hd__and3_4
X_17006_ _17006_/A VGND VGND VPWR VPWR _17006_/X sky130_fd_sc_hd__buf_2
X_14218_ _14218_/A VGND VGND VPWR VPWR _14218_/X sky130_fd_sc_hd__buf_2
XANTENNA__21236__A2 _21235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15198_ _14215_/A _15196_/X _15197_/X VGND VGND VPWR VPWR _15198_/X sky130_fd_sc_hd__and3_4
XANTENNA__22433__B2 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14149_ _14149_/A _23465_/Q VGND VGND VPWR VPWR _14149_/X sky130_fd_sc_hd__or2_4
XANTENNA__17555__A _17164_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14898__B _14898_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18957_ _18937_/X _18955_/X _18956_/X _24346_/Q VGND VGND VPWR VPWR _18957_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12699__A _15689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17908_ _17908_/A VGND VGND VPWR VPWR _17908_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19770__A HRDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18888_ _16233_/X _18884_/X _18975_/A _18885_/X VGND VGND VPWR VPWR _18888_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21805__A _21817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17839_ _17814_/X _17206_/X _17804_/X _17202_/X VGND VGND VPWR VPWR _17839_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18386__A _18204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19310__A1_N _19303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20850_ _20641_/X _20849_/X _20754_/B VGND VGND VPWR VPWR _20850_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__15803__A _12522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19509_ _19422_/X _19508_/X HRDATA[8] _19438_/X VGND VGND VPWR VPWR _19729_/B sky130_fd_sc_hd__o22a_4
X_20781_ HRDATA[9] _20821_/B VGND VGND VPWR VPWR _20781_/X sky130_fd_sc_hd__or2_4
XANTENNA__15522__B _15522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17376__B1 _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21172__B2 _21166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22520_ _22514_/Y _22519_/X _22388_/X _22519_/X VGND VGND VPWR VPWR _22520_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22636__A _22636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13042__B _23474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22451_ _20892_/A VGND VGND VPWR VPWR _22451_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16634__A _16652_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22121__B1 _23435_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21402_ _21401_/X VGND VGND VPWR VPWR _21402_/X sky130_fd_sc_hd__buf_2
X_22382_ _11705_/B VGND VGND VPWR VPWR _22382_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21475__A2 _21470_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21333_ _21300_/A VGND VGND VPWR VPWR _21333_/X sky130_fd_sc_hd__buf_2
X_24121_ _24126_/CLK _20052_/Y HRESETn VGND VGND VPWR VPWR _24121_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11778__A _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14154__A _15015_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21264_ _21263_/X _21259_/X _23916_/Q _21254_/X VGND VGND VPWR VPWR _23916_/D sky130_fd_sc_hd__o22a_4
X_24052_ _24021_/CLK _24052_/D VGND VGND VPWR VPWR _24052_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22424__B2 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20215_ _24159_/Q VGND VGND VPWR VPWR _20223_/A sky130_fd_sc_hd__buf_2
X_23003_ _23003_/A _18199_/X VGND VGND VPWR VPWR _23005_/B sky130_fd_sc_hd__nand2_4
XFILLER_116_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13993__A _12598_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21195_ _20723_/X _21190_/X _23947_/Q _21194_/X VGND VGND VPWR VPWR _23947_/D sky130_fd_sc_hd__o22a_4
XFILLER_85_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20146_ IRQ[7] VGND VGND VPWR VPWR _20146_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19680__A HRDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20077_ _20090_/D _20077_/B _20076_/X _20077_/D VGND VGND VPWR VPWR _20077_/X sky130_fd_sc_hd__or4_4
XFILLER_98_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12402__A _15774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20738__B2 _20686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24472__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23905_ _23487_/CLK _23905_/D VGND VGND VPWR VPWR _15146_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_79_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18296__A _18242_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16809__A _16622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24401__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15713__A _15712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ _11850_/A VGND VGND VPWR VPWR _13491_/A sky130_fd_sc_hd__buf_2
X_23836_ _23840_/CLK _21407_/X VGND VGND VPWR VPWR _23836_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11781_ _11780_/X _11781_/B VGND VGND VPWR VPWR _11782_/C sky130_fd_sc_hd__or2_4
X_23767_ _23316_/CLK _21523_/X VGND VGND VPWR VPWR _16171_/B sky130_fd_sc_hd__dfxtp_4
X_20979_ _20913_/A _20979_/B VGND VGND VPWR VPWR _20979_/X sky130_fd_sc_hd__or2_4
XANTENNA__14329__A _14322_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13520_ _13558_/A _13453_/B VGND VGND VPWR VPWR _13522_/B sky130_fd_sc_hd__or2_4
XANTENNA__13233__A _13257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22718_ _19108_/A VGND VGND VPWR VPWR _22967_/A sky130_fd_sc_hd__inv_2
X_23698_ _23698_/CLK _21657_/X VGND VGND VPWR VPWR _13122_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13451_ _13447_/X _13451_/B _13451_/C VGND VGND VPWR VPWR _13452_/C sky130_fd_sc_hd__and3_4
XFILLER_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22649_ _22437_/X _22643_/X _13966_/B _22647_/X VGND VGND VPWR VPWR _22649_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16544__A _11886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12402_ _15774_/A _12402_/B _12402_/C VGND VGND VPWR VPWR _12406_/B sky130_fd_sc_hd__and3_4
X_16170_ _16201_/A _16096_/B VGND VGND VPWR VPWR _16170_/X sky130_fd_sc_hd__or2_4
XANTENNA__21466__A2 _21463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13382_ _13358_/X _23664_/Q VGND VGND VPWR VPWR _13384_/B sky130_fd_sc_hd__or2_4
XFILLER_70_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22663__B2 _22626_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15121_ _14986_/X VGND VGND VPWR VPWR _15121_/X sky130_fd_sc_hd__buf_2
XANTENNA__11688__A _15774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12333_ _12747_/A _12331_/X _12332_/X VGND VGND VPWR VPWR _12333_/X sky130_fd_sc_hd__and3_4
X_24319_ _24320_/CLK _24319_/D HRESETn VGND VGND VPWR VPWR _24319_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15052_ _12341_/A _15052_/B VGND VGND VPWR VPWR _15054_/B sky130_fd_sc_hd__or2_4
X_12264_ _12255_/X _12259_/X _12263_/X VGND VGND VPWR VPWR _12264_/X sky130_fd_sc_hd__and3_4
XFILLER_108_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14999__A _15019_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22074__A2_N _22072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14003_ _14026_/A VGND VGND VPWR VPWR _14845_/A sky130_fd_sc_hd__buf_2
XFILLER_68_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12195_ _13982_/A VGND VGND VPWR VPWR _12196_/A sky130_fd_sc_hd__buf_2
X_19860_ _19585_/X _19859_/X _22017_/B _19678_/X VGND VGND VPWR VPWR _19860_/X sky130_fd_sc_hd__o22a_4
X_18811_ _12100_/X _12101_/X _12036_/X _12051_/X VGND VGND VPWR VPWR _18812_/D sky130_fd_sc_hd__or4_4
X_19791_ _19622_/Y _19785_/Y _19429_/A _19790_/X VGND VGND VPWR VPWR _19791_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13408__A _12822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15954_ _15980_/A _15946_/X _15954_/C VGND VGND VPWR VPWR _15954_/X sky130_fd_sc_hd__or3_4
X_18742_ _18728_/A _19941_/B VGND VGND VPWR VPWR _19943_/B sky130_fd_sc_hd__nor2_4
XANTENNA__12312__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21926__B1 _23548_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14905_ _15146_/A _14905_/B VGND VGND VPWR VPWR _14905_/X sky130_fd_sc_hd__or2_4
XFILLER_37_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18673_ _18392_/A _17937_/X VGND VGND VPWR VPWR _18673_/Y sky130_fd_sc_hd__nor2_4
XFILLER_97_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13127__B _24082_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15885_ _13550_/A _15883_/X _15884_/X VGND VGND VPWR VPWR _15889_/B sky130_fd_sc_hd__and3_4
XFILLER_110_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12031__B _12031_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24142__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15623__A _15623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14836_ _14050_/A _14834_/X _14835_/X VGND VGND VPWR VPWR _14836_/X sky130_fd_sc_hd__and3_4
X_17624_ _17623_/X VGND VGND VPWR VPWR _18274_/C sky130_fd_sc_hd__inv_2
XFILLER_79_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17555_ _17164_/X _17572_/B VGND VGND VPWR VPWR _18066_/B sky130_fd_sc_hd__and2_4
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14767_ _13800_/A _14765_/X _14766_/X VGND VGND VPWR VPWR _14767_/X sky130_fd_sc_hd__and3_4
X_11979_ _15812_/A VGND VGND VPWR VPWR _11980_/A sky130_fd_sc_hd__buf_2
XANTENNA__18934__A _18934_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16506_ _16506_/A _16504_/X _16506_/C VGND VGND VPWR VPWR _16506_/X sky130_fd_sc_hd__and3_4
XANTENNA__13143__A _12706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13718_ _13718_/A VGND VGND VPWR VPWR _15494_/A sky130_fd_sc_hd__buf_2
X_17486_ _11834_/A _17364_/X _17365_/X VGND VGND VPWR VPWR _17487_/B sky130_fd_sc_hd__o21a_4
XANTENNA__24332__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14698_ _11697_/A _14698_/B VGND VGND VPWR VPWR _14700_/B sky130_fd_sc_hd__or2_4
XFILLER_60_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22456__A _22456_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16437_ _16394_/X _16437_/B VGND VGND VPWR VPWR _16437_/X sky130_fd_sc_hd__or2_4
X_19225_ _19225_/A _19257_/A VGND VGND VPWR VPWR _19225_/X sky130_fd_sc_hd__and2_4
X_13649_ _13597_/X _13617_/X _13625_/X _13638_/X _13648_/X VGND VGND VPWR VPWR _13649_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12982__A _12982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19156_ _24310_/Q _19157_/A _19155_/Y VGND VGND VPWR VPWR _19156_/X sky130_fd_sc_hd__o21a_4
X_16368_ _11715_/A _16368_/B VGND VGND VPWR VPWR _16369_/C sky130_fd_sc_hd__or2_4
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18107_ _18107_/A VGND VGND VPWR VPWR _18107_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_51_0_HCLK clkbuf_5_25_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15319_ _15333_/A _15256_/B VGND VGND VPWR VPWR _15320_/C sky130_fd_sc_hd__or2_4
X_19087_ _18935_/X VGND VGND VPWR VPWR _19087_/X sky130_fd_sc_hd__buf_2
X_16299_ _15929_/X _16295_/X _16298_/X VGND VGND VPWR VPWR _16299_/X sky130_fd_sc_hd__or3_4
X_18038_ _17861_/A _18035_/X _17256_/A _18037_/X VGND VGND VPWR VPWR _18038_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21209__A2 _21204_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14702__A _14055_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20000_ _20000_/A VGND VGND VPWR VPWR _20000_/X sky130_fd_sc_hd__buf_2
XANTENNA__21090__B1 _15724_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19989_ _19988_/X VGND VGND VPWR VPWR _19989_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22709__A2 _22707_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12222__A _12221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21951_ _21838_/X _21945_/X _23530_/Q _21949_/X VGND VGND VPWR VPWR _23530_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16629__A _11754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21393__B2 _21387_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20902_ _20901_/Y _20708_/B VGND VGND VPWR VPWR _20902_/X sky130_fd_sc_hd__or2_4
XANTENNA__15533__A _15533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21882_ _21807_/X _21880_/X _23575_/Q _21877_/X VGND VGND VPWR VPWR _23575_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16348__B _16280_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _23845_/CLK _23621_/D VGND VGND VPWR VPWR _14480_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833_ _20833_/A VGND VGND VPWR VPWR _20833_/Y sky130_fd_sc_hd__inv_2
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14149__A _14149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21145__B2 _21144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13053__A _12211_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23552_ _23391_/CLK _21913_/X VGND VGND VPWR VPWR _23552_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21696__A2 _21691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22893__A1 _18700_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20764_ _20654_/X _20761_/Y _20763_/X _19056_/Y _20709_/X VGND VGND VPWR VPWR _20764_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22503_ _22444_/X _22500_/X _13824_/B _22497_/X VGND VGND VPWR VPWR _23207_/D sky130_fd_sc_hd__o22a_4
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20695_ _24204_/Q _20614_/X _20694_/Y VGND VGND VPWR VPWR _20696_/A sky130_fd_sc_hd__o21a_4
X_23483_ _24026_/CLK _22027_/X VGND VGND VPWR VPWR _23483_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12892__A _12892_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16364__A _16364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22434_ _20722_/A VGND VGND VPWR VPWR _22434_/X sky130_fd_sc_hd__buf_2
XANTENNA__22645__B2 _22640_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19675__A HRDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22365_ _22351_/A VGND VGND VPWR VPWR _22365_/X sky130_fd_sc_hd__buf_2
XFILLER_30_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24104_ _24229_/CLK _24104_/D HRESETn VGND VGND VPWR VPWR _19414_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__14335__B1 _14326_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21316_ _21316_/A VGND VGND VPWR VPWR _21316_/X sky130_fd_sc_hd__buf_2
X_22296_ _22141_/X _22293_/X _15255_/B _22290_/X VGND VGND VPWR VPWR _23330_/D sky130_fd_sc_hd__o22a_4
XFILLER_105_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16905__A1_N _16897_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20614__A _20512_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21247_ _21247_/A VGND VGND VPWR VPWR _21247_/X sky130_fd_sc_hd__buf_2
X_24035_ _23270_/CLK _21053_/X VGND VGND VPWR VPWR _14759_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17195__A _17194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15708__A _12747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20959__A1 _20872_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20959__B2 _20202_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21081__B1 _24020_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21178_ _20442_/X _21176_/X _23959_/Q _21173_/X VGND VGND VPWR VPWR _21178_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21620__A2 _21619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20129_ _18689_/Y _19936_/X _20128_/X VGND VGND VPWR VPWR _20129_/X sky130_fd_sc_hd__o21a_4
XFILLER_24_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12951_ _12951_/A _12951_/B _12950_/X VGND VGND VPWR VPWR _12951_/X sky130_fd_sc_hd__and3_4
XFILLER_100_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16539__A _12024_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21384__B2 _21380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22581__B1 _16186_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11902_ _11901_/X VGND VGND VPWR VPWR _11903_/A sky130_fd_sc_hd__buf_2
XFILLER_73_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15443__A _15443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15670_ _15693_/A _15670_/B VGND VGND VPWR VPWR _15670_/X sky130_fd_sc_hd__or2_4
X_12882_ _13960_/A VGND VGND VPWR VPWR _12883_/A sky130_fd_sc_hd__buf_2
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14621_ _14734_/A _14618_/X _14620_/X VGND VGND VPWR VPWR _14621_/X sky130_fd_sc_hd__and3_4
X_11833_ _11782_/A _11831_/X _11833_/C VGND VGND VPWR VPWR _11833_/X sky130_fd_sc_hd__and3_4
X_23819_ _23819_/CLK _23819_/D VGND VGND VPWR VPWR _15560_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14059__A _11647_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21136__B2 _21130_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17340_ _17012_/A VGND VGND VPWR VPWR _17340_/X sky130_fd_sc_hd__buf_2
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24060__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _13711_/X _14550_/X _14551_/X VGND VGND VPWR VPWR _14552_/X sky130_fd_sc_hd__and3_4
XANTENNA__18001__B2 _18000_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _14175_/A VGND VGND VPWR VPWR _14020_/A sky130_fd_sc_hd__inv_2
XFILLER_53_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22276__A _22269_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _12959_/A VGND VGND VPWR VPWR _15892_/A sky130_fd_sc_hd__buf_2
XANTENNA__23628__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21180__A _21180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17270_/X VGND VGND VPWR VPWR _17271_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13898__A _13910_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14483_ _13614_/A _14547_/B VGND VGND VPWR VPWR _14483_/X sky130_fd_sc_hd__or2_4
XANTENNA__16563__A1 _16741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _13839_/A VGND VGND VPWR VPWR _14247_/A sky130_fd_sc_hd__buf_2
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19010_ _19010_/A VGND VGND VPWR VPWR _19010_/Y sky130_fd_sc_hd__inv_2
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16222_ _16198_/A _16222_/B _16221_/X VGND VGND VPWR VPWR _16230_/B sky130_fd_sc_hd__or3_4
XFILLER_35_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13434_ _13427_/A _13434_/B VGND VGND VPWR VPWR _13434_/X sky130_fd_sc_hd__or2_4
XANTENNA__21439__A2 _21433_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16153_ _11852_/X _16153_/B VGND VGND VPWR VPWR _16153_/X sky130_fd_sc_hd__and2_4
X_13365_ _13354_/X _23760_/Q VGND VGND VPWR VPWR _13366_/C sky130_fd_sc_hd__or2_4
XANTENNA__12307__A _12307_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15104_ _15104_/A _15102_/X _15103_/X VGND VGND VPWR VPWR _15108_/B sky130_fd_sc_hd__and3_4
X_12316_ _15693_/A _12316_/B VGND VGND VPWR VPWR _12316_/X sky130_fd_sc_hd__or2_4
X_16084_ _16096_/A _16158_/B VGND VGND VPWR VPWR _16084_/X sky130_fd_sc_hd__or2_4
X_13296_ _13301_/A _13296_/B VGND VGND VPWR VPWR _13296_/X sky130_fd_sc_hd__or2_4
XFILLER_108_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16721__B _23835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15035_ _14748_/A _15035_/B _15035_/C VGND VGND VPWR VPWR _15039_/B sky130_fd_sc_hd__and3_4
X_19912_ _19909_/X _24151_/Q _19910_/X _20400_/B VGND VGND VPWR VPWR _19912_/X sky130_fd_sc_hd__o22a_4
XFILLER_68_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12247_ _12240_/A VGND VGND VPWR VPWR _12726_/A sky130_fd_sc_hd__buf_2
XANTENNA__14522__A _13747_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24394__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19843_ _19678_/A _19837_/X _19840_/Y _21162_/C _19531_/A VGND VGND VPWR VPWR _19844_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_69_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21611__A2 _21605_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12178_ _11829_/A _23645_/Q VGND VGND VPWR VPWR _12179_/C sky130_fd_sc_hd__or2_4
XFILLER_64_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13138__A _12691_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17291__A2 _17012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19774_ _19541_/A _19773_/X _19669_/Y VGND VGND VPWR VPWR _19774_/X sky130_fd_sc_hd__o21a_4
XFILLER_81_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16986_ _16942_/Y _16985_/X VGND VGND VPWR VPWR _16986_/X sky130_fd_sc_hd__or2_4
XFILLER_110_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18725_ _18650_/X _18724_/X _20180_/A _18650_/X VGND VGND VPWR VPWR _24448_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21355__A _21369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15937_ _13303_/X VGND VGND VPWR VPWR _15937_/X sky130_fd_sc_hd__buf_2
XANTENNA__21375__B2 _21373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11881__A _14283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15868_ _13548_/X _15799_/B VGND VGND VPWR VPWR _15869_/C sky130_fd_sc_hd__or2_4
X_18656_ _18656_/A _18656_/B VGND VGND VPWR VPWR _18656_/X sky130_fd_sc_hd__or2_4
X_14819_ _13872_/A _14819_/B VGND VGND VPWR VPWR _14821_/B sky130_fd_sc_hd__or2_4
X_17607_ _18621_/B _17606_/X VGND VGND VPWR VPWR _17607_/X sky130_fd_sc_hd__or2_4
X_15799_ _12865_/A _15799_/B VGND VGND VPWR VPWR _15799_/X sky130_fd_sc_hd__or2_4
X_18587_ _18499_/X _18587_/B VGND VGND VPWR VPWR _18587_/X sky130_fd_sc_hd__and2_4
XFILLER_45_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21127__B2 _21123_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17538_ _17628_/A VGND VGND VPWR VPWR _17540_/A sky130_fd_sc_hd__inv_2
XANTENNA__21678__A2 _21676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22186__A _22153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17469_ _17662_/B VGND VGND VPWR VPWR _17469_/Y sky130_fd_sc_hd__inv_2
X_19208_ _24259_/Q _19208_/B VGND VGND VPWR VPWR _19209_/B sky130_fd_sc_hd__and2_4
X_20480_ _18193_/X _20424_/X _20290_/X _20479_/Y VGND VGND VPWR VPWR _20481_/A sky130_fd_sc_hd__a211o_4
XANTENNA__20638__B1 _15697_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19139_ _19139_/A VGND VGND VPWR VPWR _20244_/A sky130_fd_sc_hd__inv_2
XANTENNA__19495__A HRDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12217__A _12217_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22150_ _21583_/A VGND VGND VPWR VPWR _22383_/C sky130_fd_sc_hd__buf_2
XFILLER_69_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17727__B _17300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21101_ _20838_/X _21096_/X _14278_/B _21100_/X VGND VGND VPWR VPWR _24006_/D sky130_fd_sc_hd__o22a_4
X_22081_ _20355_/A VGND VGND VPWR VPWR _22081_/X sky130_fd_sc_hd__buf_2
XFILLER_86_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21032_ _20553_/X _21030_/X _24050_/Q _21027_/X VGND VGND VPWR VPWR _24050_/D sky130_fd_sc_hd__o22a_4
XFILLER_87_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_58_0_HCLK clkbuf_7_58_0_HCLK/A VGND VGND VPWR VPWR _23794_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__13048__A _13048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21790__A2_N _21788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22983_ _22955_/X _17681_/A _22967_/X _22982_/X VGND VGND VPWR VPWR _22984_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16359__A _11702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11791__A _11780_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15263__A _14143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21934_ _21809_/X _21931_/X _12263_/B _21928_/X VGND VGND VPWR VPWR _21934_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16078__B _16077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21865_ _23582_/Q VGND VGND VPWR VPWR _21865_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _23315_/CLK _21815_/X VGND VGND VPWR VPWR _23604_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ _20913_/A _20815_/X VGND VGND VPWR VPWR _20816_/X sky130_fd_sc_hd__or2_4
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21796_ _21795_/X _21793_/X _23612_/Q _21788_/X VGND VGND VPWR VPWR _23612_/D sky130_fd_sc_hd__o22a_4
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22096__A _22108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23535_ _23311_/CLK _23535_/D VGND VGND VPWR VPWR _23535_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15710__B _15709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20747_ _20747_/A VGND VGND VPWR VPWR _20748_/A sky130_fd_sc_hd__buf_2
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14607__A _14113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13511__A _12951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23466_ _23819_/CLK _22051_/X VGND VGND VPWR VPWR _23466_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20678_ _22821_/A _20676_/X _20677_/X VGND VGND VPWR VPWR _20678_/X sky130_fd_sc_hd__and3_4
XFILLER_104_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22824__A _18759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22417_ _22415_/X _22416_/X _12925_/B _22411_/X VGND VGND VPWR VPWR _22417_/X sky130_fd_sc_hd__o22a_4
XANTENNA__13230__B _23985_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22094__A2 _22089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23397_ _23365_/CLK _22192_/X VGND VGND VPWR VPWR _14473_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12127__A _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13150_ _15687_/A _13150_/B _13149_/X VGND VGND VPWR VPWR _13150_/X sky130_fd_sc_hd__and3_4
X_22348_ _22088_/X _22347_/X _15952_/B _22344_/X VGND VGND VPWR VPWR _23288_/D sky130_fd_sc_hd__o22a_4
XFILLER_109_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12101_ _12008_/A VGND VGND VPWR VPWR _12101_/X sky130_fd_sc_hd__buf_2
XANTENNA__19771__A1_N _19674_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15438__A _13670_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13081_ _13096_/A _13078_/X _13081_/C VGND VGND VPWR VPWR _13082_/C sky130_fd_sc_hd__and3_4
X_22279_ _22272_/A VGND VGND VPWR VPWR _22279_/X sky130_fd_sc_hd__buf_2
XFILLER_105_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12032_ _11837_/X VGND VGND VPWR VPWR _18728_/A sky130_fd_sc_hd__inv_2
X_24018_ _24082_/CLK _21084_/X VGND VGND VPWR VPWR _24018_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_105_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17653__A _16985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16840_ _13776_/X _16840_/B _16840_/C VGND VGND VPWR VPWR _16840_/X sky130_fd_sc_hd__or3_4
XFILLER_93_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16771_ _11834_/A _16771_/B _16770_/X VGND VGND VPWR VPWR _16779_/B sky130_fd_sc_hd__or3_4
X_13983_ _13983_/A _23690_/Q VGND VGND VPWR VPWR _13985_/B sky130_fd_sc_hd__or2_4
XFILLER_77_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12797__A _12813_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16269__A _11933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21357__B2 _21352_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15722_ _13130_/A _15722_/B VGND VGND VPWR VPWR _15722_/X sky130_fd_sc_hd__or2_4
X_18510_ _17706_/X _18509_/X _17706_/X _18509_/X VGND VGND VPWR VPWR _18510_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15173__A _14161_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12934_ _12596_/A _12932_/X _12933_/X VGND VGND VPWR VPWR _12934_/X sky130_fd_sc_hd__and3_4
X_19490_ _19490_/A VGND VGND VPWR VPWR _19490_/X sky130_fd_sc_hd__buf_2
X_15653_ _12691_/A _15715_/B VGND VGND VPWR VPWR _15653_/X sky130_fd_sc_hd__or2_4
X_18441_ _18264_/A _17432_/B VGND VGND VPWR VPWR _18444_/B sky130_fd_sc_hd__and2_4
X_12865_ _12865_/A _23283_/Q VGND VGND VPWR VPWR _12865_/X sky130_fd_sc_hd__or2_4
XFILLER_76_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21109__B2 _21072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14604_ _14752_/A _14604_/B _14603_/X VGND VGND VPWR VPWR _14605_/B sky130_fd_sc_hd__or3_4
XFILLER_2_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11816_ _11824_/A _11812_/X _11815_/X VGND VGND VPWR VPWR _11816_/X sky130_fd_sc_hd__or3_4
X_18372_ _17792_/A _18274_/C _17259_/A _18153_/A VGND VGND VPWR VPWR _18373_/B sky130_fd_sc_hd__o22a_4
X_15584_ _15584_/A _23499_/Q VGND VGND VPWR VPWR _15585_/C sky130_fd_sc_hd__or2_4
XFILLER_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22857__A1 _17560_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12796_ _12803_/A _12711_/B VGND VGND VPWR VPWR _12796_/X sky130_fd_sc_hd__or2_4
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _15379_/X _17114_/A VGND VGND VPWR VPWR _17323_/X sky130_fd_sc_hd__or2_4
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14554_/A _14535_/B VGND VGND VPWR VPWR _14537_/B sky130_fd_sc_hd__or2_4
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11746_/X VGND VGND VPWR VPWR _11747_/X sky130_fd_sc_hd__buf_2
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17254_ _17249_/A _17845_/A VGND VGND VPWR VPWR _17254_/X sky130_fd_sc_hd__or2_4
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ _12885_/A _14536_/B VGND VGND VPWR VPWR _14467_/C sky130_fd_sc_hd__or2_4
XANTENNA__22609__B2 _22604_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _14816_/A VGND VGND VPWR VPWR _13908_/A sky130_fd_sc_hd__buf_2
XFILLER_105_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16205_ _16193_/A _24055_/Q VGND VGND VPWR VPWR _16206_/C sky130_fd_sc_hd__or2_4
XFILLER_30_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13417_ _13397_/X _24080_/Q VGND VGND VPWR VPWR _13417_/X sky130_fd_sc_hd__or2_4
X_17185_ _17151_/X _17177_/X _17160_/X _17184_/X VGND VGND VPWR VPWR _17185_/Y sky130_fd_sc_hd__a22oi_4
X_14397_ _14397_/A _14392_/X _14397_/C VGND VGND VPWR VPWR _14397_/X sky130_fd_sc_hd__or3_4
XANTENNA__12037__A _11924_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16732__A _12100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16136_ _16140_/A _16134_/X _16136_/C VGND VGND VPWR VPWR _16137_/C sky130_fd_sc_hd__and3_4
X_13348_ _11980_/A _13324_/X _13331_/X _13339_/X _13347_/X VGND VGND VPWR VPWR _13348_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21832__A2 _21829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20254__A _20253_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16067_ _11684_/X _16067_/B _16066_/X VGND VGND VPWR VPWR _16075_/B sky130_fd_sc_hd__or3_4
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13279_ _13202_/X _13278_/X _13273_/Y VGND VGND VPWR VPWR _13280_/B sky130_fd_sc_hd__a21o_4
XANTENNA__14252__A _14252_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15018_ _13987_/A _14995_/X _15002_/X _15009_/X _15017_/X VGND VGND VPWR VPWR _15018_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_44_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19762__B HRDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18659__A _18713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21596__B2 _21595_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19826_ _19829_/A _19826_/B VGND VGND VPWR VPWR _19827_/C sky130_fd_sc_hd__or2_4
XFILLER_69_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19757_ _19755_/Y _19789_/B _19486_/Y VGND VGND VPWR VPWR _19757_/X sky130_fd_sc_hd__o21a_4
X_16969_ _16969_/A _16969_/B VGND VGND VPWR VPWR _16970_/B sky130_fd_sc_hd__or2_4
XANTENNA__16179__A _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22545__B1 _15852_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15083__A _15107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18708_ _16925_/Y _18703_/Y _16924_/X _19356_/A VGND VGND VPWR VPWR _18708_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21899__A2 _21894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19688_ _19468_/X _19829_/A _19726_/B VGND VGND VPWR VPWR _19689_/A sky130_fd_sc_hd__o21a_4
XANTENNA__12500__A _13016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22909__A _23027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18639_ _18697_/A _17306_/A _18635_/X _18638_/Y VGND VGND VPWR VPWR _18639_/X sky130_fd_sc_hd__a211o_4
XFILLER_92_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15811__A _12891_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21650_ _21522_/X _21648_/X _16219_/B _21645_/X VGND VGND VPWR VPWR _23703_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22848__A1 _17466_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19713__A1 _20490_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16626__B _23580_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20601_ _20518_/X _20600_/X _24335_/Q _20525_/X VGND VGND VPWR VPWR _20601_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15530__B _15530_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21581_ _21581_/A VGND VGND VPWR VPWR _21684_/A sky130_fd_sc_hd__buf_2
XFILLER_60_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20323__A2 _18814_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23320_ _23320_/CLK _23320_/D VGND VGND VPWR VPWR _15960_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13331__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20532_ _20376_/X _20514_/X _20515_/X _20531_/Y VGND VGND VPWR VPWR _20532_/X sky130_fd_sc_hd__a211o_4
XFILLER_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20463_ _20463_/A VGND VGND VPWR VPWR _20464_/A sky130_fd_sc_hd__buf_2
X_23251_ _23986_/CLK _22417_/X VGND VGND VPWR VPWR _12925_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_14_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22202_ _22201_/X VGND VGND VPWR VPWR _22207_/A sky130_fd_sc_hd__buf_2
Xclkbuf_5_21_0_HCLK clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20394_ _21802_/A VGND VGND VPWR VPWR _20394_/X sky130_fd_sc_hd__buf_2
X_23182_ _23692_/CLK _22544_/X VGND VGND VPWR VPWR _15659_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_119_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22133_ _22131_/X _22125_/X _14296_/B _22132_/X VGND VGND VPWR VPWR _23430_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15258__A _14145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14162__A _14737_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24449__CLK _24203_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22064_ _21861_/X _22059_/X _23456_/Q _22020_/X VGND VGND VPWR VPWR _23456_/D sky130_fd_sc_hd__o22a_4
XFILLER_102_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21015_ _21015_/A VGND VGND VPWR VPWR _21030_/A sky130_fd_sc_hd__buf_2
XANTENNA__17473__A _12676_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16089__A _12546_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21339__B2 _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13506__A _13494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22000__A2 _21995_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22966_ _22966_/A VGND VGND VPWR VPWR HADDR[14] sky130_fd_sc_hd__inv_2
XFILLER_28_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20547__C1 _20546_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21917_ _21684_/A _21917_/B _21684_/C _21866_/D VGND VGND VPWR VPWR _21917_/X sky130_fd_sc_hd__or4_4
XFILLER_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21723__A _21702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22897_ _22886_/X _22896_/X _18610_/A _22892_/X VGND VGND VPWR VPWR _22897_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15721__A _13129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12650_ _12650_/A VGND VGND VPWR VPWR _12976_/A sky130_fd_sc_hd__buf_2
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22839__A1 _13059_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21848_ _21812_/A VGND VGND VPWR VPWR _21848_/X sky130_fd_sc_hd__buf_2
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20339__A _21795_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _11601_/A VGND VGND VPWR VPWR _18866_/B sky130_fd_sc_hd__buf_2
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _14002_/A VGND VGND VPWR VPWR _12582_/A sky130_fd_sc_hd__buf_2
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21779_ _21572_/X _21776_/X _15300_/B _21773_/X VGND VGND VPWR VPWR _23618_/D sky130_fd_sc_hd__o22a_4
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14337__A _11669_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21511__B2 _21503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14320_ _14432_/A _14320_/B VGND VGND VPWR VPWR _14321_/C sky130_fd_sc_hd__or2_4
XFILLER_15_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13241__A _13260_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ _11532_/A _11531_/X VGND VGND VPWR VPWR _11532_/X sky130_fd_sc_hd__or2_4
X_23518_ _23320_/CLK _23518_/D VGND VGND VPWR VPWR _23518_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22554__A _22533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _14251_/A _23465_/Q VGND VGND VPWR VPWR _14251_/X sky130_fd_sc_hd__or2_4
XFILLER_8_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23449_ _23354_/CLK _23449_/D VGND VGND VPWR VPWR _16267_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_32_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13202_ _12189_/X _12681_/X _13170_/X _12281_/X _13201_/X VGND VGND VPWR VPWR _13202_/X
+ sky130_fd_sc_hd__a32o_4
X_14182_ _14182_/A _23497_/Q VGND VGND VPWR VPWR _14183_/C sky130_fd_sc_hd__or2_4
XANTENNA__20074__A _11622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13133_ _13133_/A _13133_/B _13133_/C VGND VGND VPWR VPWR _13133_/X sky130_fd_sc_hd__and3_4
XANTENNA__15168__A _14145_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18691__A1 _17989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18990_ _24340_/Q _11524_/X _18983_/Y VGND VGND VPWR VPWR _18990_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__14072__A _14040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13064_ _13104_/A _13064_/B VGND VGND VPWR VPWR _13067_/B sky130_fd_sc_hd__or2_4
X_17941_ _18327_/A _17577_/X _17874_/X _17629_/Y VGND VGND VPWR VPWR _17942_/B sky130_fd_sc_hd__o22a_4
XFILLER_117_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12015_ _16536_/A _23646_/Q VGND VGND VPWR VPWR _12016_/C sky130_fd_sc_hd__or2_4
XANTENNA__17383__A _13837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17872_ _17794_/X _17853_/Y _17856_/X _17871_/X VGND VGND VPWR VPWR _17872_/X sky130_fd_sc_hd__a211o_4
XFILLER_78_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14800__A _13706_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19611_ _19537_/A _19610_/X VGND VGND VPWR VPWR _19611_/X sky130_fd_sc_hd__and2_4
XFILLER_66_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_41_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR _23079_/CLK sky130_fd_sc_hd__clkbuf_1
X_16823_ _15926_/D VGND VGND VPWR VPWR _16824_/D sky130_fd_sc_hd__buf_2
XFILLER_94_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15615__B _23947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22527__B1 _16387_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19542_ _19499_/Y _19877_/B _19582_/A VGND VGND VPWR VPWR _19542_/X sky130_fd_sc_hd__o21a_4
X_13966_ _13966_/A _13966_/B VGND VGND VPWR VPWR _13966_/X sky130_fd_sc_hd__or2_4
X_16754_ _16629_/X _16754_/B VGND VGND VPWR VPWR _16754_/X sky130_fd_sc_hd__or2_4
XFILLER_93_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12320__A _12320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20002__A1 _18196_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12917_ _12917_/A _12915_/X _12916_/X VGND VGND VPWR VPWR _12921_/B sky130_fd_sc_hd__and3_4
X_15705_ _12744_/A _15703_/X _15705_/C VGND VGND VPWR VPWR _15705_/X sky130_fd_sc_hd__and3_4
XFILLER_39_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16685_ _16718_/A _16683_/X _16685_/C VGND VGND VPWR VPWR _16685_/X sky130_fd_sc_hd__and3_4
X_19473_ _24155_/Q _19459_/X HRDATA[29] _19460_/X VGND VGND VPWR VPWR _19473_/X sky130_fd_sc_hd__o22a_4
X_13897_ _13890_/A _23367_/Q VGND VGND VPWR VPWR _13899_/B sky130_fd_sc_hd__or2_4
XFILLER_111_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21750__B2 _21745_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18424_ _18107_/A VGND VGND VPWR VPWR _18424_/X sky130_fd_sc_hd__buf_2
XFILLER_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12848_ _12444_/A _23507_/Q VGND VGND VPWR VPWR _12849_/C sky130_fd_sc_hd__or2_4
X_15636_ _15601_/A _23467_/Q VGND VGND VPWR VPWR _15636_/X sky130_fd_sc_hd__or2_4
XANTENNA__20249__A _20301_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15567_ _14432_/A _24075_/Q VGND VGND VPWR VPWR _15567_/X sky130_fd_sc_hd__or2_4
X_18355_ _18354_/X VGND VGND VPWR VPWR _18355_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12779_ _13088_/A VGND VGND VPWR VPWR _15724_/A sky130_fd_sc_hd__buf_2
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13151__A _13317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14518_ _13695_/X _14518_/B VGND VGND VPWR VPWR _14518_/X sky130_fd_sc_hd__or2_4
X_17306_ _17306_/A _17305_/Y VGND VGND VPWR VPWR _17306_/X sky130_fd_sc_hd__or2_4
XFILLER_33_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15498_ _13737_/A _15496_/X _15497_/X VGND VGND VPWR VPWR _15499_/C sky130_fd_sc_hd__and3_4
X_18286_ _18286_/A _18285_/X VGND VGND VPWR VPWR _18286_/X sky130_fd_sc_hd__and2_4
X_14449_ _13019_/A _22325_/A VGND VGND VPWR VPWR _14451_/B sky130_fd_sc_hd__or2_4
X_17237_ _17860_/A _17200_/X _17256_/A _17236_/X VGND VGND VPWR VPWR _17238_/A sky130_fd_sc_hd__o22a_4
XANTENNA__22058__A2 _22052_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12990__A _12989_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17168_ _17151_/X _17159_/X _17160_/X _17167_/X VGND VGND VPWR VPWR _17168_/Y sky130_fd_sc_hd__a22oi_4
X_16119_ _16146_/A _16189_/B VGND VGND VPWR VPWR _16120_/C sky130_fd_sc_hd__or2_4
XFILLER_66_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17099_ _17173_/A VGND VGND VPWR VPWR _17161_/A sky130_fd_sc_hd__buf_2
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21018__B1 _24060_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23496__CLK _23079_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18389__A _18266_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21569__B2 _21563_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17293__A _14565_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15806__A _12852_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22230__A2 _22229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19809_ _19524_/B VGND VGND VPWR VPWR _19809_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15525__B _23339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22820_ _22813_/X _22820_/B VGND VGND VPWR VPWR HWDATA[14] sky130_fd_sc_hd__nor2_4
XFILLER_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12230__A _13017_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22751_ _22727_/A _24097_/Q VGND VGND VPWR VPWR _22751_/X sky130_fd_sc_hd__or2_4
XFILLER_80_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21702_ _21702_/A VGND VGND VPWR VPWR _21702_/X sky130_fd_sc_hd__buf_2
XFILLER_77_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22682_ _20464_/A _22679_/X _12328_/B _22676_/X VGND VGND VPWR VPWR _23094_/D sky130_fd_sc_hd__o22a_4
XFILLER_90_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24421_ _24320_/CLK _24421_/D HRESETn VGND VGND VPWR VPWR _20855_/A sky130_fd_sc_hd__dfrtp_4
X_21633_ _23710_/Q VGND VGND VPWR VPWR _21633_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15260__B _15260_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19698__B1 _12036_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22297__A2 _22293_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14157__A _15006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13061__A _13087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24352_ _24425_/CLK _24352_/D HRESETn VGND VGND VPWR VPWR _20968_/A sky130_fd_sc_hd__dfstp_4
XFILLER_100_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21564_ _21562_/X _21556_/X _14276_/B _21563_/X VGND VGND VPWR VPWR _21564_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19667__B _19667_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23303_ _24008_/CLK _23303_/D VGND VGND VPWR VPWR _13794_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20515_ _20515_/A VGND VGND VPWR VPWR _20515_/X sky130_fd_sc_hd__buf_2
XANTENNA__13996__A _12568_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24283_ _24344_/CLK _24283_/D HRESETn VGND VGND VPWR VPWR _19232_/A sky130_fd_sc_hd__dfrtp_4
X_21495_ _21289_/X _21491_/X _15177_/B _21452_/X VGND VGND VPWR VPWR _23777_/D sky130_fd_sc_hd__o22a_4
XFILLER_14_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16372__A _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24271__CLK _24092_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23234_ _24065_/CLK _23234_/D VGND VGND VPWR VPWR _15252_/B sky130_fd_sc_hd__dfxtp_4
X_20446_ _20229_/A _20445_/X _20284_/X VGND VGND VPWR VPWR _20446_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_119_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19683__A _19784_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23165_ _24092_/CLK _23165_/D VGND VGND VPWR VPWR _12139_/B sky130_fd_sc_hd__dfxtp_4
X_20377_ _20285_/X _20754_/A _20286_/X VGND VGND VPWR VPWR _20377_/X sky130_fd_sc_hd__a21o_4
XANTENNA__19870__B1 _20206_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20480__A1 _18193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22821__B _17283_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22116_ _22115_/X _22113_/X _15864_/B _22108_/X VGND VGND VPWR VPWR _23437_/D sky130_fd_sc_hd__o22a_4
X_23096_ _24088_/CLK _22680_/X VGND VGND VPWR VPWR _23096_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22047_ _21831_/X _22045_/X _15828_/B _22042_/X VGND VGND VPWR VPWR _23469_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22221__A2 _22215_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_28_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_28_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17451__A1_N _12752_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13820_ _15435_/A _13816_/X _13820_/C VGND VGND VPWR VPWR _13820_/X sky130_fd_sc_hd__or3_4
XANTENNA__13236__A _15484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21980__B2 _21978_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23998_ _23774_/CLK _23998_/D VGND VGND VPWR VPWR _21110_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_1_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23219__CLK _23155_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13751_ _12935_/A _13664_/B VGND VGND VPWR VPWR _13753_/B sky130_fd_sc_hd__or2_4
XANTENNA__21453__A _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22949_ _22962_/A _22949_/B VGND VGND VPWR VPWR _22952_/B sky130_fd_sc_hd__nand2_4
XANTENNA__21732__B2 _21687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12702_ _15664_/A _12699_/X _12702_/C VGND VGND VPWR VPWR _12706_/B sky130_fd_sc_hd__and3_4
X_16470_ _16363_/X _16466_/X _16470_/C VGND VGND VPWR VPWR _16480_/B sky130_fd_sc_hd__or3_4
X_13682_ _13682_/A _13682_/B VGND VGND VPWR VPWR _13682_/X sky130_fd_sc_hd__and2_4
XANTENNA__16266__B _16266_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15421_ _13597_/X _15398_/X _15405_/X _15412_/X _15420_/X VGND VGND VPWR VPWR _15421_/X
+ sky130_fd_sc_hd__a32o_4
X_12633_ _12622_/X _12633_/B VGND VGND VPWR VPWR _12634_/C sky130_fd_sc_hd__or2_4
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22288__A2 _22286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18762__A _18762_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20299__A1 _20407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15352_ _14810_/A _15352_/B VGND VGND VPWR VPWR _15353_/C sky130_fd_sc_hd__or2_4
X_18140_ _18140_/A VGND VGND VPWR VPWR _18140_/Y sky130_fd_sc_hd__inv_2
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20299__B2 _20253_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12564_ _12965_/A _12564_/B VGND VGND VPWR VPWR _12564_/X sky130_fd_sc_hd__or2_4
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ _12307_/A _14301_/X _14303_/C VGND VGND VPWR VPWR _14303_/X sky130_fd_sc_hd__and3_4
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11515_ _24330_/Q _11515_/B VGND VGND VPWR VPWR _11516_/B sky130_fd_sc_hd__or2_4
X_18071_ _17864_/A _18069_/X _17975_/A _18070_/X VGND VGND VPWR VPWR _18071_/X sky130_fd_sc_hd__o22a_4
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22715__C _20576_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15283_ _14575_/X _15283_/B VGND VGND VPWR VPWR _15283_/X sky130_fd_sc_hd__or2_4
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ _12920_/A VGND VGND VPWR VPWR _12540_/A sky130_fd_sc_hd__buf_2
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17022_ _17022_/A VGND VGND VPWR VPWR _17022_/X sky130_fd_sc_hd__buf_2
X_14234_ _14225_/A _23113_/Q VGND VGND VPWR VPWR _14237_/B sky130_fd_sc_hd__or2_4
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21248__B1 _23923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14165_ _14165_/A _23785_/Q VGND VGND VPWR VPWR _14165_/X sky130_fd_sc_hd__or2_4
XANTENNA__12315__A _12315_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13116_ _13100_/A _13116_/B _13116_/C VGND VGND VPWR VPWR _13117_/C sky130_fd_sc_hd__and3_4
XFILLER_113_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14096_ _14990_/A VGND VGND VPWR VPWR _14096_/X sky130_fd_sc_hd__buf_2
X_18973_ _11527_/X VGND VGND VPWR VPWR _18973_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13047_ _13014_/A _13045_/X _13046_/X VGND VGND VPWR VPWR _13047_/X sky130_fd_sc_hd__and3_4
X_17924_ _17225_/X VGND VGND VPWR VPWR _17925_/B sky130_fd_sc_hd__inv_2
XANTENNA__18416__A1 _18011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14530__A _12612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17855_ _17854_/X VGND VGND VPWR VPWR _17933_/A sky130_fd_sc_hd__buf_2
XFILLER_26_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18937__A _18971_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16806_ _16799_/A _16806_/B VGND VGND VPWR VPWR _16806_/X sky130_fd_sc_hd__or2_4
XFILLER_93_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13146__A _12720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17786_ _18421_/A VGND VGND VPWR VPWR _18443_/A sky130_fd_sc_hd__buf_2
XFILLER_82_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14998_ _14998_/A _14998_/B _14998_/C VGND VGND VPWR VPWR _15002_/B sky130_fd_sc_hd__and3_4
X_19525_ _19522_/X _19686_/A VGND VGND VPWR VPWR _19525_/X sky130_fd_sc_hd__or2_4
XFILLER_53_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16737_ _11943_/A _23707_/Q VGND VGND VPWR VPWR _16739_/B sky130_fd_sc_hd__or2_4
X_13949_ _11925_/Y VGND VGND VPWR VPWR _13956_/A sky130_fd_sc_hd__buf_2
XANTENNA__12985__A _12947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16457__A _11727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15361__A _11638_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19456_ _19424_/A _19455_/X HRDATA[15] _19439_/X VGND VGND VPWR VPWR _19572_/B sky130_fd_sc_hd__o22a_4
X_16668_ _16599_/X _16668_/B _16667_/X VGND VGND VPWR VPWR _16668_/X sky130_fd_sc_hd__or3_4
XANTENNA__20931__C1 _20930_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18407_ _18386_/X _18391_/Y _18393_/X _18405_/X _18406_/Y VGND VGND VPWR VPWR _18407_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_22_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15619_ _15631_/A _15619_/B _15619_/C VGND VGND VPWR VPWR _15620_/C sky130_fd_sc_hd__and3_4
X_19387_ _19385_/X _18262_/X _19385_/X _24210_/Q VGND VGND VPWR VPWR _19387_/X sky130_fd_sc_hd__a2bb2o_4
X_16599_ _16598_/X VGND VGND VPWR VPWR _16599_/X sky130_fd_sc_hd__buf_2
XFILLER_15_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_29_0_HCLK_A clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24294__CLK _24299_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18338_ _18198_/X _18335_/X _18224_/X _18337_/X VGND VGND VPWR VPWR _18338_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21589__A2_N _21588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18269_ _17962_/X _17930_/X _17964_/X VGND VGND VPWR VPWR _18269_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_15_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20300_ _20300_/A VGND VGND VPWR VPWR _20300_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21280_ _20870_/A VGND VGND VPWR VPWR _21280_/X sky130_fd_sc_hd__buf_2
X_20231_ _20421_/A VGND VGND VPWR VPWR _20515_/A sky130_fd_sc_hd__inv_2
XFILLER_85_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12225__A _12688_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20462__A1 _24214_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20162_ _11564_/X _20161_/Y VGND VGND VPWR VPWR _20162_/X sky130_fd_sc_hd__or2_4
XANTENNA__17735__B _17117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20442__A _20442_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15536__A _15536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20093_ _20093_/A VGND VGND VPWR VPWR _20093_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14440__A _14463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12879__B _23923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23921_ _23342_/CLK _21252_/X VGND VGND VPWR VPWR _13162_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_57_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21411__B1 _16280_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15255__B _15255_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21962__B2 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13056__A _13056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23852_ _23698_/CLK _21379_/X VGND VGND VPWR VPWR _23852_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22803_ _22792_/X _22803_/B VGND VGND VPWR VPWR HWDATA[9] sky130_fd_sc_hd__nor2_4
XANTENNA__19907__B2 _20342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23783_ _23079_/CLK _21487_/X VGND VGND VPWR VPWR _13829_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_77_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20995_ _20825_/X _20994_/X VGND VGND VPWR VPWR _20995_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__12895__A _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16367__A _11702_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21714__B2 _21709_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22734_ _22733_/Y _24099_/Q SYSTICKCLKDIV[2] _22756_/A VGND VGND VPWR VPWR _22734_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_57_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17394__A1 _13685_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17394__B2 _17393_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22665_ _21005_/A _21582_/A _22383_/C _21060_/A VGND VGND VPWR VPWR _22665_/X sky130_fd_sc_hd__or4_4
XFILLER_40_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24404_ _23358_/CLK _24404_/D HRESETn VGND VGND VPWR VPWR _24404_/Q sky130_fd_sc_hd__dfrtp_4
X_21616_ _21602_/A VGND VGND VPWR VPWR _21616_/X sky130_fd_sc_hd__buf_2
XFILLER_16_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17146__A1 _17143_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22596_ _22432_/X _22593_/X _15473_/B _22590_/X VGND VGND VPWR VPWR _22596_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16814__B _16814_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24335_ _24092_/CLK _24335_/D HRESETn VGND VGND VPWR VPWR _24335_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_21_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21547_ _21546_/X _21544_/X _15792_/B _21539_/X VGND VGND VPWR VPWR _23757_/D sky130_fd_sc_hd__o22a_4
XFILLER_103_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18894__A1 _12990_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14615__A _11894_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12280_ _12922_/A _12226_/X _12243_/X _12265_/X _12279_/X VGND VGND VPWR VPWR _12280_/X
+ sky130_fd_sc_hd__a32o_4
X_24266_ _24305_/CLK _24266_/D HRESETn VGND VGND VPWR VPWR _19215_/A sky130_fd_sc_hd__dfrtp_4
X_21478_ _21258_/X _21477_/X _15763_/B _21474_/X VGND VGND VPWR VPWR _23790_/D sky130_fd_sc_hd__o22a_4
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23217_ _23217_/CLK _22489_/X VGND VGND VPWR VPWR _13188_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20429_ _20425_/X _20426_/Y _20428_/X _18975_/Y _20253_/X VGND VGND VPWR VPWR _20430_/A
+ sky130_fd_sc_hd__a32o_4
X_24197_ _24473_/CLK _24197_/D HRESETn VGND VGND VPWR VPWR _24197_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24017__CLK _24082_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12135__A _11675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19843__B1 _21162_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21650__B1 _16219_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23148_ _23564_/CLK _22596_/X VGND VGND VPWR VPWR _15473_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17645__B _17535_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15970_ _15948_/A _15970_/B _15970_/C VGND VGND VPWR VPWR _15971_/C sky130_fd_sc_hd__and3_4
X_23079_ _23079_/CLK _22703_/X VGND VGND VPWR VPWR _23079_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20071__B _20071_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12789__B _23572_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14921_ _14026_/A _14857_/B VGND VGND VPWR VPWR _14922_/C sky130_fd_sc_hd__or2_4
XFILLER_62_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21953__B2 _21949_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17640_ _16991_/A _17044_/Y _16991_/A _17044_/Y VGND VGND VPWR VPWR _17640_/X sky130_fd_sc_hd__a2bb2o_4
X_14852_ _14851_/X VGND VGND VPWR VPWR _14852_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22279__A _22272_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21183__A _21183_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13803_ _13654_/A _13801_/X _13803_/C VGND VGND VPWR VPWR _13803_/X sky130_fd_sc_hd__and3_4
X_14783_ _11847_/A _14783_/B VGND VGND VPWR VPWR _14783_/X sky130_fd_sc_hd__and2_4
X_17571_ _16233_/X _17564_/B VGND VGND VPWR VPWR _17571_/Y sky130_fd_sc_hd__nand2_4
XFILLER_90_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11995_ _11995_/A _11995_/B _11995_/C VGND VGND VPWR VPWR _11995_/X sky130_fd_sc_hd__and3_4
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19310_ _19303_/X _19309_/X _20210_/A _19303_/X VGND VGND VPWR VPWR _19310_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15181__A _14617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13734_ _15495_/A _13732_/X _13733_/X VGND VGND VPWR VPWR _13738_/B sky130_fd_sc_hd__and3_4
X_16522_ _16520_/B _16521_/Y VGND VGND VPWR VPWR _16522_/Y sky130_fd_sc_hd__nor2_4
XFILLER_44_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19241_ _19233_/B VGND VGND VPWR VPWR _19241_/Y sky130_fd_sc_hd__inv_2
X_13665_ _12211_/A _23400_/Q VGND VGND VPWR VPWR _13665_/X sky130_fd_sc_hd__or2_4
X_16453_ _16506_/A _16453_/B _16453_/C VGND VGND VPWR VPWR _16453_/X sky130_fd_sc_hd__and3_4
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12616_ _12970_/A _12614_/X _12615_/X VGND VGND VPWR VPWR _12625_/B sky130_fd_sc_hd__and3_4
X_15404_ _15404_/A _15402_/X _15404_/C VGND VGND VPWR VPWR _15405_/C sky130_fd_sc_hd__and3_4
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21469__B1 _23796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16384_ _16002_/A _16384_/B VGND VGND VPWR VPWR _16384_/X sky130_fd_sc_hd__or2_4
X_19172_ _24302_/Q _19123_/B _19171_/Y VGND VGND VPWR VPWR _19172_/X sky130_fd_sc_hd__o21a_4
X_13596_ _13987_/A VGND VGND VPWR VPWR _15450_/A sky130_fd_sc_hd__buf_2
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22130__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22130__B2 _22120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16724__B _16792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15335_ _14000_/A _15276_/B VGND VGND VPWR VPWR _15335_/X sky130_fd_sc_hd__or2_4
X_18123_ _17568_/Y _18121_/X _17634_/X VGND VGND VPWR VPWR _18123_/X sky130_fd_sc_hd__o21a_4
X_12547_ _12500_/X _12668_/B VGND VGND VPWR VPWR _12548_/C sky130_fd_sc_hd__or2_4
XANTENNA__22681__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15266_ _14149_/A _15266_/B VGND VGND VPWR VPWR _15266_/X sky130_fd_sc_hd__or2_4
X_18054_ _17651_/B _18003_/X _17651_/B _18003_/X VGND VGND VPWR VPWR _18054_/X sky130_fd_sc_hd__a2bb2o_4
X_12478_ _12477_/X _12607_/B VGND VGND VPWR VPWR _12478_/X sky130_fd_sc_hd__or2_4
X_14217_ _14247_/A _14217_/B VGND VGND VPWR VPWR _14217_/X sky130_fd_sc_hd__or2_4
X_17005_ _16931_/X VGND VGND VPWR VPWR _17006_/A sky130_fd_sc_hd__buf_2
XANTENNA__18637__A1 _18082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15197_ _15190_/A _15197_/B VGND VGND VPWR VPWR _15197_/X sky130_fd_sc_hd__or2_4
XANTENNA__12045__A _11888_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22433__A2 _22428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16740__A _12112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14148_ _15026_/A VGND VGND VPWR VPWR _14149_/A sky130_fd_sc_hd__buf_2
XFILLER_4_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14079_ _14906_/A VGND VGND VPWR VPWR _14089_/A sky130_fd_sc_hd__buf_2
X_18956_ _18971_/A VGND VGND VPWR VPWR _18956_/X sky130_fd_sc_hd__buf_2
XANTENNA__14260__A _11798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24355__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22197__B2 _22162_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17907_ _17817_/X _17184_/X _17911_/A _17159_/X VGND VGND VPWR VPWR _17908_/A sky130_fd_sc_hd__o22a_4
XANTENNA__15075__B _23423_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18887_ _17164_/X _18884_/X _24376_/Q _18885_/X VGND VGND VPWR VPWR _18887_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19369__A2_N _17898_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21944__A1 _21826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21944__B2 _21942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17571__A _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17838_ _17826_/X _17203_/X _17804_/A _17212_/X VGND VGND VPWR VPWR _17838_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_6_11_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21093__A _21079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17769_ _17769_/A _17263_/Y VGND VGND VPWR VPWR _17769_/X sky130_fd_sc_hd__or2_4
XFILLER_82_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ _24150_/Q _19435_/A HRDATA[24] _19431_/X VGND VGND VPWR VPWR _19508_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20780_ _20750_/X _20779_/X _24073_/Q _20724_/X VGND VGND VPWR VPWR _24073_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17376__A1 _15910_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21172__A2 _21169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17376__B2 _17375_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22917__A _22899_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21821__A _20574_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19439_ _19438_/X VGND VGND VPWR VPWR _19439_/X sky130_fd_sc_hd__buf_2
XFILLER_22_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22450_ _22449_/X _22440_/X _14431_/B _22447_/X VGND VGND VPWR VPWR _22450_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17128__A1 _15050_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17128__B2 _17127_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22121__B2 _22120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21401_ _21416_/A VGND VGND VPWR VPWR _21401_/X sky130_fd_sc_hd__buf_2
X_22381_ _22147_/X _22354_/A _23263_/Q _22344_/A VGND VGND VPWR VPWR _23263_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14435__A _12441_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24120_ _24202_/CLK _20056_/Y HRESETn VGND VGND VPWR VPWR _16956_/A sky130_fd_sc_hd__dfrtp_4
X_21332_ _21268_/X _21326_/X _23882_/Q _21330_/X VGND VGND VPWR VPWR _23882_/D sky130_fd_sc_hd__o22a_4
XFILLER_50_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24051_ _23311_/CLK _21031_/X VGND VGND VPWR VPWR _24051_/Q sky130_fd_sc_hd__dfxtp_4
X_21263_ _21263_/A VGND VGND VPWR VPWR _21263_/X sky130_fd_sc_hd__buf_2
XANTENNA__22424__A2 _22416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19825__B1 _21112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23002_ _23001_/X VGND VGND VPWR VPWR HADDR[20] sky130_fd_sc_hd__inv_2
XANTENNA__20435__A1 _18124_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20214_ _11579_/X VGND VGND VPWR VPWR _20214_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21632__B1 _23711_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21194_ _21180_/A VGND VGND VPWR VPWR _21194_/X sky130_fd_sc_hd__buf_2
XFILLER_104_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15266__A _14149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11794__A _11772_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20145_ _24422_/Q VGND VGND VPWR VPWR _20145_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19961__A _19985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14170__A _14617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22188__B2 _22183_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19589__C1 _19554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20076_ _20076_/A _20076_/B _18940_/A VGND VGND VPWR VPWR _20076_/X sky130_fd_sc_hd__or3_4
XFILLER_85_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18577__A _16929_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17481__A _13591_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23904_ _23840_/CLK _21292_/X VGND VGND VPWR VPWR _14879_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18800__A1 _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23835_ _23867_/CLK _23835_/D VGND VGND VPWR VPWR _23835_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13514__A _12640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11780_ _11758_/X VGND VGND VPWR VPWR _11780_/X sky130_fd_sc_hd__buf_2
X_23766_ _23920_/CLK _21525_/X VGND VGND VPWR VPWR _12229_/B sky130_fd_sc_hd__dfxtp_4
X_20978_ _24224_/Q _20444_/A _20977_/X VGND VGND VPWR VPWR _20979_/B sky130_fd_sc_hd__o21a_4
XFILLER_41_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22360__B2 _22358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22717_ _19674_/X _22714_/X _22714_/X _23064_/C VGND VGND VPWR VPWR _24106_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23697_ _23564_/CLK _23697_/D VGND VGND VPWR VPWR _13196_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13450_ _13450_/A _23535_/Q VGND VGND VPWR VPWR _13451_/C sky130_fd_sc_hd__or2_4
XANTENNA__19201__A _19108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22648_ _22434_/X _22643_/X _23115_/Q _22647_/X VGND VGND VPWR VPWR _23115_/D sky130_fd_sc_hd__o22a_4
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12401_ _12828_/A _12294_/B VGND VGND VPWR VPWR _12402_/C sky130_fd_sc_hd__or2_4
X_13381_ _13370_/A _13381_/B _13380_/X VGND VGND VPWR VPWR _13381_/X sky130_fd_sc_hd__or3_4
X_22579_ _22586_/A VGND VGND VPWR VPWR _22579_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14345__A _14345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22663__A2 _22636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15120_ _14918_/X VGND VGND VPWR VPWR _15120_/Y sky130_fd_sc_hd__inv_2
X_12332_ _12315_/A _12332_/B VGND VGND VPWR VPWR _12332_/X sky130_fd_sc_hd__or2_4
X_24318_ _24290_/CLK _24318_/D HRESETn VGND VGND VPWR VPWR _19139_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15051_ _15050_/Y VGND VGND VPWR VPWR _15051_/X sky130_fd_sc_hd__buf_2
X_12263_ _15667_/A _12263_/B VGND VGND VPWR VPWR _12263_/X sky130_fd_sc_hd__or2_4
X_24249_ _24216_/CLK _24249_/D HRESETn VGND VGND VPWR VPWR _24249_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16560__A _12020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14002_ _14002_/A VGND VGND VPWR VPWR _14026_/A sky130_fd_sc_hd__buf_2
XANTENNA__14999__B _23999_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12194_ _11606_/A VGND VGND VPWR VPWR _13982_/A sky130_fd_sc_hd__buf_2
XANTENNA__20082__A _20090_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18810_ _15119_/X _18781_/A _11540_/A _18782_/A VGND VGND VPWR VPWR _24415_/D sky130_fd_sc_hd__o22a_4
XANTENNA__15176__A _14992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19790_ _19500_/X _19788_/X _19872_/B _19789_/X VGND VGND VPWR VPWR _19790_/X sky130_fd_sc_hd__a211o_4
X_18741_ _12031_/B _17016_/X _18864_/C _17023_/X VGND VGND VPWR VPWR _19941_/B sky130_fd_sc_hd__o22a_4
X_15953_ _15994_/A _15953_/B _15952_/X VGND VGND VPWR VPWR _15954_/C sky130_fd_sc_hd__and3_4
XFILLER_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12312__B _12312_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21926__B2 _21921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14904_ _14998_/A _14902_/X _14903_/X VGND VGND VPWR VPWR _14904_/X sky130_fd_sc_hd__and3_4
XANTENNA__15904__A _13507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18672_ _17324_/X _18670_/Y VGND VGND VPWR VPWR _18672_/Y sky130_fd_sc_hd__nand2_4
XFILLER_64_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15884_ _15884_/A _23821_/Q VGND VGND VPWR VPWR _15884_/X sky130_fd_sc_hd__or2_4
XFILLER_114_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17623_ _17370_/X _17594_/Y _17602_/Y _17622_/Y VGND VGND VPWR VPWR _17623_/X sky130_fd_sc_hd__or4_4
X_14835_ _14811_/A _14777_/B VGND VGND VPWR VPWR _14835_/X sky130_fd_sc_hd__or2_4
XFILLER_40_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13424__A _11800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17554_ _16008_/Y _17015_/X _17015_/X _17652_/B VGND VGND VPWR VPWR _17572_/B sky130_fd_sc_hd__a2bb2o_4
X_11978_ _11977_/X VGND VGND VPWR VPWR _15812_/A sky130_fd_sc_hd__buf_2
X_14766_ _13799_/A _14766_/B VGND VGND VPWR VPWR _14766_/X sky130_fd_sc_hd__or2_4
X_16505_ _16473_/X _24090_/Q VGND VGND VPWR VPWR _16506_/C sky130_fd_sc_hd__or2_4
XFILLER_32_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21641__A _21662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13717_ _15493_/A _24008_/Q VGND VGND VPWR VPWR _13720_/B sky130_fd_sc_hd__or2_4
X_14697_ _15114_/A _14695_/X _14697_/C VGND VGND VPWR VPWR _14697_/X sky130_fd_sc_hd__and3_4
X_17485_ _18274_/A VGND VGND VPWR VPWR _17513_/A sky130_fd_sc_hd__inv_2
XANTENNA__16735__A _11921_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19224_ _24275_/Q _19223_/X VGND VGND VPWR VPWR _19257_/A sky130_fd_sc_hd__and2_4
XANTENNA__24111__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16436_ _11872_/X _16434_/X _16435_/X VGND VGND VPWR VPWR _16436_/X sky130_fd_sc_hd__and3_4
X_13648_ _15420_/A _13648_/B VGND VGND VPWR VPWR _13648_/X sky130_fd_sc_hd__and2_4
XFILLER_60_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11879__A _11879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19155_ _19132_/B VGND VGND VPWR VPWR _19155_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18858__A1 _17297_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13579_ _13350_/Y _13425_/X VGND VGND VPWR VPWR _13579_/X sky130_fd_sc_hd__or2_4
X_16367_ _11702_/A _16289_/B VGND VGND VPWR VPWR _16369_/B sky130_fd_sc_hd__or2_4
XFILLER_34_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_2_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18106_ _18106_/A VGND VGND VPWR VPWR _18106_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15318_ _11707_/A VGND VGND VPWR VPWR _15333_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21862__B1 _23584_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16298_ _15937_/X _16296_/X _16298_/C VGND VGND VPWR VPWR _16298_/X sky130_fd_sc_hd__and3_4
X_19086_ _19074_/X _19085_/X _19074_/X _11509_/A VGND VGND VPWR VPWR _24324_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18037_ _17845_/X _17865_/X _17837_/A _18036_/X VGND VGND VPWR VPWR _18037_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17566__A _16235_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15249_ _11652_/X _15249_/B _15248_/X VGND VGND VPWR VPWR _15249_/X sky130_fd_sc_hd__and3_4
XANTENNA__19807__B1 _18759_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15086__A _14039_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21090__B2 _21086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19988_ _19970_/X _18012_/X _19976_/X _19987_/X VGND VGND VPWR VPWR _19988_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12503__A _12503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18939_ _19027_/A VGND VGND VPWR VPWR _18940_/A sky130_fd_sc_hd__inv_2
XFILLER_45_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20720__A _20534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21950_ _21835_/X _21945_/X _23531_/Q _21949_/X VGND VGND VPWR VPWR _23531_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15814__A _12443_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21393__A2 _21390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20901_ _20901_/A VGND VGND VPWR VPWR _20901_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21881_ _21804_/X _21880_/X _23576_/Q _21877_/X VGND VGND VPWR VPWR _21881_/X sky130_fd_sc_hd__o22a_4
XFILLER_23_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23620_ _23363_/CLK _23620_/D VGND VGND VPWR VPWR _14714_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_36_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20832_ _18594_/Y _20680_/X _20731_/X _20831_/Y VGND VGND VPWR VPWR _20832_/X sky130_fd_sc_hd__a211o_4
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21145__A2 _21140_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18546__B1 _17878_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22647__A _22633_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22342__B2 _22337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21551__A _21527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23551_ _23487_/CLK _21914_/X VGND VGND VPWR VPWR _23551_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20763_ _20762_/Y _20708_/B VGND VGND VPWR VPWR _20763_/X sky130_fd_sc_hd__or2_4
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16645__A _16624_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22502_ _22442_/X _22500_/X _13766_/B _22497_/X VGND VGND VPWR VPWR _23208_/D sky130_fd_sc_hd__o22a_4
XFILLER_51_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23482_ _23699_/CLK _23482_/D VGND VGND VPWR VPWR _16427_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_18_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR _24239_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20694_ _20634_/A _20693_/X VGND VGND VPWR VPWR _20694_/Y sky130_fd_sc_hd__nand2_4
XFILLER_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22433_ _22432_/X _22428_/X _15454_/B _22423_/X VGND VGND VPWR VPWR _23244_/D sky130_fd_sc_hd__o22a_4
XFILLER_13_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14165__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22645__A2 _22643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22364_ _22117_/X _22361_/X _15403_/B _22358_/X VGND VGND VPWR VPWR _22364_/X sky130_fd_sc_hd__o22a_4
X_24103_ _24320_/CLK _24103_/D HRESETn VGND VGND VPWR VPWR _22772_/A sky130_fd_sc_hd__dfrtp_4
X_21315_ _21239_/X _21312_/X _12285_/B _21309_/X VGND VGND VPWR VPWR _21315_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14335__A1 _11977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22295_ _22139_/X _22293_/X _14790_/B _22290_/X VGND VGND VPWR VPWR _23331_/D sky130_fd_sc_hd__o22a_4
XANTENNA__16380__A _15959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24034_ _24066_/CLK _24034_/D VGND VGND VPWR VPWR _15352_/B sky130_fd_sc_hd__dfxtp_4
X_21246_ _21246_/A VGND VGND VPWR VPWR _21246_/X sky130_fd_sc_hd__buf_2
XFILLER_105_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13509__A _15884_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21081__B2 _21079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21177_ _20419_/X _21176_/X _23960_/Q _21173_/X VGND VGND VPWR VPWR _21177_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12413__A _12596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20128_ _20176_/A _20128_/B VGND VGND VPWR VPWR _20128_/X sky130_fd_sc_hd__or2_4
XFILLER_63_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21726__A _21690_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12132__B _12132_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12950_ _12974_/A _23987_/Q VGND VGND VPWR VPWR _12950_/X sky130_fd_sc_hd__or2_4
XANTENNA__15724__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20059_ _18531_/X _20057_/X _20058_/Y _20044_/X VGND VGND VPWR VPWR _20059_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21384__A2 _21383_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18785__B1 _24434_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11901_ _15952_/A VGND VGND VPWR VPWR _11901_/X sky130_fd_sc_hd__buf_2
X_12881_ _13951_/A VGND VGND VPWR VPWR _13960_/A sky130_fd_sc_hd__buf_2
XFILLER_46_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15443__B _23084_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13244__A _12367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ _11780_/X _23646_/Q VGND VGND VPWR VPWR _11833_/C sky130_fd_sc_hd__or2_4
X_14620_ _14756_/A _14620_/B VGND VGND VPWR VPWR _14620_/X sky130_fd_sc_hd__or2_4
X_23818_ _23564_/CLK _21432_/X VGND VGND VPWR VPWR _23818_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22557__A _22521_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21136__A2 _21133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14059__B _23690_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14519_/X _14487_/B VGND VGND VPWR VPWR _14551_/X sky130_fd_sc_hd__or2_4
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11675_/X _11736_/X _11763_/C VGND VGND VPWR VPWR _11763_/X sky130_fd_sc_hd__and3_4
X_23749_ _23973_/CLK _21566_/X VGND VGND VPWR VPWR _14506_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18001__A2 _17953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16555__A _12022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _15879_/A _13502_/B VGND VGND VPWR VPWR _13502_/X sky130_fd_sc_hd__or2_4
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _13025_/A _14482_/B _14482_/C VGND VGND VPWR VPWR _14482_/X sky130_fd_sc_hd__or3_4
X_17270_ _17267_/X _17270_/B VGND VGND VPWR VPWR _17270_/X sky130_fd_sc_hd__or2_4
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _14178_/A VGND VGND VPWR VPWR _13839_/A sky130_fd_sc_hd__buf_2
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20077__A _20090_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13433_ _11861_/X _13433_/B _13433_/C VGND VGND VPWR VPWR _13433_/X sky130_fd_sc_hd__or3_4
X_16221_ _16162_/X _16221_/B _16220_/X VGND VGND VPWR VPWR _16221_/X sky130_fd_sc_hd__and3_4
XANTENNA__11699__A _13256_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19386__A1_N _19374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14075__A _14074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16152_ _16152_/A _16147_/X _16151_/X VGND VGND VPWR VPWR _16153_/B sky130_fd_sc_hd__or3_4
X_13364_ _13352_/X _13291_/B VGND VGND VPWR VPWR _13364_/X sky130_fd_sc_hd__or2_4
X_12315_ _12315_/A VGND VGND VPWR VPWR _15693_/A sky130_fd_sc_hd__buf_2
X_15103_ _15110_/A _23775_/Q VGND VGND VPWR VPWR _15103_/X sky130_fd_sc_hd__or2_4
X_16083_ _16083_/A VGND VGND VPWR VPWR _16109_/A sky130_fd_sc_hd__buf_2
X_13295_ _12730_/A VGND VGND VPWR VPWR _13301_/A sky130_fd_sc_hd__buf_2
XANTENNA__14803__A _13862_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15034_ _13927_/A _24063_/Q VGND VGND VPWR VPWR _15035_/C sky130_fd_sc_hd__or2_4
X_19911_ _19909_/X _24152_/Q _19910_/X _20754_/A VGND VGND VPWR VPWR _24152_/D sky130_fd_sc_hd__o22a_4
XFILLER_108_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12246_ _12725_/A _12246_/B VGND VGND VPWR VPWR _12246_/X sky130_fd_sc_hd__or2_4
XFILLER_114_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15618__B _15556_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19842_ _21297_/A VGND VGND VPWR VPWR _21162_/C sky130_fd_sc_hd__buf_2
X_12177_ _11827_/A _12177_/B VGND VGND VPWR VPWR _12177_/X sky130_fd_sc_hd__or2_4
XFILLER_111_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12323__A _12738_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21636__A _21636_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19773_ _19722_/A _19742_/X _19592_/A VGND VGND VPWR VPWR _19773_/X sky130_fd_sc_hd__o21a_4
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16985_ _16985_/A _16984_/X VGND VGND VPWR VPWR _16985_/X sky130_fd_sc_hd__or2_4
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12042__B _23517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18724_ _18480_/X _18722_/X _18508_/X _18723_/X VGND VGND VPWR VPWR _18724_/X sky130_fd_sc_hd__o22a_4
XFILLER_77_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15936_ _15936_/A _15936_/B _15935_/X VGND VGND VPWR VPWR _15942_/B sky130_fd_sc_hd__and3_4
XFILLER_42_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17579__A1 _17132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21375__A2 _21369_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12977__B _23859_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18655_ _18498_/A _18655_/B VGND VGND VPWR VPWR _18655_/X sky130_fd_sc_hd__or2_4
X_15867_ _13546_/X _15798_/B VGND VGND VPWR VPWR _15867_/X sky130_fd_sc_hd__or2_4
XFILLER_58_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18945__A _19027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17606_ _18655_/B _17306_/A _17305_/A VGND VGND VPWR VPWR _17606_/X sky130_fd_sc_hd__o21a_4
XANTENNA__13154__A _12730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14818_ _14039_/A _14818_/B _14818_/C VGND VGND VPWR VPWR _14818_/X sky130_fd_sc_hd__or3_4
X_18586_ _17618_/C _18585_/B VGND VGND VPWR VPWR _18586_/X sky130_fd_sc_hd__or2_4
X_15798_ _12462_/A _15798_/B VGND VGND VPWR VPWR _15798_/X sky130_fd_sc_hd__or2_4
XFILLER_33_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18528__B1 _18523_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22467__A _22471_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17537_ _17144_/Y _17570_/A VGND VGND VPWR VPWR _17628_/A sky130_fd_sc_hd__or2_4
X_14749_ _13959_/A _23139_/Q VGND VGND VPWR VPWR _14751_/B sky130_fd_sc_hd__or2_4
XANTENNA__12993__A _12924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17468_ _17039_/A _17467_/X _17043_/A VGND VGND VPWR VPWR _17662_/B sky130_fd_sc_hd__o21a_4
X_19207_ _24258_/Q _19207_/B VGND VGND VPWR VPWR _19208_/B sky130_fd_sc_hd__and2_4
X_16419_ _16121_/A _16415_/X _16418_/X VGND VGND VPWR VPWR _16419_/X sky130_fd_sc_hd__or3_4
XFILLER_34_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22627__A2 _22622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19776__A _19775_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17399_ _17603_/B VGND VGND VPWR VPWR _17422_/B sky130_fd_sc_hd__buf_2
XANTENNA__18680__A _18679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20638__A1 _20613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19138_ _19138_/A _19137_/X VGND VGND VPWR VPWR _19138_/X sky130_fd_sc_hd__and2_4
XANTENNA__20638__B2 _20592_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19069_ _19052_/X _19067_/X _19068_/Y _19057_/X VGND VGND VPWR VPWR _19069_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15809__A _12886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21100_ _21079_/A VGND VGND VPWR VPWR _21100_/X sky130_fd_sc_hd__buf_2
XFILLER_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22080_ _22079_/X _22077_/X _16559_/B _22072_/X VGND VGND VPWR VPWR _23452_/D sky130_fd_sc_hd__o22a_4
XANTENNA__23872__CLK _23840_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21031_ _20537_/X _21030_/X _24051_/Q _21027_/X VGND VGND VPWR VPWR _21031_/X sky130_fd_sc_hd__o22a_4
XFILLER_102_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20271__C1 _20270_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22012__B1 _15253_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19016__A _19002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22982_ _22982_/A _22979_/Y _22981_/X VGND VGND VPWR VPWR _22982_/X sky130_fd_sc_hd__and3_4
XFILLER_83_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22563__B2 _22518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21933_ _21807_/X _21931_/X _23543_/Q _21928_/X VGND VGND VPWR VPWR _23543_/D sky130_fd_sc_hd__o22a_4
XFILLER_95_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13064__A _13104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21864_ _21863_/X _21817_/A _23583_/Q _21787_/X VGND VGND VPWR VPWR _23583_/D sky130_fd_sc_hd__o22a_4
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23603_ _23987_/CLK _21818_/X VGND VGND VPWR VPWR _23603_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23252__CLK _24047_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20815_ _24231_/Q _20639_/X _20814_/X VGND VGND VPWR VPWR _20815_/X sky130_fd_sc_hd__o21a_4
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13999__A _11645_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21795_ _21795_/A VGND VGND VPWR VPWR _21795_/X sky130_fd_sc_hd__buf_2
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16375__A _16374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23534_ _23692_/CLK _21946_/X VGND VGND VPWR VPWR _15670_/B sky130_fd_sc_hd__dfxtp_4
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20746_ _24202_/Q _20614_/X _20745_/Y VGND VGND VPWR VPWR _20747_/A sky130_fd_sc_hd__o21a_4
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23465_ _23910_/CLK _22053_/X VGND VGND VPWR VPWR _23465_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20677_ _20317_/B _20822_/B VGND VGND VPWR VPWR _20677_/X sky130_fd_sc_hd__or2_4
XANTENNA__12408__A _11671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22824__B _22824_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22416_ _22416_/A VGND VGND VPWR VPWR _22416_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23396_ _24066_/CLK _23396_/D VGND VGND VPWR VPWR _14620_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_13_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20625__A _20407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22347_ _22354_/A VGND VGND VPWR VPWR _22347_/X sky130_fd_sc_hd__buf_2
XFILLER_100_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15719__A _12765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14623__A _15036_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12100_ _16541_/A VGND VGND VPWR VPWR _12100_/X sky130_fd_sc_hd__buf_2
X_13080_ _13080_/A _23282_/Q VGND VGND VPWR VPWR _13081_/C sky130_fd_sc_hd__or2_4
X_22278_ _22110_/X _22272_/X _13502_/B _22276_/X VGND VGND VPWR VPWR _23343_/D sky130_fd_sc_hd__o22a_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12031_ _11837_/X _12031_/B VGND VGND VPWR VPWR _12034_/A sky130_fd_sc_hd__and2_4
X_24017_ _24082_/CLK _24017_/D VGND VGND VPWR VPWR _24017_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21229_ _21799_/A VGND VGND VPWR VPWR _21229_/X sky130_fd_sc_hd__buf_2
XANTENNA__21054__B2 _21048_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19798__A2 _19793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21456__A _21470_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17653__B _17653_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11982__A _11982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16770_ _16757_/X _16767_/X _16769_/X VGND VGND VPWR VPWR _16770_/X sky130_fd_sc_hd__and3_4
X_13982_ _13982_/A _13982_/B _13982_/C VGND VGND VPWR VPWR _13986_/B sky130_fd_sc_hd__and3_4
XANTENNA__14492__B1 _11596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15721_ _13129_/A _15659_/B VGND VGND VPWR VPWR _15721_/X sky130_fd_sc_hd__or2_4
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12933_ _12926_/A _12858_/B VGND VGND VPWR VPWR _12933_/X sky130_fd_sc_hd__or2_4
XANTENNA__15173__B _23617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18765__A _18781_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18440_ _18204_/A _17361_/X VGND VGND VPWR VPWR _18440_/X sky130_fd_sc_hd__or2_4
XFILLER_74_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15652_ _12221_/X _15652_/B VGND VGND VPWR VPWR _15652_/X sky130_fd_sc_hd__or2_4
X_12864_ _12518_/X _24019_/Q VGND VGND VPWR VPWR _12866_/B sky130_fd_sc_hd__or2_4
XFILLER_34_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21109__A2 _21075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14603_ _14603_/A _14601_/X _14602_/X VGND VGND VPWR VPWR _14603_/X sky130_fd_sc_hd__and3_4
X_11815_ _11730_/X _11815_/B _11814_/X VGND VGND VPWR VPWR _11815_/X sky130_fd_sc_hd__and3_4
X_18371_ _18107_/X _18367_/Y _18249_/X _18370_/Y VGND VGND VPWR VPWR _18371_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15901__B _15831_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12795_ _12795_/A VGND VGND VPWR VPWR _12803_/A sky130_fd_sc_hd__buf_2
X_15583_ _15614_/A _15522_/B VGND VGND VPWR VPWR _15585_/B sky130_fd_sc_hd__or2_4
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _15381_/X _17322_/B VGND VGND VPWR VPWR _17322_/X sky130_fd_sc_hd__or2_4
XFILLER_42_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _11745_/X VGND VGND VPWR VPWR _11746_/X sky130_fd_sc_hd__buf_2
X_14534_ _14556_/A _14532_/X _14534_/C VGND VGND VPWR VPWR _14534_/X sky130_fd_sc_hd__and3_4
XFILLER_57_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _17244_/X _17250_/X _17252_/X VGND VGND VPWR VPWR _17253_/X sky130_fd_sc_hd__o21a_4
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _13992_/A VGND VGND VPWR VPWR _14816_/A sky130_fd_sc_hd__buf_2
X_14465_ _12878_/A _14535_/B VGND VGND VPWR VPWR _14467_/B sky130_fd_sc_hd__or2_4
XANTENNA__22609__A2 _22607_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12318__A _12196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16204_ _16223_/A _23607_/Q VGND VGND VPWR VPWR _16206_/B sky130_fd_sc_hd__or2_4
X_13416_ _13395_/X _23472_/Q VGND VGND VPWR VPWR _13416_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_64_0_HCLK clkbuf_7_65_0_HCLK/A VGND VGND VPWR VPWR _24293_/CLK sky130_fd_sc_hd__clkbuf_1
X_14396_ _15607_/A _14393_/X _14396_/C VGND VGND VPWR VPWR _14397_/C sky130_fd_sc_hd__and3_4
X_17184_ _17130_/X _17180_/X _17163_/X _17183_/X VGND VGND VPWR VPWR _17184_/X sky130_fd_sc_hd__o22a_4
XFILLER_6_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21220__A2_N _21218_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13347_ _12682_/X _13346_/X VGND VGND VPWR VPWR _13347_/X sky130_fd_sc_hd__and2_4
X_16135_ _16139_/A _16135_/B VGND VGND VPWR VPWR _16136_/C sky130_fd_sc_hd__or2_4
X_13278_ _13272_/B VGND VGND VPWR VPWR _13278_/X sky130_fd_sc_hd__buf_2
X_16066_ _16058_/A _16066_/B _16065_/X VGND VGND VPWR VPWR _16066_/X sky130_fd_sc_hd__and3_4
XFILLER_68_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12229_ _12691_/A _12229_/B VGND VGND VPWR VPWR _12230_/C sky130_fd_sc_hd__or2_4
X_15017_ _13957_/A _15017_/B VGND VGND VPWR VPWR _15017_/X sky130_fd_sc_hd__and2_4
XANTENNA__13149__A _15667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21045__B2 _21041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23125__CLK _23699_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19825_ _19449_/X _19672_/D _19822_/Y _21112_/A _19490_/X VGND VGND VPWR VPWR _24169_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21366__A _21373_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12988__A _12392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19756_ _19661_/A _19631_/Y _19689_/A VGND VGND VPWR VPWR _19789_/B sky130_fd_sc_hd__or3_4
X_16968_ _18558_/A _18557_/A VGND VGND VPWR VPWR _16969_/B sky130_fd_sc_hd__or2_4
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18707_ _18704_/Y _18706_/X _18704_/Y _18706_/X VGND VGND VPWR VPWR _19356_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22545__B2 _22540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15919_ _15919_/A VGND VGND VPWR VPWR _15919_/Y sky130_fd_sc_hd__inv_2
X_19687_ _19873_/B _19867_/C VGND VGND VPWR VPWR _19687_/X sky130_fd_sc_hd__or2_4
XANTENNA__19410__B2 _24193_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16899_ _16899_/A _16899_/B VGND VGND VPWR VPWR _16899_/X sky130_fd_sc_hd__or2_4
XFILLER_65_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18638_ _18638_/A VGND VGND VPWR VPWR _18638_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17972__B2 _17805_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18569_ _18568_/X VGND VGND VPWR VPWR _18569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16195__A _16219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14708__A _15592_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20600_ _20468_/X _20599_/Y _19220_/A _20562_/X VGND VGND VPWR VPWR _20600_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13612__A _13800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21580_ _23742_/Q VGND VGND VPWR VPWR _21580_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22925__A _23048_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20531_ _20531_/A VGND VGND VPWR VPWR _20531_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12228__A _12221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23250_ _23314_/CLK _22419_/X VGND VGND VPWR VPWR _13064_/B sky130_fd_sc_hd__dfxtp_4
X_20462_ _24214_/Q _20398_/X _20461_/Y VGND VGND VPWR VPWR _20463_/A sky130_fd_sc_hd__o21a_4
XFILLER_53_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20445__A _20342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22201_ _21112_/B _21348_/C _21634_/D VGND VGND VPWR VPWR _22201_/X sky130_fd_sc_hd__or3_4
XFILLER_10_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16642__B _23548_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17488__B1 _17021_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21284__A1 _21282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23181_ _23564_/CLK _23181_/D VGND VGND VPWR VPWR _15852_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_88_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21284__B2 _21278_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22481__B1 _16226_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20393_ _20393_/A VGND VGND VPWR VPWR _21802_/A sky130_fd_sc_hd__buf_2
XFILLER_88_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22132_ _22108_/A VGND VGND VPWR VPWR _22132_/X sky130_fd_sc_hd__buf_2
XFILLER_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18472__A1_N _17261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22063_ _21859_/X _22059_/X _15240_/B _22020_/X VGND VGND VPWR VPWR _22063_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21036__B2 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21014_ _21004_/Y _21013_/X _20277_/X _21013_/X VGND VGND VPWR VPWR _21014_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12898__A _12520_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15274__A _14165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21339__A2 _21333_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22965_ _22955_/X _17699_/X _22937_/X _22964_/X VGND VGND VPWR VPWR _22966_/A sky130_fd_sc_hd__a211o_4
XFILLER_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19401__B2 _24200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21916_ _21296_/A VGND VGND VPWR VPWR _21917_/B sky130_fd_sc_hd__buf_2
XFILLER_55_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22896_ _19901_/X _24112_/Q _18701_/X _18679_/X _22889_/X VGND VGND VPWR VPWR _22896_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_3_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16817__B _16816_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21847_ _20838_/A VGND VGND VPWR VPWR _21847_/X sky130_fd_sc_hd__buf_2
XFILLER_110_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15721__B _15659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14618__A _12439_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _17533_/A _17543_/A _17552_/A VGND VGND VPWR VPWR _11601_/A sky130_fd_sc_hd__or3_4
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13522__A _13522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12980_/A _12580_/B VGND VGND VPWR VPWR _12580_/X sky130_fd_sc_hd__or2_4
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21778_ _21570_/X _21776_/X _14773_/B _21773_/X VGND VGND VPWR VPWR _23619_/D sky130_fd_sc_hd__o22a_4
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21511__A2 _21508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _24346_/Q _11530_/X VGND VGND VPWR VPWR _11531_/X sky130_fd_sc_hd__or2_4
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20729_ _20642_/X _20727_/X _20728_/X VGND VGND VPWR VPWR _20729_/X sky130_fd_sc_hd__and3_4
X_23517_ _23514_/CLK _23517_/D VGND VGND VPWR VPWR _23517_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _13686_/A _14250_/B _14249_/X VGND VGND VPWR VPWR _14259_/B sky130_fd_sc_hd__or3_4
XANTENNA__18751__C _18751_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23448_ _23383_/CLK _22090_/X VGND VGND VPWR VPWR _15969_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13201__A1 _12716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20355__A _20355_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _12716_/X _13177_/X _13184_/X _13192_/X _13200_/X VGND VGND VPWR VPWR _13201_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16552__B _23548_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11977__A _15420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20078__A2 _18600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14181_ _11708_/A VGND VGND VPWR VPWR _14182_/A sky130_fd_sc_hd__buf_2
XANTENNA__15449__A _15449_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23379_ _23311_/CLK _22223_/X VGND VGND VPWR VPWR _23379_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_99_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23148__CLK _23564_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14353__A _14345_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13132_ _13082_/A _13132_/B _13131_/X VGND VGND VPWR VPWR _13133_/C sky130_fd_sc_hd__or3_4
XFILLER_98_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13063_ _15480_/A VGND VGND VPWR VPWR _13104_/A sky130_fd_sc_hd__buf_2
X_17940_ _17858_/X VGND VGND VPWR VPWR _18327_/A sky130_fd_sc_hd__buf_2
XFILLER_97_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12014_ _12008_/A _12014_/B VGND VGND VPWR VPWR _12016_/B sky130_fd_sc_hd__or2_4
XFILLER_105_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23298__CLK _23812_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17871_ _17871_/A _17871_/B VGND VGND VPWR VPWR _17871_/X sky130_fd_sc_hd__and2_4
Xclkbuf_4_6_0_HCLK clkbuf_4_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19610_ _19607_/X _19862_/A _19578_/X _19609_/X VGND VGND VPWR VPWR _19610_/X sky130_fd_sc_hd__a211o_4
XFILLER_117_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16822_ _12188_/Y _16819_/X _12188_/Y _16819_/X VGND VGND VPWR VPWR _16822_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12601__A _12646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19541_ _19541_/A _19541_/B VGND VGND VPWR VPWR _19582_/A sky130_fd_sc_hd__or2_4
X_16753_ _16598_/X _16746_/X _16752_/X VGND VGND VPWR VPWR _16753_/X sky130_fd_sc_hd__or3_4
X_13965_ _12302_/A _13961_/X _13965_/C VGND VGND VPWR VPWR _13965_/X sky130_fd_sc_hd__or3_4
XFILLER_24_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18495__A _17422_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15704_ _12743_/A _15763_/B VGND VGND VPWR VPWR _15705_/C sky130_fd_sc_hd__or2_4
XANTENNA__15912__A _15910_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20002__A2 _19985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12916_ _13009_/A _12974_/B VGND VGND VPWR VPWR _12916_/X sky130_fd_sc_hd__or2_4
X_19472_ _19468_/X _19754_/A VGND VGND VPWR VPWR _19526_/B sky130_fd_sc_hd__or2_4
XFILLER_74_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16684_ _16583_/A _23515_/Q VGND VGND VPWR VPWR _16685_/C sky130_fd_sc_hd__or2_4
X_13896_ _13896_/A _13896_/B _13895_/X VGND VGND VPWR VPWR _13896_/X sky130_fd_sc_hd__and3_4
XFILLER_74_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21750__A2 _21748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18423_ _18422_/X VGND VGND VPWR VPWR _18423_/Y sky130_fd_sc_hd__inv_2
X_15635_ _13884_/A _15635_/B _15635_/C VGND VGND VPWR VPWR _15643_/B sky130_fd_sc_hd__or3_4
X_12847_ _12443_/A _12925_/B VGND VGND VPWR VPWR _12849_/B sky130_fd_sc_hd__or2_4
XFILLER_22_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14528__A _13711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13432__A _11913_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18354_ _18354_/A _18354_/B VGND VGND VPWR VPWR _18354_/X sky130_fd_sc_hd__and2_4
X_15566_ _14431_/A _23467_/Q VGND VGND VPWR VPWR _15566_/X sky130_fd_sc_hd__or2_4
X_12778_ _12777_/X VGND VGND VPWR VPWR _12813_/A sky130_fd_sc_hd__buf_2
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17305_/A VGND VGND VPWR VPWR _17305_/Y sky130_fd_sc_hd__inv_2
X_14517_ _14556_/A _14515_/X _14517_/C VGND VGND VPWR VPWR _14517_/X sky130_fd_sc_hd__and3_4
XFILLER_30_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11729_ _16048_/A VGND VGND VPWR VPWR _11729_/X sky130_fd_sc_hd__buf_2
X_18285_ _17758_/X _17759_/X _18285_/C VGND VGND VPWR VPWR _18285_/X sky130_fd_sc_hd__or3_4
X_15497_ _15497_/A _23404_/Q VGND VGND VPWR VPWR _15497_/X sky130_fd_sc_hd__or2_4
XFILLER_30_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17236_ _17863_/A _17216_/X _17845_/A _17235_/X VGND VGND VPWR VPWR _17236_/X sky130_fd_sc_hd__o22a_4
X_14448_ _12862_/A _14446_/X _14447_/X VGND VGND VPWR VPWR _14448_/X sky130_fd_sc_hd__and3_4
XFILLER_80_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15359__A _14810_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11887__A _11886_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17167_ _17130_/X _17162_/X _17163_/X _17166_/X VGND VGND VPWR VPWR _17167_/X sky130_fd_sc_hd__o22a_4
X_14379_ _14379_/A _14379_/B VGND VGND VPWR VPWR _14380_/C sky130_fd_sc_hd__or2_4
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16118_ _16145_/A _16186_/B VGND VGND VPWR VPWR _16118_/X sky130_fd_sc_hd__or2_4
XFILLER_31_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17098_ _17063_/A VGND VGND VPWR VPWR _17173_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17574__A _16374_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21018__B2 _21013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16049_ _16037_/A _23608_/Q VGND VGND VPWR VPWR _16051_/B sky130_fd_sc_hd__or2_4
XFILLER_44_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21569__A2 _21568_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21096__A _21067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19808_ _19808_/A _19718_/B VGND VGND VPWR VPWR _19808_/X sky130_fd_sc_hd__or2_4
XFILLER_84_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12511__A _13623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21824__A _21812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19739_ _19670_/X VGND VGND VPWR VPWR _19740_/A sky130_fd_sc_hd__buf_2
XFILLER_38_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22750_ _22750_/A _22747_/X VGND VGND VPWR VPWR _22750_/X sky130_fd_sc_hd__and2_4
XFILLER_65_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15822__A _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21701_ _21524_/X _21698_/X _12246_/B _21695_/X VGND VGND VPWR VPWR _23670_/D sky130_fd_sc_hd__o22a_4
XANTENNA__17945__B2 _17944_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22681_ _20442_/A _22679_/X _23095_/Q _22676_/X VGND VGND VPWR VPWR _23095_/D sky130_fd_sc_hd__o22a_4
XANTENNA__14438__A _12533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24420_ _24425_/CLK _24420_/D HRESETn VGND VGND VPWR VPWR _24420_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13342__A _12740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21632_ _21578_/X _21605_/A _23711_/Q _21595_/A VGND VGND VPWR VPWR _23711_/D sky130_fd_sc_hd__o22a_4
XFILLER_55_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24351_ _24425_/CLK _24351_/D HRESETn VGND VGND VPWR VPWR _24351_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_90_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21563_ _21527_/A VGND VGND VPWR VPWR _21563_/X sky130_fd_sc_hd__buf_2
XANTENNA__16653__A _16622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23302_ _23845_/CLK _22324_/X VGND VGND VPWR VPWR _14287_/B sky130_fd_sc_hd__dfxtp_4
X_20514_ _20422_/X _20895_/B _20286_/X VGND VGND VPWR VPWR _20514_/X sky130_fd_sc_hd__a21o_4
X_24282_ _24344_/CLK _24282_/D HRESETn VGND VGND VPWR VPWR _19231_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_53_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15184__A1 _12267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21494_ _21287_/X _21491_/X _15304_/B _21488_/X VGND VGND VPWR VPWR _23778_/D sky130_fd_sc_hd__o22a_4
XFILLER_88_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23233_ _23233_/CLK _22459_/X VGND VGND VPWR VPWR _15125_/B sky130_fd_sc_hd__dfxtp_4
X_20445_ _20342_/A _20445_/B VGND VGND VPWR VPWR _20445_/X sky130_fd_sc_hd__and2_4
XFILLER_10_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15269__A _14158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21257__B2 _21254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23164_ _23324_/CLK _23164_/D VGND VGND VPWR VPWR _16631_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20376_ _20212_/X VGND VGND VPWR VPWR _20376_/X sky130_fd_sc_hd__buf_2
XANTENNA__19683__B _19754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22390__A _20314_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22115_ _20670_/A VGND VGND VPWR VPWR _22115_/X sky130_fd_sc_hd__buf_2
X_23095_ _23699_/CLK _23095_/D VGND VGND VPWR VPWR _23095_/Q sky130_fd_sc_hd__dfxtp_4
X_22046_ _21828_/X _22045_/X _15769_/B _22042_/X VGND VGND VPWR VPWR _23470_/D sky130_fd_sc_hd__o22a_4
XFILLER_47_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13517__A _13507_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12421__A _12421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22509__B2 _22504_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21980__A2 _21974_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23997_ _24026_/CLK _21120_/X VGND VGND VPWR VPWR _23997_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12140__B _12140_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15732__A _12792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13750_ _13699_/A _13750_/B _13749_/X VGND VGND VPWR VPWR _13750_/X sky130_fd_sc_hd__and3_4
XFILLER_44_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19204__A _20190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22948_ _22948_/A VGND VGND VPWR VPWR HADDR[11] sky130_fd_sc_hd__inv_2
XFILLER_43_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21732__A2 _21705_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16547__B _23996_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12701_ _12722_/A _23988_/Q VGND VGND VPWR VPWR _12702_/C sky130_fd_sc_hd__or2_4
XFILLER_56_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13681_ _15449_/A _13681_/B _13681_/C VGND VGND VPWR VPWR _13682_/B sky130_fd_sc_hd__or3_4
X_22879_ _19893_/X _22821_/X _15713_/Y _22855_/A VGND VGND VPWR VPWR _22879_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_70_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15420_ _15420_/A _15419_/X VGND VGND VPWR VPWR _15420_/X sky130_fd_sc_hd__and2_4
XANTENNA__13252__A _15484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12632_ _12660_/A _23317_/Q VGND VGND VPWR VPWR _12632_/X sky130_fd_sc_hd__or2_4
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12563_ _13738_/A VGND VGND VPWR VPWR _12655_/A sky130_fd_sc_hd__buf_2
X_15351_ _15332_/A _15285_/B VGND VGND VPWR VPWR _15351_/X sky130_fd_sc_hd__or2_4
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21496__B2 _21452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ _24329_/Q _11514_/B VGND VGND VPWR VPWR _11515_/B sky130_fd_sc_hd__or2_4
X_14302_ _12260_/X _14302_/B VGND VGND VPWR VPWR _14303_/C sky130_fd_sc_hd__or2_4
XFILLER_106_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18070_ _17824_/X _17832_/Y _17921_/A _17840_/Y VGND VGND VPWR VPWR _18070_/X sky130_fd_sc_hd__o22a_4
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _12494_/A VGND VGND VPWR VPWR _12920_/A sky130_fd_sc_hd__buf_2
X_15282_ _15142_/A _15282_/B VGND VGND VPWR VPWR _15282_/X sky130_fd_sc_hd__or2_4
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16282__B _16282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17021_ _17021_/A VGND VGND VPWR VPWR _17022_/A sky130_fd_sc_hd__buf_2
X_14233_ _14201_/A _14233_/B _14232_/X VGND VGND VPWR VPWR _14243_/B sky130_fd_sc_hd__or3_4
XANTENNA__15179__A _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21248__B2 _21242_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14164_ _14992_/A _23081_/Q VGND VGND VPWR VPWR _14166_/B sky130_fd_sc_hd__or2_4
X_13115_ _13115_/A _13039_/B VGND VGND VPWR VPWR _13116_/C sky130_fd_sc_hd__or2_4
XANTENNA__24136__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14095_ _15011_/A VGND VGND VPWR VPWR _14990_/A sky130_fd_sc_hd__buf_2
X_18972_ _11528_/A VGND VGND VPWR VPWR _18972_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15907__A _11657_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13046_ _13046_/A _13046_/B VGND VGND VPWR VPWR _13046_/X sky130_fd_sc_hd__or2_4
X_17923_ _17910_/X _17919_/Y _17921_/X _17922_/Y VGND VGND VPWR VPWR _17923_/X sky130_fd_sc_hd__o22a_4
XFILLER_80_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17854_ _18249_/A VGND VGND VPWR VPWR _17854_/X sky130_fd_sc_hd__buf_2
XANTENNA__21420__B2 _21416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12331__A _12745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16805_ _16747_/X _16805_/B _16805_/C VGND VGND VPWR VPWR _16809_/B sky130_fd_sc_hd__and3_4
X_17785_ _18206_/A _17785_/B VGND VGND VPWR VPWR _17789_/C sky130_fd_sc_hd__and2_4
X_14997_ _14997_/A _23743_/Q VGND VGND VPWR VPWR _14998_/C sky130_fd_sc_hd__or2_4
XANTENNA__16738__A _11997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19524_ _19481_/A _19524_/B VGND VGND VPWR VPWR _19686_/A sky130_fd_sc_hd__or2_4
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16736_ _11875_/X _16736_/B _16736_/C VGND VGND VPWR VPWR _16740_/B sky130_fd_sc_hd__and3_4
X_13948_ _13972_/A _13944_/X _13948_/C VGND VGND VPWR VPWR _13948_/X sky130_fd_sc_hd__or3_4
Xclkbuf_1_1_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_1_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19455_ _24157_/Q _19435_/X _20224_/B _19432_/X VGND VGND VPWR VPWR _19455_/X sky130_fd_sc_hd__o22a_4
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16667_ _16640_/X _16665_/X _16666_/X VGND VGND VPWR VPWR _16667_/X sky130_fd_sc_hd__and3_4
X_13879_ _13879_/A _13792_/B VGND VGND VPWR VPWR _13879_/X sky130_fd_sc_hd__or2_4
XANTENNA__14258__A _14367_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18406_ _18405_/A _18404_/X _18160_/X VGND VGND VPWR VPWR _18406_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__13162__A _12710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15618_ _15618_/A _15556_/B VGND VGND VPWR VPWR _15619_/C sky130_fd_sc_hd__or2_4
X_19386_ _19374_/X _18238_/X _19385_/X _24211_/Q VGND VGND VPWR VPWR _24211_/D sky130_fd_sc_hd__a2bb2o_4
X_16598_ _11685_/X VGND VGND VPWR VPWR _16598_/X sky130_fd_sc_hd__buf_2
XFILLER_50_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18337_ _17758_/X _18336_/X _17758_/X _18336_/X VGND VGND VPWR VPWR _18337_/X sky130_fd_sc_hd__a2bb2o_4
X_15549_ _12459_/A _15545_/X _15548_/X VGND VGND VPWR VPWR _15549_/X sky130_fd_sc_hd__or3_4
XANTENNA__21487__B2 _21481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24378__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18268_ _18268_/A VGND VGND VPWR VPWR _18268_/Y sky130_fd_sc_hd__inv_2
X_17219_ _17141_/X _17217_/X _17154_/X _17218_/X VGND VGND VPWR VPWR _17219_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22436__B1 _15522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18199_ _24130_/Q _18174_/B _16982_/X VGND VGND VPWR VPWR _18199_/X sky130_fd_sc_hd__o21a_4
XFILLER_102_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_34_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_34_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12506__A _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12924__B1 _11596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20230_ _18759_/A _20224_/B _20229_/X VGND VGND VPWR VPWR _20230_/X sky130_fd_sc_hd__a21o_4
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21819__A _21249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20161_ _24438_/Q IRQ[23] _20160_/X VGND VGND VPWR VPWR _20161_/Y sky130_fd_sc_hd__a21boi_4
X_20092_ _20076_/X _20091_/Y _11628_/X _18604_/X _18649_/X VGND VGND VPWR VPWR _20092_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_83_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15536__B _23659_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23920_ _23920_/CLK _23920_/D VGND VGND VPWR VPWR _13308_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13337__A _13428_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21411__B2 _21409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12241__A _12240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21962__A2 _21959_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13056__B _13055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23851_ _24044_/CLK _23851_/D VGND VGND VPWR VPWR _15577_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22802_ _13685_/Y _22794_/X _22796_/X _22801_/X VGND VGND VPWR VPWR _22803_/B sky130_fd_sc_hd__o22a_4
XFILLER_2_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15552__A _15552_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19024__A _18994_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19907__A2 _24154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20994_ _20493_/A _20993_/X _19108_/B _20500_/A VGND VGND VPWR VPWR _20994_/X sky130_fd_sc_hd__o22a_4
X_23782_ _23781_/CLK _21489_/X VGND VGND VPWR VPWR _14328_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_96_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21714__A2 _21712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16367__B _16289_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22733_ SYSTICKCLKDIV[3] VGND VGND VPWR VPWR _22733_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17394__A2 _17340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14168__A _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22664_ _23102_/Q VGND VGND VPWR VPWR _22664_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22385__A _22384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21066__A2_N _21065_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21615_ _21548_/X _21612_/X _15459_/B _21609_/X VGND VGND VPWR VPWR _21615_/X sky130_fd_sc_hd__o22a_4
X_24403_ _23326_/CLK _24403_/D HRESETn VGND VGND VPWR VPWR _20519_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_116_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR _24084_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__21478__B2 _21474_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22595_ _22430_/X _22593_/X _15863_/B _22590_/X VGND VGND VPWR VPWR _22595_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16383__A _15999_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13800__A _13800_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21546_ _21831_/A VGND VGND VPWR VPWR _21546_/X sky130_fd_sc_hd__buf_2
X_24334_ _24334_/CLK _19029_/X HRESETn VGND VGND VPWR VPWR _11519_/A sky130_fd_sc_hd__dfstp_4
XFILLER_33_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24265_ _24305_/CLK _19278_/X HRESETn VGND VGND VPWR VPWR _24265_/Q sky130_fd_sc_hd__dfrtp_4
X_21477_ _21470_/A VGND VGND VPWR VPWR _21477_/X sky130_fd_sc_hd__buf_2
XFILLER_14_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12416__A _12413_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23216_ _23473_/CLK _23216_/D VGND VGND VPWR VPWR _13336_/B sky130_fd_sc_hd__dfxtp_4
X_20428_ _20427_/Y _20258_/X VGND VGND VPWR VPWR _20428_/X sky130_fd_sc_hd__or2_4
X_24196_ _24199_/CLK _24196_/D HRESETn VGND VGND VPWR VPWR _24196_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18646__A2 _18641_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23147_ _23336_/CLK _22598_/X VGND VGND VPWR VPWR _23147_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20359_ _20229_/X _20358_/X _20213_/X VGND VGND VPWR VPWR _20359_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21650__B2 _21645_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14631__A _15006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23078_ _23781_/CLK _23078_/D VGND VGND VPWR VPWR _14327_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_103_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14920_ _11646_/A _14856_/B VGND VGND VPWR VPWR _14922_/B sky130_fd_sc_hd__or2_4
X_22029_ _21799_/X _22024_/X _16427_/B _22028_/X VGND VGND VPWR VPWR _23482_/D sky130_fd_sc_hd__o22a_4
XFILLER_76_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12151__A _16045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21953__A2 _21952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14851_ _14851_/A VGND VGND VPWR VPWR _14851_/X sky130_fd_sc_hd__buf_2
XANTENNA__17661__B _17459_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11990__A _11982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13802_ _13641_/A _13875_/B VGND VGND VPWR VPWR _13803_/C sky130_fd_sc_hd__or2_4
XFILLER_29_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17570_ _17570_/A VGND VGND VPWR VPWR _17570_/Y sky130_fd_sc_hd__inv_2
X_14782_ _14782_/A _14778_/X _14782_/C VGND VGND VPWR VPWR _14783_/B sky130_fd_sc_hd__or3_4
XFILLER_99_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11994_ _11994_/A _21161_/A VGND VGND VPWR VPWR _11995_/C sky130_fd_sc_hd__or2_4
XFILLER_99_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16521_ _16081_/A _16237_/Y _16080_/A VGND VGND VPWR VPWR _16521_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_72_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13733_ _15494_/A _13630_/B VGND VGND VPWR VPWR _13733_/X sky130_fd_sc_hd__or2_4
XFILLER_95_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14078__A _12202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19240_ _24284_/Q _19233_/B _19239_/Y VGND VGND VPWR VPWR _24284_/D sky130_fd_sc_hd__o21a_4
X_16452_ _16465_/A _16384_/B VGND VGND VPWR VPWR _16453_/C sky130_fd_sc_hd__or2_4
X_13664_ _15432_/A _13664_/B VGND VGND VPWR VPWR _13666_/B sky130_fd_sc_hd__or2_4
XANTENNA__19588__B HRDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15403_ _13623_/A _15403_/B VGND VGND VPWR VPWR _15404_/C sky130_fd_sc_hd__or2_4
X_12615_ _12643_/A _12505_/B VGND VGND VPWR VPWR _12615_/X sky130_fd_sc_hd__or2_4
X_19171_ _19124_/B VGND VGND VPWR VPWR _19171_/Y sky130_fd_sc_hd__inv_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17389__A _13918_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21469__B2 _21467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16383_ _15999_/X _16383_/B VGND VGND VPWR VPWR _16383_/X sky130_fd_sc_hd__or2_4
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ _13595_/A VGND VGND VPWR VPWR _13595_/X sky130_fd_sc_hd__buf_2
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16293__A _11884_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14806__A _14845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22130__A2 _22125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18122_ _17568_/Y _18121_/X VGND VGND VPWR VPWR _18122_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__13710__A _13710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15334_ _15334_/A _15332_/X _15334_/C VGND VGND VPWR VPWR _15338_/B sky130_fd_sc_hd__and3_4
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24388__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12546_ _12546_/A _12667_/B VGND VGND VPWR VPWR _12546_/X sky130_fd_sc_hd__or2_4
XFILLER_8_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18053_ _18224_/A VGND VGND VPWR VPWR _18053_/X sky130_fd_sc_hd__buf_2
XANTENNA__24317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15265_ _14136_/A _15265_/B _15264_/X VGND VGND VPWR VPWR _15265_/X sky130_fd_sc_hd__or3_4
XFILLER_32_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12477_ _13029_/A VGND VGND VPWR VPWR _12477_/X sky130_fd_sc_hd__buf_2
XANTENNA__12326__A _13317_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17004_ _16993_/X _17003_/A _16937_/X _17003_/Y VGND VGND VPWR VPWR _17004_/X sky130_fd_sc_hd__o22a_4
X_14216_ _13709_/A VGND VGND VPWR VPWR _14345_/A sky130_fd_sc_hd__buf_2
X_15196_ _15201_/A _15196_/B VGND VGND VPWR VPWR _15196_/X sky130_fd_sc_hd__or2_4
XANTENNA__19834__A1 _19775_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14147_ _15010_/A VGND VGND VPWR VPWR _15026_/A sky130_fd_sc_hd__buf_2
XFILLER_99_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14078_ _12202_/A _14078_/B VGND VGND VPWR VPWR _14081_/B sky130_fd_sc_hd__or2_4
X_18955_ _18941_/X _18953_/Y _18954_/Y _18946_/X VGND VGND VPWR VPWR _18955_/X sky130_fd_sc_hd__o22a_4
XFILLER_45_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22197__A2 _22193_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13157__A _15696_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13029_ _13029_/A _23954_/Q VGND VGND VPWR VPWR _13030_/C sky130_fd_sc_hd__or2_4
X_17906_ _17801_/X _17167_/X _17807_/X _17147_/X VGND VGND VPWR VPWR _17906_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18886_ _16374_/X _18884_/X _18961_/A _18885_/X VGND VGND VPWR VPWR _24377_/D sky130_fd_sc_hd__o22a_4
XANTENNA__21944__A2 _21938_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17837_ _17837_/A VGND VGND VPWR VPWR _17837_/X sky130_fd_sc_hd__buf_2
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16468__A _16159_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17768_ _17767_/X VGND VGND VPWR VPWR _17768_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16719_ _16542_/A _16719_/B _16719_/C VGND VGND VPWR VPWR _16719_/X sky130_fd_sc_hd__or3_4
X_19507_ _19718_/A VGND VGND VPWR VPWR _19877_/B sky130_fd_sc_hd__buf_2
XANTENNA__15091__B _15023_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17699_ _17699_/A VGND VGND VPWR VPWR _17699_/X sky130_fd_sc_hd__buf_2
XANTENNA__17376__A2 _17013_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19438_ _19462_/A VGND VGND VPWR VPWR _19438_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19369_ _19367_/X _17898_/X _19367_/X _24219_/Q VGND VGND VPWR VPWR _24219_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21400_ _21400_/A VGND VGND VPWR VPWR _21416_/A sky130_fd_sc_hd__inv_2
XANTENNA__22121__A2 _22113_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13620__A _13620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22380_ _22145_/X _22375_/X _14868_/B _22344_/A VGND VGND VPWR VPWR _23264_/D sky130_fd_sc_hd__o22a_4
XANTENNA__22933__A _18548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21331_ _21265_/X _21326_/X _23883_/Q _21330_/X VGND VGND VPWR VPWR _21331_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12236__A _12693_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16931__A _17062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24050_ _23986_/CLK _24050_/D VGND VGND VPWR VPWR _24050_/Q sky130_fd_sc_hd__dfxtp_4
X_21262_ _21261_/X _21259_/X _15805_/B _21254_/X VGND VGND VPWR VPWR _23917_/D sky130_fd_sc_hd__o22a_4
XFILLER_116_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23209__CLK _23433_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20453__A _20453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23001_ _22985_/X _17667_/A _22997_/X _23000_/X VGND VGND VPWR VPWR _23001_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16650__B _23612_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20213_ _20212_/X VGND VGND VPWR VPWR _20213_/X sky130_fd_sc_hd__buf_2
XFILLER_89_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21193_ _20697_/X _21190_/X _15487_/B _21187_/X VGND VGND VPWR VPWR _23948_/D sky130_fd_sc_hd__o22a_4
XFILLER_46_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21632__B2 _21595_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14451__A _12494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20144_ IRQ[9] VGND VGND VPWR VPWR _20144_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15311__A1 _12267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22188__A2 _22186_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20075_ NMI _20074_/Y VGND VGND VPWR VPWR _20076_/B sky130_fd_sc_hd__or2_4
XANTENNA__21396__B1 _23839_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20900__B _20556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23903_ _23217_/CLK _21294_/X VGND VGND VPWR VPWR _23903_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23834_ _23706_/CLK _23834_/D VGND VGND VPWR VPWR _16421_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_22_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19689__A _19689_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20977_ _20616_/X _20964_/X _20757_/X _20976_/Y VGND VGND VPWR VPWR _20977_/X sky130_fd_sc_hd__a211o_4
X_23765_ _24021_/CLK _21528_/X VGND VGND VPWR VPWR _12463_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__21699__B2 _21695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22896__B1 _18679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22360__A2 _22354_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22716_ _22932_/A _22723_/B VGND VGND VPWR VPWR _23064_/C sky130_fd_sc_hd__and2_4
XFILLER_0_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23696_ _23157_/CLK _23696_/D VGND VGND VPWR VPWR _23696_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23004__A _18222_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22648__B1 _23115_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22647_ _22633_/A VGND VGND VPWR VPWR _22647_/X sky130_fd_sc_hd__buf_2
XFILLER_9_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12400_ _12826_/A _12293_/B VGND VGND VPWR VPWR _12402_/B sky130_fd_sc_hd__or2_4
X_13380_ _13399_/A _13377_/X _13380_/C VGND VGND VPWR VPWR _13380_/X sky130_fd_sc_hd__and3_4
XFILLER_22_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22578_ _22401_/X _22572_/X _16266_/B _22576_/X VGND VGND VPWR VPWR _23161_/D sky130_fd_sc_hd__o22a_4
XFILLER_70_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24361__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12331_ _12745_/A _12331_/B VGND VGND VPWR VPWR _12331_/X sky130_fd_sc_hd__or2_4
X_24317_ _24290_/CLK _24317_/D HRESETn VGND VGND VPWR VPWR _19138_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21529_ _20509_/A VGND VGND VPWR VPWR _21529_/X sky130_fd_sc_hd__buf_2
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12262_ _12743_/A VGND VGND VPWR VPWR _15667_/A sky130_fd_sc_hd__buf_2
X_15050_ _15050_/A VGND VGND VPWR VPWR _15050_/Y sky130_fd_sc_hd__inv_2
X_24248_ _24216_/CLK _24248_/D HRESETn VGND VGND VPWR VPWR _20414_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19816__B2 _19531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14001_ _14021_/A _23338_/Q VGND VGND VPWR VPWR _14001_/X sky130_fd_sc_hd__or2_4
XFILLER_68_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12193_ _13055_/A VGND VGND VPWR VPWR _12556_/A sky130_fd_sc_hd__buf_2
X_24179_ _23584_/CLK _19717_/X HRESETn VGND VGND VPWR VPWR _11905_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_64_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20082__B _20071_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15176__B _15176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18768__A _18782_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18740_ _17084_/A VGND VGND VPWR VPWR _18750_/B sky130_fd_sc_hd__inv_2
XANTENNA__17672__A _17672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15952_ _15952_/A _15952_/B VGND VGND VPWR VPWR _15952_/X sky130_fd_sc_hd__or2_4
XFILLER_89_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21926__A2 _21924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14903_ _14906_/A _14903_/B VGND VGND VPWR VPWR _14903_/X sky130_fd_sc_hd__or2_4
XANTENNA__21194__A _21180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18671_ _17324_/X _18670_/Y VGND VGND VPWR VPWR _18671_/X sky130_fd_sc_hd__or2_4
XFILLER_37_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15883_ _15876_/A _15821_/B VGND VGND VPWR VPWR _15883_/X sky130_fd_sc_hd__or2_4
X_17622_ _17595_/X _17622_/B VGND VGND VPWR VPWR _17622_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14834_ _14841_/A _14776_/B VGND VGND VPWR VPWR _14834_/X sky130_fd_sc_hd__or2_4
XANTENNA__13705__A _13754_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17553_ _17039_/A _17552_/X _17043_/A VGND VGND VPWR VPWR _17652_/B sky130_fd_sc_hd__o21a_4
X_14765_ _13606_/A _14765_/B VGND VGND VPWR VPWR _14765_/X sky130_fd_sc_hd__or2_4
X_11977_ _15420_/A VGND VGND VPWR VPWR _11977_/X sky130_fd_sc_hd__buf_2
X_16504_ _16471_/X _16427_/B VGND VGND VPWR VPWR _16504_/X sky130_fd_sc_hd__or2_4
X_13716_ _12578_/A VGND VGND VPWR VPWR _15493_/A sky130_fd_sc_hd__buf_2
XFILLER_75_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17484_ _17484_/A _17483_/X VGND VGND VPWR VPWR _18274_/A sky130_fd_sc_hd__or2_4
X_14696_ _14672_/A _14696_/B VGND VGND VPWR VPWR _14697_/C sky130_fd_sc_hd__or2_4
XFILLER_32_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19223_ _19223_/A _19261_/A VGND VGND VPWR VPWR _19223_/X sky130_fd_sc_hd__and2_4
XANTENNA__16735__B _23803_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16435_ _16100_/X _16435_/B VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__or2_4
X_13647_ _13647_/A _13647_/B _13646_/X VGND VGND VPWR VPWR _13648_/B sky130_fd_sc_hd__or3_4
XFILLER_32_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13440__A _13467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19154_ _19132_/A _19132_/B _19153_/Y VGND VGND VPWR VPWR _24311_/D sky130_fd_sc_hd__o21a_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16366_ _16366_/A _16366_/B _16366_/C VGND VGND VPWR VPWR _16366_/X sky130_fd_sc_hd__and3_4
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _13578_/A VGND VGND VPWR VPWR _13578_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21311__B1 _16272_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18105_ _18180_/A _18100_/Y _18105_/C _18105_/D VGND VGND VPWR VPWR _18106_/A sky130_fd_sc_hd__or4_4
X_15317_ _13871_/A _15255_/B VGND VGND VPWR VPWR _15317_/X sky130_fd_sc_hd__or2_4
XANTENNA__24151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12529_ _12529_/A VGND VGND VPWR VPWR _15032_/A sky130_fd_sc_hd__buf_2
X_19085_ _18965_/A _19082_/Y _19083_/Y _19084_/X VGND VGND VPWR VPWR _19085_/X sky130_fd_sc_hd__o22a_4
XFILLER_118_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16297_ _15956_/A _16297_/B VGND VGND VPWR VPWR _16298_/C sky130_fd_sc_hd__or2_4
XFILLER_69_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12056__A _11943_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21862__B2 _21787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18036_ _17244_/X _17215_/Y _17921_/A _17234_/Y VGND VGND VPWR VPWR _18036_/X sky130_fd_sc_hd__o22a_4
X_15248_ _11798_/A _15232_/X _15248_/C VGND VGND VPWR VPWR _15248_/X sky130_fd_sc_hd__or3_4
XANTENNA__21369__A _21369_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11895__A _15393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15367__A _12567_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21614__B2 _21609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15179_ _15026_/A _23681_/Q VGND VGND VPWR VPWR _15181_/B sky130_fd_sc_hd__or2_4
XFILLER_113_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14271__A _12257_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21090__A2 _21089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19987_ _18091_/X _19985_/X _19986_/Y _19972_/X VGND VGND VPWR VPWR _19987_/X sky130_fd_sc_hd__o22a_4
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18938_ _11533_/X VGND VGND VPWR VPWR _19027_/A sky130_fd_sc_hd__buf_2
.ends

