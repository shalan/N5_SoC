VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NfiVe32_SYS
  CLASS BLOCK ;
  FOREIGN NfiVe32_SYS ;
  ORIGIN 0.000 0.000 ;
  SIZE 794.740 BY 349.510 ;
  PIN HADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.760 0.000 55.040 4.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.280 0.000 60.560 4.000 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.340 0.000 65.620 4.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.860 0.000 71.140 4.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.380 0.000 76.660 4.000 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.900 0.000 82.180 4.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.420 0.000 87.700 4.000 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.940 0.000 93.220 4.000 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.460 0.000 98.740 4.000 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.980 0.000 104.260 4.000 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.080 0.000 5.360 4.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.500 0.000 109.780 4.000 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.020 0.000 115.300 4.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.540 0.000 120.820 4.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.600 0.000 125.880 4.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.120 0.000 131.400 4.000 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.640 0.000 136.920 4.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.160 0.000 142.440 4.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.680 0.000 147.960 4.000 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.200 0.000 153.480 4.000 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.720 0.000 159.000 4.000 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.600 0.000 10.880 4.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.240 0.000 164.520 4.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.760 0.000 170.040 4.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.120 0.000 16.400 4.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.640 0.000 21.920 4.000 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.160 0.000 27.440 4.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.680 0.000 32.960 4.000 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.200 0.000 38.480 4.000 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.720 0.000 44.000 4.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.240 0.000 49.520 4.000 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.500 0.000 569.780 4.000 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.280 0.000 175.560 4.000 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.020 0.000 230.300 4.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.540 0.000 235.820 4.000 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.060 0.000 241.340 4.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.120 0.000 246.400 4.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.640 0.000 251.920 4.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.160 0.000 257.440 4.000 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.680 0.000 262.960 4.000 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.200 0.000 268.480 4.000 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.720 0.000 274.000 4.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.240 0.000 279.520 4.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.800 0.000 181.080 4.000 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.760 0.000 285.040 4.000 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.280 0.000 290.560 4.000 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.800 0.000 296.080 4.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.320 0.000 301.600 4.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.840 0.000 307.120 4.000 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.900 0.000 312.180 4.000 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.420 0.000 317.700 4.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.940 0.000 323.220 4.000 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.460 0.000 328.740 4.000 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.980 0.000 334.260 4.000 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.860 0.000 186.140 4.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.500 0.000 339.780 4.000 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.020 0.000 345.300 4.000 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.380 0.000 191.660 4.000 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.900 0.000 197.180 4.000 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.420 0.000 202.700 4.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.940 0.000 208.220 4.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.460 0.000 213.740 4.000 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.980 0.000 219.260 4.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.500 0.000 224.780 4.000 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.060 0.000 586.340 4.000 ;
    END
  END HREADY
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.020 0.000 575.300 4.000 ;
    END
  END HRESETn
  PIN HSIZE[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.100 0.000 597.380 4.000 ;
    END
  END HSIZE[0]
  PIN HSIZE[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.620 0.000 602.900 4.000 ;
    END
  END HSIZE[1]
  PIN HSIZE[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.140 0.000 608.420 4.000 ;
    END
  END HSIZE[2]
  PIN HTRANS[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.660 0.000 613.940 4.000 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.720 0.000 619.000 4.000 ;
    END
  END HTRANS[1]
  PIN HWDATA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.540 0.000 350.820 4.000 ;
    END
  END HWDATA[0]
  PIN HWDATA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.280 0.000 405.560 4.000 ;
    END
  END HWDATA[10]
  PIN HWDATA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.800 0.000 411.080 4.000 ;
    END
  END HWDATA[11]
  PIN HWDATA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.320 0.000 416.600 4.000 ;
    END
  END HWDATA[12]
  PIN HWDATA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.840 0.000 422.120 4.000 ;
    END
  END HWDATA[13]
  PIN HWDATA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.360 0.000 427.640 4.000 ;
    END
  END HWDATA[14]
  PIN HWDATA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.420 0.000 432.700 4.000 ;
    END
  END HWDATA[15]
  PIN HWDATA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.940 0.000 438.220 4.000 ;
    END
  END HWDATA[16]
  PIN HWDATA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.460 0.000 443.740 4.000 ;
    END
  END HWDATA[17]
  PIN HWDATA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.980 0.000 449.260 4.000 ;
    END
  END HWDATA[18]
  PIN HWDATA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.500 0.000 454.780 4.000 ;
    END
  END HWDATA[19]
  PIN HWDATA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.060 0.000 356.340 4.000 ;
    END
  END HWDATA[1]
  PIN HWDATA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.020 0.000 460.300 4.000 ;
    END
  END HWDATA[20]
  PIN HWDATA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.540 0.000 465.820 4.000 ;
    END
  END HWDATA[21]
  PIN HWDATA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.060 0.000 471.340 4.000 ;
    END
  END HWDATA[22]
  PIN HWDATA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.580 0.000 476.860 4.000 ;
    END
  END HWDATA[23]
  PIN HWDATA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.100 0.000 482.380 4.000 ;
    END
  END HWDATA[24]
  PIN HWDATA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.620 0.000 487.900 4.000 ;
    END
  END HWDATA[25]
  PIN HWDATA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.680 0.000 492.960 4.000 ;
    END
  END HWDATA[26]
  PIN HWDATA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.200 0.000 498.480 4.000 ;
    END
  END HWDATA[27]
  PIN HWDATA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.720 0.000 504.000 4.000 ;
    END
  END HWDATA[28]
  PIN HWDATA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.240 0.000 509.520 4.000 ;
    END
  END HWDATA[29]
  PIN HWDATA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.580 0.000 361.860 4.000 ;
    END
  END HWDATA[2]
  PIN HWDATA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.760 0.000 515.040 4.000 ;
    END
  END HWDATA[30]
  PIN HWDATA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.280 0.000 520.560 4.000 ;
    END
  END HWDATA[31]
  PIN HWDATA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.100 0.000 367.380 4.000 ;
    END
  END HWDATA[3]
  PIN HWDATA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.160 0.000 372.440 4.000 ;
    END
  END HWDATA[4]
  PIN HWDATA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.680 0.000 377.960 4.000 ;
    END
  END HWDATA[5]
  PIN HWDATA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.200 0.000 383.480 4.000 ;
    END
  END HWDATA[6]
  PIN HWDATA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.720 0.000 389.000 4.000 ;
    END
  END HWDATA[7]
  PIN HWDATA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.240 0.000 394.520 4.000 ;
    END
  END HWDATA[8]
  PIN HWDATA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.760 0.000 400.040 4.000 ;
    END
  END HWDATA[9]
  PIN HWRITE
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.540 0.000 580.820 4.000 ;
    END
  END HWRITE
  PIN IRQ[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.240 0.000 624.520 4.000 ;
    END
  END IRQ[0]
  PIN IRQ[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.980 0.000 679.260 4.000 ;
    END
  END IRQ[10]
  PIN IRQ[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.500 0.000 684.780 4.000 ;
    END
  END IRQ[11]
  PIN IRQ[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.020 0.000 690.300 4.000 ;
    END
  END IRQ[12]
  PIN IRQ[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.540 0.000 695.820 4.000 ;
    END
  END IRQ[13]
  PIN IRQ[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.060 0.000 701.340 4.000 ;
    END
  END IRQ[14]
  PIN IRQ[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.580 0.000 706.860 4.000 ;
    END
  END IRQ[15]
  PIN IRQ[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.100 0.000 712.380 4.000 ;
    END
  END IRQ[16]
  PIN IRQ[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.620 0.000 717.900 4.000 ;
    END
  END IRQ[17]
  PIN IRQ[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.140 0.000 723.420 4.000 ;
    END
  END IRQ[18]
  PIN IRQ[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.660 0.000 728.940 4.000 ;
    END
  END IRQ[19]
  PIN IRQ[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.760 0.000 630.040 4.000 ;
    END
  END IRQ[1]
  PIN IRQ[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.180 0.000 734.460 4.000 ;
    END
  END IRQ[20]
  PIN IRQ[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.240 0.000 739.520 4.000 ;
    END
  END IRQ[21]
  PIN IRQ[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.760 0.000 745.040 4.000 ;
    END
  END IRQ[22]
  PIN IRQ[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.280 0.000 750.560 4.000 ;
    END
  END IRQ[23]
  PIN IRQ[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.800 0.000 756.080 4.000 ;
    END
  END IRQ[24]
  PIN IRQ[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.320 0.000 761.600 4.000 ;
    END
  END IRQ[25]
  PIN IRQ[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.840 0.000 767.120 4.000 ;
    END
  END IRQ[26]
  PIN IRQ[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.360 0.000 772.640 4.000 ;
    END
  END IRQ[27]
  PIN IRQ[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.880 0.000 778.160 4.000 ;
    END
  END IRQ[28]
  PIN IRQ[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.400 0.000 783.680 4.000 ;
    END
  END IRQ[29]
  PIN IRQ[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.280 0.000 635.560 4.000 ;
    END
  END IRQ[2]
  PIN IRQ[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.920 0.000 789.200 4.000 ;
    END
  END IRQ[30]
  PIN IRQ[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.440 0.000 794.720 4.000 ;
    END
  END IRQ[31]
  PIN IRQ[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.800 0.000 641.080 4.000 ;
    END
  END IRQ[3]
  PIN IRQ[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.320 0.000 646.600 4.000 ;
    END
  END IRQ[4]
  PIN IRQ[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.840 0.000 652.120 4.000 ;
    END
  END IRQ[5]
  PIN IRQ[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.360 0.000 657.640 4.000 ;
    END
  END IRQ[6]
  PIN IRQ[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.880 0.000 663.160 4.000 ;
    END
  END IRQ[7]
  PIN IRQ[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.400 0.000 668.680 4.000 ;
    END
  END IRQ[8]
  PIN IRQ[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.920 0.000 674.200 4.000 ;
    END
  END IRQ[9]
  PIN NMI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.580 0.000 591.860 4.000 ;
    END
  END NMI
  PIN SYSTICKCLKDIV[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.800 0.000 526.080 4.000 ;
    END
  END SYSTICKCLKDIV[0]
  PIN SYSTICKCLKDIV[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.320 0.000 531.600 4.000 ;
    END
  END SYSTICKCLKDIV[1]
  PIN SYSTICKCLKDIV[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.840 0.000 537.120 4.000 ;
    END
  END SYSTICKCLKDIV[2]
  PIN SYSTICKCLKDIV[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.360 0.000 542.640 4.000 ;
    END
  END SYSTICKCLKDIV[3]
  PIN SYSTICKCLKDIV[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.880 0.000 548.160 4.000 ;
    END
  END SYSTICKCLKDIV[4]
  PIN SYSTICKCLKDIV[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.400 0.000 553.680 4.000 ;
    END
  END SYSTICKCLKDIV[5]
  PIN SYSTICKCLKDIV[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.460 0.000 558.740 4.000 ;
    END
  END SYSTICKCLKDIV[6]
  PIN SYSTICKCLKDIV[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.980 0.000 564.260 4.000 ;
    END
  END SYSTICKCLKDIV[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 786.670 10.640 788.270 337.520 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 633.070 10.640 634.670 337.520 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 479.470 10.640 481.070 337.520 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 325.870 10.640 327.470 337.520 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 172.270 10.640 173.870 337.520 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.670 10.640 20.270 337.520 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 709.870 10.640 711.470 337.520 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 556.270 10.640 557.870 337.520 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 402.670 10.640 404.270 337.520 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 249.070 10.640 250.670 337.520 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.470 10.640 97.070 337.520 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 3.150 7.225 792.050 342.635 ;
      LAYER met1 ;
        RECT 0.000 0.040 794.740 349.480 ;
      LAYER met2 ;
        RECT 0.030 4.280 794.710 349.510 ;
        RECT 0.580 0.010 4.800 4.280 ;
        RECT 5.640 0.010 10.320 4.280 ;
        RECT 11.160 0.010 15.840 4.280 ;
        RECT 16.680 0.010 21.360 4.280 ;
        RECT 22.200 0.010 26.880 4.280 ;
        RECT 27.720 0.010 32.400 4.280 ;
        RECT 33.240 0.010 37.920 4.280 ;
        RECT 38.760 0.010 43.440 4.280 ;
        RECT 44.280 0.010 48.960 4.280 ;
        RECT 49.800 0.010 54.480 4.280 ;
        RECT 55.320 0.010 60.000 4.280 ;
        RECT 60.840 0.010 65.060 4.280 ;
        RECT 65.900 0.010 70.580 4.280 ;
        RECT 71.420 0.010 76.100 4.280 ;
        RECT 76.940 0.010 81.620 4.280 ;
        RECT 82.460 0.010 87.140 4.280 ;
        RECT 87.980 0.010 92.660 4.280 ;
        RECT 93.500 0.010 98.180 4.280 ;
        RECT 99.020 0.010 103.700 4.280 ;
        RECT 104.540 0.010 109.220 4.280 ;
        RECT 110.060 0.010 114.740 4.280 ;
        RECT 115.580 0.010 120.260 4.280 ;
        RECT 121.100 0.010 125.320 4.280 ;
        RECT 126.160 0.010 130.840 4.280 ;
        RECT 131.680 0.010 136.360 4.280 ;
        RECT 137.200 0.010 141.880 4.280 ;
        RECT 142.720 0.010 147.400 4.280 ;
        RECT 148.240 0.010 152.920 4.280 ;
        RECT 153.760 0.010 158.440 4.280 ;
        RECT 159.280 0.010 163.960 4.280 ;
        RECT 164.800 0.010 169.480 4.280 ;
        RECT 170.320 0.010 175.000 4.280 ;
        RECT 175.840 0.010 180.520 4.280 ;
        RECT 181.360 0.010 185.580 4.280 ;
        RECT 186.420 0.010 191.100 4.280 ;
        RECT 191.940 0.010 196.620 4.280 ;
        RECT 197.460 0.010 202.140 4.280 ;
        RECT 202.980 0.010 207.660 4.280 ;
        RECT 208.500 0.010 213.180 4.280 ;
        RECT 214.020 0.010 218.700 4.280 ;
        RECT 219.540 0.010 224.220 4.280 ;
        RECT 225.060 0.010 229.740 4.280 ;
        RECT 230.580 0.010 235.260 4.280 ;
        RECT 236.100 0.010 240.780 4.280 ;
        RECT 241.620 0.010 245.840 4.280 ;
        RECT 246.680 0.010 251.360 4.280 ;
        RECT 252.200 0.010 256.880 4.280 ;
        RECT 257.720 0.010 262.400 4.280 ;
        RECT 263.240 0.010 267.920 4.280 ;
        RECT 268.760 0.010 273.440 4.280 ;
        RECT 274.280 0.010 278.960 4.280 ;
        RECT 279.800 0.010 284.480 4.280 ;
        RECT 285.320 0.010 290.000 4.280 ;
        RECT 290.840 0.010 295.520 4.280 ;
        RECT 296.360 0.010 301.040 4.280 ;
        RECT 301.880 0.010 306.560 4.280 ;
        RECT 307.400 0.010 311.620 4.280 ;
        RECT 312.460 0.010 317.140 4.280 ;
        RECT 317.980 0.010 322.660 4.280 ;
        RECT 323.500 0.010 328.180 4.280 ;
        RECT 329.020 0.010 333.700 4.280 ;
        RECT 334.540 0.010 339.220 4.280 ;
        RECT 340.060 0.010 344.740 4.280 ;
        RECT 345.580 0.010 350.260 4.280 ;
        RECT 351.100 0.010 355.780 4.280 ;
        RECT 356.620 0.010 361.300 4.280 ;
        RECT 362.140 0.010 366.820 4.280 ;
        RECT 367.660 0.010 371.880 4.280 ;
        RECT 372.720 0.010 377.400 4.280 ;
        RECT 378.240 0.010 382.920 4.280 ;
        RECT 383.760 0.010 388.440 4.280 ;
        RECT 389.280 0.010 393.960 4.280 ;
        RECT 394.800 0.010 399.480 4.280 ;
        RECT 400.320 0.010 405.000 4.280 ;
        RECT 405.840 0.010 410.520 4.280 ;
        RECT 411.360 0.010 416.040 4.280 ;
        RECT 416.880 0.010 421.560 4.280 ;
        RECT 422.400 0.010 427.080 4.280 ;
        RECT 427.920 0.010 432.140 4.280 ;
        RECT 432.980 0.010 437.660 4.280 ;
        RECT 438.500 0.010 443.180 4.280 ;
        RECT 444.020 0.010 448.700 4.280 ;
        RECT 449.540 0.010 454.220 4.280 ;
        RECT 455.060 0.010 459.740 4.280 ;
        RECT 460.580 0.010 465.260 4.280 ;
        RECT 466.100 0.010 470.780 4.280 ;
        RECT 471.620 0.010 476.300 4.280 ;
        RECT 477.140 0.010 481.820 4.280 ;
        RECT 482.660 0.010 487.340 4.280 ;
        RECT 488.180 0.010 492.400 4.280 ;
        RECT 493.240 0.010 497.920 4.280 ;
        RECT 498.760 0.010 503.440 4.280 ;
        RECT 504.280 0.010 508.960 4.280 ;
        RECT 509.800 0.010 514.480 4.280 ;
        RECT 515.320 0.010 520.000 4.280 ;
        RECT 520.840 0.010 525.520 4.280 ;
        RECT 526.360 0.010 531.040 4.280 ;
        RECT 531.880 0.010 536.560 4.280 ;
        RECT 537.400 0.010 542.080 4.280 ;
        RECT 542.920 0.010 547.600 4.280 ;
        RECT 548.440 0.010 553.120 4.280 ;
        RECT 553.960 0.010 558.180 4.280 ;
        RECT 559.020 0.010 563.700 4.280 ;
        RECT 564.540 0.010 569.220 4.280 ;
        RECT 570.060 0.010 574.740 4.280 ;
        RECT 575.580 0.010 580.260 4.280 ;
        RECT 581.100 0.010 585.780 4.280 ;
        RECT 586.620 0.010 591.300 4.280 ;
        RECT 592.140 0.010 596.820 4.280 ;
        RECT 597.660 0.010 602.340 4.280 ;
        RECT 603.180 0.010 607.860 4.280 ;
        RECT 608.700 0.010 613.380 4.280 ;
        RECT 614.220 0.010 618.440 4.280 ;
        RECT 619.280 0.010 623.960 4.280 ;
        RECT 624.800 0.010 629.480 4.280 ;
        RECT 630.320 0.010 635.000 4.280 ;
        RECT 635.840 0.010 640.520 4.280 ;
        RECT 641.360 0.010 646.040 4.280 ;
        RECT 646.880 0.010 651.560 4.280 ;
        RECT 652.400 0.010 657.080 4.280 ;
        RECT 657.920 0.010 662.600 4.280 ;
        RECT 663.440 0.010 668.120 4.280 ;
        RECT 668.960 0.010 673.640 4.280 ;
        RECT 674.480 0.010 678.700 4.280 ;
        RECT 679.540 0.010 684.220 4.280 ;
        RECT 685.060 0.010 689.740 4.280 ;
        RECT 690.580 0.010 695.260 4.280 ;
        RECT 696.100 0.010 700.780 4.280 ;
        RECT 701.620 0.010 706.300 4.280 ;
        RECT 707.140 0.010 711.820 4.280 ;
        RECT 712.660 0.010 717.340 4.280 ;
        RECT 718.180 0.010 722.860 4.280 ;
        RECT 723.700 0.010 728.380 4.280 ;
        RECT 729.220 0.010 733.900 4.280 ;
        RECT 734.740 0.010 738.960 4.280 ;
        RECT 739.800 0.010 744.480 4.280 ;
        RECT 745.320 0.010 750.000 4.280 ;
        RECT 750.840 0.010 755.520 4.280 ;
        RECT 756.360 0.010 761.040 4.280 ;
        RECT 761.880 0.010 766.560 4.280 ;
        RECT 767.400 0.010 772.080 4.280 ;
        RECT 772.920 0.010 777.600 4.280 ;
        RECT 778.440 0.010 783.120 4.280 ;
        RECT 783.960 0.010 788.640 4.280 ;
        RECT 789.480 0.010 794.160 4.280 ;
      LAYER met3 ;
        RECT 6.895 1.535 788.270 344.580 ;
      LAYER met4 ;
        RECT 82.565 337.920 765.535 344.585 ;
        RECT 82.565 10.240 95.070 337.920 ;
        RECT 97.470 10.240 171.870 337.920 ;
        RECT 174.270 10.240 248.670 337.920 ;
        RECT 251.070 10.240 325.470 337.920 ;
        RECT 327.870 10.240 402.270 337.920 ;
        RECT 404.670 10.240 479.070 337.920 ;
        RECT 481.470 10.240 555.870 337.920 ;
        RECT 558.270 10.240 632.670 337.920 ;
        RECT 635.070 10.240 709.470 337.920 ;
        RECT 711.870 10.240 765.535 337.920 ;
        RECT 82.565 2.215 765.535 10.240 ;
  END
END NfiVe32_SYS
END LIBRARY

