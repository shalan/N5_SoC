VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM_4K
  CLASS BLOCK ;
  FOREIGN DFFRAM_4K ;
  ORIGIN 0.000 0.000 ;
  SIZE 1239.805 BY 1289.790 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.680 1285.790 501.960 1289.790 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.320 1285.790 517.600 1289.790 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.960 1285.790 533.240 1289.790 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.600 1285.790 548.880 1289.790 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.240 1285.790 564.520 1289.790 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.880 1285.790 580.160 1289.790 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.520 1285.790 595.800 1289.790 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.160 1285.790 611.440 1289.790 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.800 1285.790 627.080 1289.790 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.440 1285.790 642.720 1289.790 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.080 1285.790 658.360 1289.790 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.920 1285.790 752.200 1289.790 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.860 1285.790 908.140 1289.790 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.500 1285.790 923.780 1289.790 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.140 1285.790 939.420 1289.790 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.780 1285.790 955.060 1289.790 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.420 1285.790 970.700 1289.790 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.060 1285.790 986.340 1289.790 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.700 1285.790 1001.980 1289.790 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.340 1285.790 1017.620 1289.790 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.980 1285.790 1033.260 1289.790 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.620 1285.790 1048.900 1289.790 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.560 1285.790 767.840 1289.790 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.260 1285.790 1064.540 1289.790 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.900 1285.790 1080.180 1289.790 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.540 1285.790 1095.820 1289.790 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.180 1285.790 1111.460 1289.790 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.820 1285.790 1127.100 1289.790 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.460 1285.790 1142.740 1289.790 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.100 1285.790 1158.380 1289.790 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.740 1285.790 1174.020 1289.790 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.380 1285.790 1189.660 1289.790 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.020 1285.790 1205.300 1289.790 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.200 1285.790 783.480 1289.790 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.660 1285.790 1220.940 1289.790 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.300 1285.790 1236.580 1289.790 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.840 1285.790 799.120 1289.790 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.480 1285.790 814.760 1289.790 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.120 1285.790 830.400 1289.790 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.300 1285.790 845.580 1289.790 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.940 1285.790 861.220 1289.790 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.580 1285.790 876.860 1289.790 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.220 1285.790 892.500 1289.790 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.120 1285.790 2.400 1289.790 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.060 1285.790 158.340 1289.790 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.700 1285.790 173.980 1289.790 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.340 1285.790 189.620 1289.790 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.980 1285.790 205.260 1289.790 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.620 1285.790 220.900 1289.790 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.260 1285.790 236.540 1289.790 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.900 1285.790 252.180 1289.790 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.540 1285.790 267.820 1289.790 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.180 1285.790 283.460 1289.790 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.820 1285.790 299.100 1289.790 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.300 1285.790 17.580 1289.790 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.460 1285.790 314.740 1289.790 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.100 1285.790 330.380 1289.790 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.740 1285.790 346.020 1289.790 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.380 1285.790 361.660 1289.790 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.020 1285.790 377.300 1289.790 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.660 1285.790 392.940 1289.790 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.300 1285.790 408.580 1289.790 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.480 1285.790 423.760 1289.790 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.120 1285.790 439.400 1289.790 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.760 1285.790 455.040 1289.790 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.940 1285.790 33.220 1289.790 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.400 1285.790 470.680 1289.790 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.040 1285.790 486.320 1289.790 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.580 1285.790 48.860 1289.790 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.220 1285.790 64.500 1289.790 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.860 1285.790 80.140 1289.790 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.500 1285.790 95.780 1289.790 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.140 1285.790 111.420 1289.790 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.780 1285.790 127.060 1289.790 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.420 1285.790 142.700 1289.790 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.280 1285.790 736.560 1289.790 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.720 1285.790 674.000 1289.790 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.360 1285.790 689.640 1289.790 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.000 1285.790 705.280 1289.790 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.640 1285.790 720.920 1289.790 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1215.710 0.430 1217.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1095.710 0.430 1097.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 975.710 0.430 977.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 855.710 0.430 857.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 735.710 0.430 737.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 615.710 0.430 617.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 495.710 0.430 497.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 375.710 0.430 377.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 255.710 0.430 257.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 135.710 0.430 137.310 1276.590 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 0.430 17.310 1276.590 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1155.710 0.430 1157.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1035.710 0.430 1037.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 915.710 0.430 917.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 795.710 0.430 797.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 675.710 0.430 677.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 555.710 0.430 557.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 435.710 0.430 437.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 315.710 0.430 317.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 195.710 0.430 197.310 1276.590 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 75.710 0.430 77.310 1276.590 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 0.585 1239.745 1276.435 ;
      LAYER met1 ;
        RECT 0.190 0.030 1239.805 1280.050 ;
      LAYER met2 ;
        RECT 1.670 1285.510 1.840 1285.790 ;
        RECT 2.680 1285.510 17.020 1285.790 ;
        RECT 17.860 1285.510 32.660 1285.790 ;
        RECT 33.500 1285.510 48.300 1285.790 ;
        RECT 49.140 1285.510 63.940 1285.790 ;
        RECT 64.780 1285.510 79.580 1285.790 ;
        RECT 80.420 1285.510 95.220 1285.790 ;
        RECT 96.060 1285.510 110.860 1285.790 ;
        RECT 111.700 1285.510 126.500 1285.790 ;
        RECT 127.340 1285.510 142.140 1285.790 ;
        RECT 142.980 1285.510 157.780 1285.790 ;
        RECT 158.620 1285.510 173.420 1285.790 ;
        RECT 174.260 1285.510 189.060 1285.790 ;
        RECT 189.900 1285.510 204.700 1285.790 ;
        RECT 205.540 1285.510 220.340 1285.790 ;
        RECT 221.180 1285.510 235.980 1285.790 ;
        RECT 236.820 1285.510 251.620 1285.790 ;
        RECT 252.460 1285.510 267.260 1285.790 ;
        RECT 268.100 1285.510 282.900 1285.790 ;
        RECT 283.740 1285.510 298.540 1285.790 ;
        RECT 299.380 1285.510 314.180 1285.790 ;
        RECT 315.020 1285.510 329.820 1285.790 ;
        RECT 330.660 1285.510 345.460 1285.790 ;
        RECT 346.300 1285.510 361.100 1285.790 ;
        RECT 361.940 1285.510 376.740 1285.790 ;
        RECT 377.580 1285.510 392.380 1285.790 ;
        RECT 393.220 1285.510 408.020 1285.790 ;
        RECT 408.860 1285.510 423.200 1285.790 ;
        RECT 424.040 1285.510 438.840 1285.790 ;
        RECT 439.680 1285.510 454.480 1285.790 ;
        RECT 455.320 1285.510 470.120 1285.790 ;
        RECT 470.960 1285.510 485.760 1285.790 ;
        RECT 486.600 1285.510 501.400 1285.790 ;
        RECT 502.240 1285.510 517.040 1285.790 ;
        RECT 517.880 1285.510 532.680 1285.790 ;
        RECT 533.520 1285.510 548.320 1285.790 ;
        RECT 549.160 1285.510 563.960 1285.790 ;
        RECT 564.800 1285.510 579.600 1285.790 ;
        RECT 580.440 1285.510 595.240 1285.790 ;
        RECT 596.080 1285.510 610.880 1285.790 ;
        RECT 611.720 1285.510 626.520 1285.790 ;
        RECT 627.360 1285.510 642.160 1285.790 ;
        RECT 643.000 1285.510 657.800 1285.790 ;
        RECT 658.640 1285.510 673.440 1285.790 ;
        RECT 674.280 1285.510 689.080 1285.790 ;
        RECT 689.920 1285.510 704.720 1285.790 ;
        RECT 705.560 1285.510 720.360 1285.790 ;
        RECT 721.200 1285.510 736.000 1285.790 ;
        RECT 736.840 1285.510 751.640 1285.790 ;
        RECT 752.480 1285.510 767.280 1285.790 ;
        RECT 768.120 1285.510 782.920 1285.790 ;
        RECT 783.760 1285.510 798.560 1285.790 ;
        RECT 799.400 1285.510 814.200 1285.790 ;
        RECT 815.040 1285.510 829.840 1285.790 ;
        RECT 830.680 1285.510 845.020 1285.790 ;
        RECT 845.860 1285.510 860.660 1285.790 ;
        RECT 861.500 1285.510 876.300 1285.790 ;
        RECT 877.140 1285.510 891.940 1285.790 ;
        RECT 892.780 1285.510 907.580 1285.790 ;
        RECT 908.420 1285.510 923.220 1285.790 ;
        RECT 924.060 1285.510 938.860 1285.790 ;
        RECT 939.700 1285.510 954.500 1285.790 ;
        RECT 955.340 1285.510 970.140 1285.790 ;
        RECT 970.980 1285.510 985.780 1285.790 ;
        RECT 986.620 1285.510 1001.420 1285.790 ;
        RECT 1002.260 1285.510 1017.060 1285.790 ;
        RECT 1017.900 1285.510 1032.700 1285.790 ;
        RECT 1033.540 1285.510 1048.340 1285.790 ;
        RECT 1049.180 1285.510 1063.980 1285.790 ;
        RECT 1064.820 1285.510 1079.620 1285.790 ;
        RECT 1080.460 1285.510 1095.260 1285.790 ;
        RECT 1096.100 1285.510 1110.900 1285.790 ;
        RECT 1111.740 1285.510 1126.540 1285.790 ;
        RECT 1127.380 1285.510 1142.180 1285.790 ;
        RECT 1143.020 1285.510 1157.820 1285.790 ;
        RECT 1158.660 1285.510 1173.460 1285.790 ;
        RECT 1174.300 1285.510 1189.100 1285.790 ;
        RECT 1189.940 1285.510 1204.740 1285.790 ;
        RECT 1205.580 1285.510 1220.380 1285.790 ;
        RECT 1221.220 1285.510 1236.020 1285.790 ;
        RECT 1236.860 1285.510 1237.490 1285.790 ;
        RECT 1.670 0.000 1237.490 1285.510 ;
      LAYER met3 ;
        RECT 4.855 0.505 1236.605 1276.515 ;
      LAYER met4 ;
        RECT 36.365 89.925 75.310 1273.455 ;
        RECT 77.710 89.925 135.310 1273.455 ;
        RECT 137.710 89.925 195.310 1273.455 ;
        RECT 197.710 89.925 255.310 1273.455 ;
        RECT 257.710 89.925 315.310 1273.455 ;
        RECT 317.710 89.925 375.310 1273.455 ;
        RECT 377.710 89.925 435.310 1273.455 ;
        RECT 437.710 89.925 495.310 1273.455 ;
        RECT 497.710 89.925 555.310 1273.455 ;
        RECT 557.710 89.925 615.310 1273.455 ;
        RECT 617.710 89.925 675.310 1273.455 ;
        RECT 677.710 89.925 735.310 1273.455 ;
        RECT 737.710 89.925 795.310 1273.455 ;
        RECT 797.710 89.925 855.310 1273.455 ;
        RECT 857.710 89.925 915.310 1273.455 ;
        RECT 917.710 89.925 975.310 1273.455 ;
        RECT 977.710 89.925 1035.310 1273.455 ;
        RECT 1037.710 89.925 1095.310 1273.455 ;
        RECT 1097.710 89.925 1155.310 1273.455 ;
        RECT 1157.710 89.925 1215.310 1273.455 ;
        RECT 1217.710 89.925 1218.895 1273.455 ;
        RECT 0.300 0.300 1258.680 1295.880 ;
  END
END DFFRAM_4K
END LIBRARY

