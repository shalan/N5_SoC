VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO apb_sys_0
  CLASS BLOCK ;
  FOREIGN apb_sys_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 398.265 ;
  PIN HADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 0.000 700.000 0.600 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 33.320 700.000 33.920 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 36.720 700.000 37.320 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 40.120 700.000 40.720 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 43.520 700.000 44.120 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 46.920 700.000 47.520 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 50.320 700.000 50.920 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 53.720 700.000 54.320 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 57.120 700.000 57.720 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 59.840 700.000 60.440 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 63.240 700.000 63.840 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2.720 700.000 3.320 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 66.640 700.000 67.240 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 70.040 700.000 70.640 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 73.440 700.000 74.040 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 76.840 700.000 77.440 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 80.240 700.000 80.840 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 83.640 700.000 84.240 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 87.040 700.000 87.640 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 90.440 700.000 91.040 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 93.840 700.000 94.440 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 97.240 700.000 97.840 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 6.120 700.000 6.720 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 100.640 700.000 101.240 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 104.040 700.000 104.640 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 9.520 700.000 10.120 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 12.920 700.000 13.520 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 16.320 700.000 16.920 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 19.720 700.000 20.320 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 23.120 700.000 23.720 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 26.520 700.000 27.120 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 29.920 700.000 30.520 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 339.320 700.000 339.920 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 107.440 700.000 108.040 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 140.760 700.000 141.360 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 144.160 700.000 144.760 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 147.560 700.000 148.160 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 150.960 700.000 151.560 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 154.360 700.000 154.960 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 157.760 700.000 158.360 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 161.160 700.000 161.760 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 164.560 700.000 165.160 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 167.960 700.000 168.560 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 171.360 700.000 171.960 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 110.840 700.000 111.440 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 174.080 700.000 174.680 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 177.480 700.000 178.080 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 180.880 700.000 181.480 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 184.280 700.000 184.880 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 187.680 700.000 188.280 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 191.080 700.000 191.680 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 194.480 700.000 195.080 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 197.880 700.000 198.480 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 201.280 700.000 201.880 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 204.680 700.000 205.280 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 114.240 700.000 114.840 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 208.080 700.000 208.680 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 211.480 700.000 212.080 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 116.960 700.000 117.560 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 120.360 700.000 120.960 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 123.760 700.000 124.360 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 127.160 700.000 127.760 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 130.560 700.000 131.160 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 133.960 700.000 134.560 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 137.360 700.000 137.960 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 332.520 700.000 333.120 ;
    END
  END HREADY
  PIN HREADYOUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.320 4.000 390.920 ;
    END
  END HREADYOUT
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 342.720 700.000 343.320 ;
    END
  END HRESETn
  PIN HSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 335.920 700.000 336.520 ;
    END
  END HSEL
  PIN HTRANS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 322.320 700.000 322.920 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 325.720 700.000 326.320 ;
    END
  END HTRANS[1]
  PIN HWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 214.880 700.000 215.480 ;
    END
  END HWDATA[0]
  PIN HWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 248.200 700.000 248.800 ;
    END
  END HWDATA[10]
  PIN HWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 251.600 700.000 252.200 ;
    END
  END HWDATA[11]
  PIN HWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 255.000 700.000 255.600 ;
    END
  END HWDATA[12]
  PIN HWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 258.400 700.000 259.000 ;
    END
  END HWDATA[13]
  PIN HWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 261.800 700.000 262.400 ;
    END
  END HWDATA[14]
  PIN HWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 265.200 700.000 265.800 ;
    END
  END HWDATA[15]
  PIN HWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 268.600 700.000 269.200 ;
    END
  END HWDATA[16]
  PIN HWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 272.000 700.000 272.600 ;
    END
  END HWDATA[17]
  PIN HWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 275.400 700.000 276.000 ;
    END
  END HWDATA[18]
  PIN HWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 278.800 700.000 279.400 ;
    END
  END HWDATA[19]
  PIN HWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 218.280 700.000 218.880 ;
    END
  END HWDATA[1]
  PIN HWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 282.200 700.000 282.800 ;
    END
  END HWDATA[20]
  PIN HWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 285.600 700.000 286.200 ;
    END
  END HWDATA[21]
  PIN HWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 288.320 700.000 288.920 ;
    END
  END HWDATA[22]
  PIN HWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 291.720 700.000 292.320 ;
    END
  END HWDATA[23]
  PIN HWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 295.120 700.000 295.720 ;
    END
  END HWDATA[24]
  PIN HWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 298.520 700.000 299.120 ;
    END
  END HWDATA[25]
  PIN HWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 301.920 700.000 302.520 ;
    END
  END HWDATA[26]
  PIN HWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 305.320 700.000 305.920 ;
    END
  END HWDATA[27]
  PIN HWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 308.720 700.000 309.320 ;
    END
  END HWDATA[28]
  PIN HWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 312.120 700.000 312.720 ;
    END
  END HWDATA[29]
  PIN HWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 221.680 700.000 222.280 ;
    END
  END HWDATA[2]
  PIN HWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 315.520 700.000 316.120 ;
    END
  END HWDATA[30]
  PIN HWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 318.920 700.000 319.520 ;
    END
  END HWDATA[31]
  PIN HWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 225.080 700.000 225.680 ;
    END
  END HWDATA[3]
  PIN HWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 228.480 700.000 229.080 ;
    END
  END HWDATA[4]
  PIN HWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 231.200 700.000 231.800 ;
    END
  END HWDATA[5]
  PIN HWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 234.600 700.000 235.200 ;
    END
  END HWDATA[6]
  PIN HWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 238.000 700.000 238.600 ;
    END
  END HWDATA[7]
  PIN HWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 241.400 700.000 242.000 ;
    END
  END HWDATA[8]
  PIN HWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 244.800 700.000 245.400 ;
    END
  END HWDATA[9]
  PIN HWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 329.120 700.000 329.720 ;
    END
  END HWRITE
  PIN IRQ[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 345.440 700.000 346.040 ;
    END
  END IRQ[0]
  PIN IRQ[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 379.440 700.000 380.040 ;
    END
  END IRQ[10]
  PIN IRQ[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 382.840 700.000 383.440 ;
    END
  END IRQ[11]
  PIN IRQ[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 386.240 700.000 386.840 ;
    END
  END IRQ[12]
  PIN IRQ[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 389.640 700.000 390.240 ;
    END
  END IRQ[13]
  PIN IRQ[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 393.040 700.000 393.640 ;
    END
  END IRQ[14]
  PIN IRQ[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 396.440 700.000 397.040 ;
    END
  END IRQ[15]
  PIN IRQ[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 348.840 700.000 349.440 ;
    END
  END IRQ[1]
  PIN IRQ[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 352.240 700.000 352.840 ;
    END
  END IRQ[2]
  PIN IRQ[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 355.640 700.000 356.240 ;
    END
  END IRQ[3]
  PIN IRQ[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 359.040 700.000 359.640 ;
    END
  END IRQ[4]
  PIN IRQ[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 362.440 700.000 363.040 ;
    END
  END IRQ[5]
  PIN IRQ[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 365.840 700.000 366.440 ;
    END
  END IRQ[6]
  PIN IRQ[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 369.240 700.000 369.840 ;
    END
  END IRQ[7]
  PIN IRQ[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 372.640 700.000 373.240 ;
    END
  END IRQ[8]
  PIN IRQ[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 376.040 700.000 376.640 ;
    END
  END IRQ[9]
  PIN MSI_S2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.600 4.000 65.200 ;
    END
  END MSI_S2
  PIN MSI_S3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.760 4.000 124.360 ;
    END
  END MSI_S3
  PIN MSO_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.880 4.000 79.480 ;
    END
  END MSO_S2
  PIN MSO_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.720 4.000 139.320 ;
    END
  END MSO_S3
  PIN RsRx_S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.440 4.000 6.040 ;
    END
  END RsRx_S0
  PIN RsRx_S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.680 4.000 35.280 ;
    END
  END RsRx_S1
  PIN RsTx_S0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.720 4.000 20.320 ;
    END
  END RsTx_S0
  PIN RsTx_S1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.640 4.000 50.240 ;
    END
  END RsTx_S1
  PIN SCLK_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.800 4.000 109.400 ;
    END
  END SCLK_S2
  PIN SCLK_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.960 4.000 168.560 ;
    END
  END SCLK_S3
  PIN SSn_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.840 4.000 94.440 ;
    END
  END SSn_S2
  PIN SSn_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.000 4.000 153.600 ;
    END
  END SSn_S3
  PIN pwm_S6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.400 4.000 361.000 ;
    END
  END pwm_S6
  PIN pwm_S7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.360 4.000 375.960 ;
    END
  END pwm_S7
  PIN scl_i_S4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.920 4.000 183.520 ;
    END
  END scl_i_S4
  PIN scl_i_S5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.000 4.000 272.600 ;
    END
  END scl_i_S5
  PIN scl_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.880 4.000 198.480 ;
    END
  END scl_o_S4
  PIN scl_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.280 4.000 286.880 ;
    END
  END scl_o_S5
  PIN scl_oen_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.160 4.000 212.760 ;
    END
  END scl_oen_o_S4
  PIN scl_oen_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.240 4.000 301.840 ;
    END
  END scl_oen_o_S5
  PIN sda_i_S4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.120 4.000 227.720 ;
    END
  END sda_i_S4
  PIN sda_i_S5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.200 4.000 316.800 ;
    END
  END sda_i_S5
  PIN sda_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.080 4.000 242.680 ;
    END
  END sda_o_S4
  PIN sda_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.160 4.000 331.760 ;
    END
  END sda_o_S5
  PIN sda_oen_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.040 4.000 257.640 ;
    END
  END sda_oen_o_S4
  PIN sda_oen_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.440 4.000 346.040 ;
    END
  END sda_oen_o_S5
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 9.240 637.040 387.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 9.240 483.440 387.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 9.240 329.840 387.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 9.240 176.240 387.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 9.240 22.640 387.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 9.240 560.240 387.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 9.240 406.640 387.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 9.240 253.040 387.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 9.240 99.440 387.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 6.845 694.915 387.645 ;
      LAYER met1 ;
        RECT 5.520 4.760 694.990 391.260 ;
      LAYER met2 ;
        RECT 6.990 0.115 694.970 397.605 ;
      LAYER met3 ;
        RECT 3.990 397.440 696.130 398.260 ;
        RECT 3.990 396.040 695.600 397.440 ;
        RECT 3.990 394.040 696.130 396.040 ;
        RECT 3.990 392.640 695.600 394.040 ;
        RECT 3.990 391.320 696.130 392.640 ;
        RECT 4.400 390.640 696.130 391.320 ;
        RECT 4.400 389.920 695.600 390.640 ;
        RECT 3.990 389.240 695.600 389.920 ;
        RECT 3.990 387.240 696.130 389.240 ;
        RECT 3.990 385.840 695.600 387.240 ;
        RECT 3.990 383.840 696.130 385.840 ;
        RECT 3.990 382.440 695.600 383.840 ;
        RECT 3.990 380.440 696.130 382.440 ;
        RECT 3.990 379.040 695.600 380.440 ;
        RECT 3.990 377.040 696.130 379.040 ;
        RECT 3.990 376.360 695.600 377.040 ;
        RECT 4.400 375.640 695.600 376.360 ;
        RECT 4.400 374.960 696.130 375.640 ;
        RECT 3.990 373.640 696.130 374.960 ;
        RECT 3.990 372.240 695.600 373.640 ;
        RECT 3.990 370.240 696.130 372.240 ;
        RECT 3.990 368.840 695.600 370.240 ;
        RECT 3.990 366.840 696.130 368.840 ;
        RECT 3.990 365.440 695.600 366.840 ;
        RECT 3.990 363.440 696.130 365.440 ;
        RECT 3.990 362.040 695.600 363.440 ;
        RECT 3.990 361.400 696.130 362.040 ;
        RECT 4.400 360.040 696.130 361.400 ;
        RECT 4.400 360.000 695.600 360.040 ;
        RECT 3.990 358.640 695.600 360.000 ;
        RECT 3.990 356.640 696.130 358.640 ;
        RECT 3.990 355.240 695.600 356.640 ;
        RECT 3.990 353.240 696.130 355.240 ;
        RECT 3.990 351.840 695.600 353.240 ;
        RECT 3.990 349.840 696.130 351.840 ;
        RECT 3.990 348.440 695.600 349.840 ;
        RECT 3.990 346.440 696.130 348.440 ;
        RECT 4.400 345.040 695.600 346.440 ;
        RECT 3.990 343.720 696.130 345.040 ;
        RECT 3.990 342.320 695.600 343.720 ;
        RECT 3.990 340.320 696.130 342.320 ;
        RECT 3.990 338.920 695.600 340.320 ;
        RECT 3.990 336.920 696.130 338.920 ;
        RECT 3.990 335.520 695.600 336.920 ;
        RECT 3.990 333.520 696.130 335.520 ;
        RECT 3.990 332.160 695.600 333.520 ;
        RECT 4.400 332.120 695.600 332.160 ;
        RECT 4.400 330.760 696.130 332.120 ;
        RECT 3.990 330.120 696.130 330.760 ;
        RECT 3.990 328.720 695.600 330.120 ;
        RECT 3.990 326.720 696.130 328.720 ;
        RECT 3.990 325.320 695.600 326.720 ;
        RECT 3.990 323.320 696.130 325.320 ;
        RECT 3.990 321.920 695.600 323.320 ;
        RECT 3.990 319.920 696.130 321.920 ;
        RECT 3.990 318.520 695.600 319.920 ;
        RECT 3.990 317.200 696.130 318.520 ;
        RECT 4.400 316.520 696.130 317.200 ;
        RECT 4.400 315.800 695.600 316.520 ;
        RECT 3.990 315.120 695.600 315.800 ;
        RECT 3.990 313.120 696.130 315.120 ;
        RECT 3.990 311.720 695.600 313.120 ;
        RECT 3.990 309.720 696.130 311.720 ;
        RECT 3.990 308.320 695.600 309.720 ;
        RECT 3.990 306.320 696.130 308.320 ;
        RECT 3.990 304.920 695.600 306.320 ;
        RECT 3.990 302.920 696.130 304.920 ;
        RECT 3.990 302.240 695.600 302.920 ;
        RECT 4.400 301.520 695.600 302.240 ;
        RECT 4.400 300.840 696.130 301.520 ;
        RECT 3.990 299.520 696.130 300.840 ;
        RECT 3.990 298.120 695.600 299.520 ;
        RECT 3.990 296.120 696.130 298.120 ;
        RECT 3.990 294.720 695.600 296.120 ;
        RECT 3.990 292.720 696.130 294.720 ;
        RECT 3.990 291.320 695.600 292.720 ;
        RECT 3.990 289.320 696.130 291.320 ;
        RECT 3.990 287.920 695.600 289.320 ;
        RECT 3.990 287.280 696.130 287.920 ;
        RECT 4.400 286.600 696.130 287.280 ;
        RECT 4.400 285.880 695.600 286.600 ;
        RECT 3.990 285.200 695.600 285.880 ;
        RECT 3.990 283.200 696.130 285.200 ;
        RECT 3.990 281.800 695.600 283.200 ;
        RECT 3.990 279.800 696.130 281.800 ;
        RECT 3.990 278.400 695.600 279.800 ;
        RECT 3.990 276.400 696.130 278.400 ;
        RECT 3.990 275.000 695.600 276.400 ;
        RECT 3.990 273.000 696.130 275.000 ;
        RECT 4.400 271.600 695.600 273.000 ;
        RECT 3.990 269.600 696.130 271.600 ;
        RECT 3.990 268.200 695.600 269.600 ;
        RECT 3.990 266.200 696.130 268.200 ;
        RECT 3.990 264.800 695.600 266.200 ;
        RECT 3.990 262.800 696.130 264.800 ;
        RECT 3.990 261.400 695.600 262.800 ;
        RECT 3.990 259.400 696.130 261.400 ;
        RECT 3.990 258.040 695.600 259.400 ;
        RECT 4.400 258.000 695.600 258.040 ;
        RECT 4.400 256.640 696.130 258.000 ;
        RECT 3.990 256.000 696.130 256.640 ;
        RECT 3.990 254.600 695.600 256.000 ;
        RECT 3.990 252.600 696.130 254.600 ;
        RECT 3.990 251.200 695.600 252.600 ;
        RECT 3.990 249.200 696.130 251.200 ;
        RECT 3.990 247.800 695.600 249.200 ;
        RECT 3.990 245.800 696.130 247.800 ;
        RECT 3.990 244.400 695.600 245.800 ;
        RECT 3.990 243.080 696.130 244.400 ;
        RECT 4.400 242.400 696.130 243.080 ;
        RECT 4.400 241.680 695.600 242.400 ;
        RECT 3.990 241.000 695.600 241.680 ;
        RECT 3.990 239.000 696.130 241.000 ;
        RECT 3.990 237.600 695.600 239.000 ;
        RECT 3.990 235.600 696.130 237.600 ;
        RECT 3.990 234.200 695.600 235.600 ;
        RECT 3.990 232.200 696.130 234.200 ;
        RECT 3.990 230.800 695.600 232.200 ;
        RECT 3.990 229.480 696.130 230.800 ;
        RECT 3.990 228.120 695.600 229.480 ;
        RECT 4.400 228.080 695.600 228.120 ;
        RECT 4.400 226.720 696.130 228.080 ;
        RECT 3.990 226.080 696.130 226.720 ;
        RECT 3.990 224.680 695.600 226.080 ;
        RECT 3.990 222.680 696.130 224.680 ;
        RECT 3.990 221.280 695.600 222.680 ;
        RECT 3.990 219.280 696.130 221.280 ;
        RECT 3.990 217.880 695.600 219.280 ;
        RECT 3.990 215.880 696.130 217.880 ;
        RECT 3.990 214.480 695.600 215.880 ;
        RECT 3.990 213.160 696.130 214.480 ;
        RECT 4.400 212.480 696.130 213.160 ;
        RECT 4.400 211.760 695.600 212.480 ;
        RECT 3.990 211.080 695.600 211.760 ;
        RECT 3.990 209.080 696.130 211.080 ;
        RECT 3.990 207.680 695.600 209.080 ;
        RECT 3.990 205.680 696.130 207.680 ;
        RECT 3.990 204.280 695.600 205.680 ;
        RECT 3.990 202.280 696.130 204.280 ;
        RECT 3.990 200.880 695.600 202.280 ;
        RECT 3.990 198.880 696.130 200.880 ;
        RECT 4.400 197.480 695.600 198.880 ;
        RECT 3.990 195.480 696.130 197.480 ;
        RECT 3.990 194.080 695.600 195.480 ;
        RECT 3.990 192.080 696.130 194.080 ;
        RECT 3.990 190.680 695.600 192.080 ;
        RECT 3.990 188.680 696.130 190.680 ;
        RECT 3.990 187.280 695.600 188.680 ;
        RECT 3.990 185.280 696.130 187.280 ;
        RECT 3.990 183.920 695.600 185.280 ;
        RECT 4.400 183.880 695.600 183.920 ;
        RECT 4.400 182.520 696.130 183.880 ;
        RECT 3.990 181.880 696.130 182.520 ;
        RECT 3.990 180.480 695.600 181.880 ;
        RECT 3.990 178.480 696.130 180.480 ;
        RECT 3.990 177.080 695.600 178.480 ;
        RECT 3.990 175.080 696.130 177.080 ;
        RECT 3.990 173.680 695.600 175.080 ;
        RECT 3.990 172.360 696.130 173.680 ;
        RECT 3.990 170.960 695.600 172.360 ;
        RECT 3.990 168.960 696.130 170.960 ;
        RECT 4.400 167.560 695.600 168.960 ;
        RECT 3.990 165.560 696.130 167.560 ;
        RECT 3.990 164.160 695.600 165.560 ;
        RECT 3.990 162.160 696.130 164.160 ;
        RECT 3.990 160.760 695.600 162.160 ;
        RECT 3.990 158.760 696.130 160.760 ;
        RECT 3.990 157.360 695.600 158.760 ;
        RECT 3.990 155.360 696.130 157.360 ;
        RECT 3.990 154.000 695.600 155.360 ;
        RECT 4.400 153.960 695.600 154.000 ;
        RECT 4.400 152.600 696.130 153.960 ;
        RECT 3.990 151.960 696.130 152.600 ;
        RECT 3.990 150.560 695.600 151.960 ;
        RECT 3.990 148.560 696.130 150.560 ;
        RECT 3.990 147.160 695.600 148.560 ;
        RECT 3.990 145.160 696.130 147.160 ;
        RECT 3.990 143.760 695.600 145.160 ;
        RECT 3.990 141.760 696.130 143.760 ;
        RECT 3.990 140.360 695.600 141.760 ;
        RECT 3.990 139.720 696.130 140.360 ;
        RECT 4.400 138.360 696.130 139.720 ;
        RECT 4.400 138.320 695.600 138.360 ;
        RECT 3.990 136.960 695.600 138.320 ;
        RECT 3.990 134.960 696.130 136.960 ;
        RECT 3.990 133.560 695.600 134.960 ;
        RECT 3.990 131.560 696.130 133.560 ;
        RECT 3.990 130.160 695.600 131.560 ;
        RECT 3.990 128.160 696.130 130.160 ;
        RECT 3.990 126.760 695.600 128.160 ;
        RECT 3.990 124.760 696.130 126.760 ;
        RECT 4.400 123.360 695.600 124.760 ;
        RECT 3.990 121.360 696.130 123.360 ;
        RECT 3.990 119.960 695.600 121.360 ;
        RECT 3.990 117.960 696.130 119.960 ;
        RECT 3.990 116.560 695.600 117.960 ;
        RECT 3.990 115.240 696.130 116.560 ;
        RECT 3.990 113.840 695.600 115.240 ;
        RECT 3.990 111.840 696.130 113.840 ;
        RECT 3.990 110.440 695.600 111.840 ;
        RECT 3.990 109.800 696.130 110.440 ;
        RECT 4.400 108.440 696.130 109.800 ;
        RECT 4.400 108.400 695.600 108.440 ;
        RECT 3.990 107.040 695.600 108.400 ;
        RECT 3.990 105.040 696.130 107.040 ;
        RECT 3.990 103.640 695.600 105.040 ;
        RECT 3.990 101.640 696.130 103.640 ;
        RECT 3.990 100.240 695.600 101.640 ;
        RECT 3.990 98.240 696.130 100.240 ;
        RECT 3.990 96.840 695.600 98.240 ;
        RECT 3.990 94.840 696.130 96.840 ;
        RECT 4.400 93.440 695.600 94.840 ;
        RECT 3.990 91.440 696.130 93.440 ;
        RECT 3.990 90.040 695.600 91.440 ;
        RECT 3.990 88.040 696.130 90.040 ;
        RECT 3.990 86.640 695.600 88.040 ;
        RECT 3.990 84.640 696.130 86.640 ;
        RECT 3.990 83.240 695.600 84.640 ;
        RECT 3.990 81.240 696.130 83.240 ;
        RECT 3.990 79.880 695.600 81.240 ;
        RECT 4.400 79.840 695.600 79.880 ;
        RECT 4.400 78.480 696.130 79.840 ;
        RECT 3.990 77.840 696.130 78.480 ;
        RECT 3.990 76.440 695.600 77.840 ;
        RECT 3.990 74.440 696.130 76.440 ;
        RECT 3.990 73.040 695.600 74.440 ;
        RECT 3.990 71.040 696.130 73.040 ;
        RECT 3.990 69.640 695.600 71.040 ;
        RECT 3.990 67.640 696.130 69.640 ;
        RECT 3.990 66.240 695.600 67.640 ;
        RECT 3.990 65.600 696.130 66.240 ;
        RECT 4.400 64.240 696.130 65.600 ;
        RECT 4.400 64.200 695.600 64.240 ;
        RECT 3.990 62.840 695.600 64.200 ;
        RECT 3.990 60.840 696.130 62.840 ;
        RECT 3.990 59.440 695.600 60.840 ;
        RECT 3.990 58.120 696.130 59.440 ;
        RECT 3.990 56.720 695.600 58.120 ;
        RECT 3.990 54.720 696.130 56.720 ;
        RECT 3.990 53.320 695.600 54.720 ;
        RECT 3.990 51.320 696.130 53.320 ;
        RECT 3.990 50.640 695.600 51.320 ;
        RECT 4.400 49.920 695.600 50.640 ;
        RECT 4.400 49.240 696.130 49.920 ;
        RECT 3.990 47.920 696.130 49.240 ;
        RECT 3.990 46.520 695.600 47.920 ;
        RECT 3.990 44.520 696.130 46.520 ;
        RECT 3.990 43.120 695.600 44.520 ;
        RECT 3.990 41.120 696.130 43.120 ;
        RECT 3.990 39.720 695.600 41.120 ;
        RECT 3.990 37.720 696.130 39.720 ;
        RECT 3.990 36.320 695.600 37.720 ;
        RECT 3.990 35.680 696.130 36.320 ;
        RECT 4.400 34.320 696.130 35.680 ;
        RECT 4.400 34.280 695.600 34.320 ;
        RECT 3.990 32.920 695.600 34.280 ;
        RECT 3.990 30.920 696.130 32.920 ;
        RECT 3.990 29.520 695.600 30.920 ;
        RECT 3.990 27.520 696.130 29.520 ;
        RECT 3.990 26.120 695.600 27.520 ;
        RECT 3.990 24.120 696.130 26.120 ;
        RECT 3.990 22.720 695.600 24.120 ;
        RECT 3.990 20.720 696.130 22.720 ;
        RECT 4.400 19.320 695.600 20.720 ;
        RECT 3.990 17.320 696.130 19.320 ;
        RECT 3.990 15.920 695.600 17.320 ;
        RECT 3.990 13.920 696.130 15.920 ;
        RECT 3.990 12.520 695.600 13.920 ;
        RECT 3.990 10.520 696.130 12.520 ;
        RECT 3.990 9.120 695.600 10.520 ;
        RECT 3.990 7.120 696.130 9.120 ;
        RECT 3.990 6.440 695.600 7.120 ;
        RECT 4.400 5.720 695.600 6.440 ;
        RECT 4.400 5.040 696.130 5.720 ;
        RECT 3.990 3.720 696.130 5.040 ;
        RECT 3.990 2.320 695.600 3.720 ;
        RECT 3.990 1.000 696.130 2.320 ;
        RECT 3.990 0.135 695.600 1.000 ;
      LAYER met4 ;
        RECT 100.575 388.200 686.945 398.265 ;
        RECT 100.575 8.840 174.240 388.200 ;
        RECT 176.640 8.840 251.040 388.200 ;
        RECT 253.440 8.840 327.840 388.200 ;
        RECT 330.240 8.840 404.640 388.200 ;
        RECT 407.040 8.840 481.440 388.200 ;
        RECT 483.840 8.840 558.240 388.200 ;
        RECT 560.640 8.840 635.040 388.200 ;
        RECT 637.440 8.840 686.945 388.200 ;
        RECT 100.575 6.255 686.945 8.840 ;
  END
END apb_sys_0
END LIBRARY

