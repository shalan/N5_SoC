magic
tech sky130A
magscale 1 2
timestamp 1609330474
<< obsli1 >>
rect 38 117 247949 255287
<< obsm1 >>
rect 38 6 247961 256554
<< metal2 >>
rect 424 257158 480 257958
rect 3460 257158 3516 257958
rect 6588 257158 6644 257958
rect 9716 257158 9772 257958
rect 12844 257158 12900 257958
rect 15972 257158 16028 257958
rect 19100 257158 19156 257958
rect 22228 257158 22284 257958
rect 25356 257158 25412 257958
rect 28484 257158 28540 257958
rect 31612 257158 31668 257958
rect 34740 257158 34796 257958
rect 37868 257158 37924 257958
rect 40996 257158 41052 257958
rect 44124 257158 44180 257958
rect 47252 257158 47308 257958
rect 50380 257158 50436 257958
rect 53508 257158 53564 257958
rect 56636 257158 56692 257958
rect 59764 257158 59820 257958
rect 62892 257158 62948 257958
rect 66020 257158 66076 257958
rect 69148 257158 69204 257958
rect 72276 257158 72332 257958
rect 75404 257158 75460 257958
rect 78532 257158 78588 257958
rect 81660 257158 81716 257958
rect 84696 257158 84752 257958
rect 87824 257158 87880 257958
rect 90952 257158 91008 257958
rect 94080 257158 94136 257958
rect 97208 257158 97264 257958
rect 100336 257158 100392 257958
rect 103464 257158 103520 257958
rect 106592 257158 106648 257958
rect 109720 257158 109776 257958
rect 112848 257158 112904 257958
rect 115976 257158 116032 257958
rect 119104 257158 119160 257958
rect 122232 257158 122288 257958
rect 125360 257158 125416 257958
rect 128488 257158 128544 257958
rect 131616 257158 131672 257958
rect 134744 257158 134800 257958
rect 137872 257158 137928 257958
rect 141000 257158 141056 257958
rect 144128 257158 144184 257958
rect 147256 257158 147312 257958
rect 150384 257158 150440 257958
rect 153512 257158 153568 257958
rect 156640 257158 156696 257958
rect 159768 257158 159824 257958
rect 162896 257158 162952 257958
rect 166024 257158 166080 257958
rect 169060 257158 169116 257958
rect 172188 257158 172244 257958
rect 175316 257158 175372 257958
rect 178444 257158 178500 257958
rect 181572 257158 181628 257958
rect 184700 257158 184756 257958
rect 187828 257158 187884 257958
rect 190956 257158 191012 257958
rect 194084 257158 194140 257958
rect 197212 257158 197268 257958
rect 200340 257158 200396 257958
rect 203468 257158 203524 257958
rect 206596 257158 206652 257958
rect 209724 257158 209780 257958
rect 212852 257158 212908 257958
rect 215980 257158 216036 257958
rect 219108 257158 219164 257958
rect 222236 257158 222292 257958
rect 225364 257158 225420 257958
rect 228492 257158 228548 257958
rect 231620 257158 231676 257958
rect 234748 257158 234804 257958
rect 237876 257158 237932 257958
rect 241004 257158 241060 257958
rect 244132 257158 244188 257958
rect 247260 257158 247316 257958
<< obsm2 >>
rect 334 257102 368 257158
rect 536 257102 3404 257158
rect 3572 257102 6532 257158
rect 6700 257102 9660 257158
rect 9828 257102 12788 257158
rect 12956 257102 15916 257158
rect 16084 257102 19044 257158
rect 19212 257102 22172 257158
rect 22340 257102 25300 257158
rect 25468 257102 28428 257158
rect 28596 257102 31556 257158
rect 31724 257102 34684 257158
rect 34852 257102 37812 257158
rect 37980 257102 40940 257158
rect 41108 257102 44068 257158
rect 44236 257102 47196 257158
rect 47364 257102 50324 257158
rect 50492 257102 53452 257158
rect 53620 257102 56580 257158
rect 56748 257102 59708 257158
rect 59876 257102 62836 257158
rect 63004 257102 65964 257158
rect 66132 257102 69092 257158
rect 69260 257102 72220 257158
rect 72388 257102 75348 257158
rect 75516 257102 78476 257158
rect 78644 257102 81604 257158
rect 81772 257102 84640 257158
rect 84808 257102 87768 257158
rect 87936 257102 90896 257158
rect 91064 257102 94024 257158
rect 94192 257102 97152 257158
rect 97320 257102 100280 257158
rect 100448 257102 103408 257158
rect 103576 257102 106536 257158
rect 106704 257102 109664 257158
rect 109832 257102 112792 257158
rect 112960 257102 115920 257158
rect 116088 257102 119048 257158
rect 119216 257102 122176 257158
rect 122344 257102 125304 257158
rect 125472 257102 128432 257158
rect 128600 257102 131560 257158
rect 131728 257102 134688 257158
rect 134856 257102 137816 257158
rect 137984 257102 140944 257158
rect 141112 257102 144072 257158
rect 144240 257102 147200 257158
rect 147368 257102 150328 257158
rect 150496 257102 153456 257158
rect 153624 257102 156584 257158
rect 156752 257102 159712 257158
rect 159880 257102 162840 257158
rect 163008 257102 165968 257158
rect 166136 257102 169004 257158
rect 169172 257102 172132 257158
rect 172300 257102 175260 257158
rect 175428 257102 178388 257158
rect 178556 257102 181516 257158
rect 181684 257102 184644 257158
rect 184812 257102 187772 257158
rect 187940 257102 190900 257158
rect 191068 257102 194028 257158
rect 194196 257102 197156 257158
rect 197324 257102 200284 257158
rect 200452 257102 203412 257158
rect 203580 257102 206540 257158
rect 206708 257102 209668 257158
rect 209836 257102 212796 257158
rect 212964 257102 215924 257158
rect 216092 257102 219052 257158
rect 219220 257102 222180 257158
rect 222348 257102 225308 257158
rect 225476 257102 228436 257158
rect 228604 257102 231564 257158
rect 231732 257102 234692 257158
rect 234860 257102 237820 257158
rect 237988 257102 240948 257158
rect 241116 257102 244076 257158
rect 244244 257102 247204 257158
rect 247372 257102 247498 257158
rect 334 0 247498 257102
<< obsm3 >>
rect 603 101 247229 255303
<< metal4 >>
rect 3142 86 3462 255318
rect 15142 86 15462 255318
rect 27142 86 27462 255318
rect 39142 86 39462 255318
rect 51142 86 51462 255318
rect 63142 86 63462 255318
rect 75142 86 75462 255318
rect 87142 86 87462 255318
rect 99142 86 99462 255318
rect 111142 86 111462 255318
rect 123142 86 123462 255318
rect 135142 86 135462 255318
rect 147142 86 147462 255318
rect 159142 86 159462 255318
rect 171142 86 171462 255318
rect 183142 86 183462 255318
rect 195142 86 195462 255318
rect 207142 86 207462 255318
rect 219142 86 219462 255318
rect 231142 86 231462 255318
rect 243142 86 243462 255318
<< obsm4 >>
rect 1017 3569 3062 254555
rect 3542 3569 15062 254555
rect 15542 3569 27062 254555
rect 27542 3569 39062 254555
rect 39542 3569 51062 254555
rect 51542 3569 63062 254555
rect 63542 3569 75062 254555
rect 75542 3569 87062 254555
rect 87542 3569 99062 254555
rect 99542 3569 111062 254555
rect 111542 3569 123062 254555
rect 123542 3569 135062 254555
rect 135542 3569 147062 254555
rect 147542 3569 159062 254555
rect 159542 3569 171062 254555
rect 171542 3569 183062 254555
rect 183542 3569 195062 254555
rect 195542 3569 207062 254555
rect 207542 3569 219062 254555
rect 219542 3569 231062 254555
rect 231542 3569 242859 254555
<< labels >>
rlabel metal2 s 100336 257158 100392 257958 6 A[0]
port 1 nsew signal input
rlabel metal2 s 103464 257158 103520 257958 6 A[1]
port 2 nsew signal input
rlabel metal2 s 106592 257158 106648 257958 6 A[2]
port 3 nsew signal input
rlabel metal2 s 109720 257158 109776 257958 6 A[3]
port 4 nsew signal input
rlabel metal2 s 112848 257158 112904 257958 6 A[4]
port 5 nsew signal input
rlabel metal2 s 115976 257158 116032 257958 6 A[5]
port 6 nsew signal input
rlabel metal2 s 119104 257158 119160 257958 6 A[6]
port 7 nsew signal input
rlabel metal2 s 122232 257158 122288 257958 6 A[7]
port 8 nsew signal input
rlabel metal2 s 125360 257158 125416 257958 6 A[8]
port 9 nsew signal input
rlabel metal2 s 128488 257158 128544 257958 6 A[9]
port 10 nsew signal input
rlabel metal2 s 131616 257158 131672 257958 6 CLK
port 11 nsew signal input
rlabel metal2 s 150384 257158 150440 257958 6 Di[0]
port 12 nsew signal input
rlabel metal2 s 181572 257158 181628 257958 6 Di[10]
port 13 nsew signal input
rlabel metal2 s 184700 257158 184756 257958 6 Di[11]
port 14 nsew signal input
rlabel metal2 s 187828 257158 187884 257958 6 Di[12]
port 15 nsew signal input
rlabel metal2 s 190956 257158 191012 257958 6 Di[13]
port 16 nsew signal input
rlabel metal2 s 194084 257158 194140 257958 6 Di[14]
port 17 nsew signal input
rlabel metal2 s 197212 257158 197268 257958 6 Di[15]
port 18 nsew signal input
rlabel metal2 s 200340 257158 200396 257958 6 Di[16]
port 19 nsew signal input
rlabel metal2 s 203468 257158 203524 257958 6 Di[17]
port 20 nsew signal input
rlabel metal2 s 206596 257158 206652 257958 6 Di[18]
port 21 nsew signal input
rlabel metal2 s 209724 257158 209780 257958 6 Di[19]
port 22 nsew signal input
rlabel metal2 s 153512 257158 153568 257958 6 Di[1]
port 23 nsew signal input
rlabel metal2 s 212852 257158 212908 257958 6 Di[20]
port 24 nsew signal input
rlabel metal2 s 215980 257158 216036 257958 6 Di[21]
port 25 nsew signal input
rlabel metal2 s 219108 257158 219164 257958 6 Di[22]
port 26 nsew signal input
rlabel metal2 s 222236 257158 222292 257958 6 Di[23]
port 27 nsew signal input
rlabel metal2 s 225364 257158 225420 257958 6 Di[24]
port 28 nsew signal input
rlabel metal2 s 228492 257158 228548 257958 6 Di[25]
port 29 nsew signal input
rlabel metal2 s 231620 257158 231676 257958 6 Di[26]
port 30 nsew signal input
rlabel metal2 s 234748 257158 234804 257958 6 Di[27]
port 31 nsew signal input
rlabel metal2 s 237876 257158 237932 257958 6 Di[28]
port 32 nsew signal input
rlabel metal2 s 241004 257158 241060 257958 6 Di[29]
port 33 nsew signal input
rlabel metal2 s 156640 257158 156696 257958 6 Di[2]
port 34 nsew signal input
rlabel metal2 s 244132 257158 244188 257958 6 Di[30]
port 35 nsew signal input
rlabel metal2 s 247260 257158 247316 257958 6 Di[31]
port 36 nsew signal input
rlabel metal2 s 159768 257158 159824 257958 6 Di[3]
port 37 nsew signal input
rlabel metal2 s 162896 257158 162952 257958 6 Di[4]
port 38 nsew signal input
rlabel metal2 s 166024 257158 166080 257958 6 Di[5]
port 39 nsew signal input
rlabel metal2 s 169060 257158 169116 257958 6 Di[6]
port 40 nsew signal input
rlabel metal2 s 172188 257158 172244 257958 6 Di[7]
port 41 nsew signal input
rlabel metal2 s 175316 257158 175372 257958 6 Di[8]
port 42 nsew signal input
rlabel metal2 s 178444 257158 178500 257958 6 Di[9]
port 43 nsew signal input
rlabel metal2 s 424 257158 480 257958 6 Do[0]
port 44 nsew signal output
rlabel metal2 s 31612 257158 31668 257958 6 Do[10]
port 45 nsew signal output
rlabel metal2 s 34740 257158 34796 257958 6 Do[11]
port 46 nsew signal output
rlabel metal2 s 37868 257158 37924 257958 6 Do[12]
port 47 nsew signal output
rlabel metal2 s 40996 257158 41052 257958 6 Do[13]
port 48 nsew signal output
rlabel metal2 s 44124 257158 44180 257958 6 Do[14]
port 49 nsew signal output
rlabel metal2 s 47252 257158 47308 257958 6 Do[15]
port 50 nsew signal output
rlabel metal2 s 50380 257158 50436 257958 6 Do[16]
port 51 nsew signal output
rlabel metal2 s 53508 257158 53564 257958 6 Do[17]
port 52 nsew signal output
rlabel metal2 s 56636 257158 56692 257958 6 Do[18]
port 53 nsew signal output
rlabel metal2 s 59764 257158 59820 257958 6 Do[19]
port 54 nsew signal output
rlabel metal2 s 3460 257158 3516 257958 6 Do[1]
port 55 nsew signal output
rlabel metal2 s 62892 257158 62948 257958 6 Do[20]
port 56 nsew signal output
rlabel metal2 s 66020 257158 66076 257958 6 Do[21]
port 57 nsew signal output
rlabel metal2 s 69148 257158 69204 257958 6 Do[22]
port 58 nsew signal output
rlabel metal2 s 72276 257158 72332 257958 6 Do[23]
port 59 nsew signal output
rlabel metal2 s 75404 257158 75460 257958 6 Do[24]
port 60 nsew signal output
rlabel metal2 s 78532 257158 78588 257958 6 Do[25]
port 61 nsew signal output
rlabel metal2 s 81660 257158 81716 257958 6 Do[26]
port 62 nsew signal output
rlabel metal2 s 84696 257158 84752 257958 6 Do[27]
port 63 nsew signal output
rlabel metal2 s 87824 257158 87880 257958 6 Do[28]
port 64 nsew signal output
rlabel metal2 s 90952 257158 91008 257958 6 Do[29]
port 65 nsew signal output
rlabel metal2 s 6588 257158 6644 257958 6 Do[2]
port 66 nsew signal output
rlabel metal2 s 94080 257158 94136 257958 6 Do[30]
port 67 nsew signal output
rlabel metal2 s 97208 257158 97264 257958 6 Do[31]
port 68 nsew signal output
rlabel metal2 s 9716 257158 9772 257958 6 Do[3]
port 69 nsew signal output
rlabel metal2 s 12844 257158 12900 257958 6 Do[4]
port 70 nsew signal output
rlabel metal2 s 15972 257158 16028 257958 6 Do[5]
port 71 nsew signal output
rlabel metal2 s 19100 257158 19156 257958 6 Do[6]
port 72 nsew signal output
rlabel metal2 s 22228 257158 22284 257958 6 Do[7]
port 73 nsew signal output
rlabel metal2 s 25356 257158 25412 257958 6 Do[8]
port 74 nsew signal output
rlabel metal2 s 28484 257158 28540 257958 6 Do[9]
port 75 nsew signal output
rlabel metal2 s 147256 257158 147312 257958 6 EN
port 76 nsew signal input
rlabel metal2 s 134744 257158 134800 257958 6 WE[0]
port 77 nsew signal input
rlabel metal2 s 137872 257158 137928 257958 6 WE[1]
port 78 nsew signal input
rlabel metal2 s 141000 257158 141056 257958 6 WE[2]
port 79 nsew signal input
rlabel metal2 s 144128 257158 144184 257958 6 WE[3]
port 80 nsew signal input
rlabel metal4 s 243142 86 243462 255318 6 VPWR
port 81 nsew power bidirectional
rlabel metal4 s 219142 86 219462 255318 6 VPWR
port 82 nsew power bidirectional
rlabel metal4 s 195142 86 195462 255318 6 VPWR
port 83 nsew power bidirectional
rlabel metal4 s 171142 86 171462 255318 6 VPWR
port 84 nsew power bidirectional
rlabel metal4 s 147142 86 147462 255318 6 VPWR
port 85 nsew power bidirectional
rlabel metal4 s 123142 86 123462 255318 6 VPWR
port 86 nsew power bidirectional
rlabel metal4 s 99142 86 99462 255318 6 VPWR
port 87 nsew power bidirectional
rlabel metal4 s 75142 86 75462 255318 6 VPWR
port 88 nsew power bidirectional
rlabel metal4 s 51142 86 51462 255318 6 VPWR
port 89 nsew power bidirectional
rlabel metal4 s 27142 86 27462 255318 6 VPWR
port 90 nsew power bidirectional
rlabel metal4 s 3142 86 3462 255318 6 VPWR
port 91 nsew power bidirectional
rlabel metal4 s 231142 86 231462 255318 6 VGND
port 92 nsew ground bidirectional
rlabel metal4 s 207142 86 207462 255318 6 VGND
port 93 nsew ground bidirectional
rlabel metal4 s 183142 86 183462 255318 6 VGND
port 94 nsew ground bidirectional
rlabel metal4 s 159142 86 159462 255318 6 VGND
port 95 nsew ground bidirectional
rlabel metal4 s 135142 86 135462 255318 6 VGND
port 96 nsew ground bidirectional
rlabel metal4 s 111142 86 111462 255318 6 VGND
port 97 nsew ground bidirectional
rlabel metal4 s 87142 86 87462 255318 6 VGND
port 98 nsew ground bidirectional
rlabel metal4 s 63142 86 63462 255318 6 VGND
port 99 nsew ground bidirectional
rlabel metal4 s 39142 86 39462 255318 6 VGND
port 100 nsew ground bidirectional
rlabel metal4 s 15142 86 15462 255318 6 VGND
port 101 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 247961 257958
string LEFview TRUE
<< end >>
