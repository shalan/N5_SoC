* NGSPICE file created from apb_sys_0.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt apb_sys_0 HADDR[0] HADDR[10] HADDR[11] HADDR[12] HADDR[13] HADDR[14] HADDR[15]
+ HADDR[16] HADDR[17] HADDR[18] HADDR[19] HADDR[1] HADDR[20] HADDR[21] HADDR[22] HADDR[23]
+ HADDR[24] HADDR[25] HADDR[26] HADDR[27] HADDR[28] HADDR[29] HADDR[2] HADDR[30] HADDR[31]
+ HADDR[3] HADDR[4] HADDR[5] HADDR[6] HADDR[7] HADDR[8] HADDR[9] HCLK HRDATA[0] HRDATA[10]
+ HRDATA[11] HRDATA[12] HRDATA[13] HRDATA[14] HRDATA[15] HRDATA[16] HRDATA[17] HRDATA[18]
+ HRDATA[19] HRDATA[1] HRDATA[20] HRDATA[21] HRDATA[22] HRDATA[23] HRDATA[24] HRDATA[25]
+ HRDATA[26] HRDATA[27] HRDATA[28] HRDATA[29] HRDATA[2] HRDATA[30] HRDATA[31] HRDATA[3]
+ HRDATA[4] HRDATA[5] HRDATA[6] HRDATA[7] HRDATA[8] HRDATA[9] HREADY HREADYOUT HRESETn
+ HSEL HTRANS[0] HTRANS[1] HWDATA[0] HWDATA[10] HWDATA[11] HWDATA[12] HWDATA[13] HWDATA[14]
+ HWDATA[15] HWDATA[16] HWDATA[17] HWDATA[18] HWDATA[19] HWDATA[1] HWDATA[20] HWDATA[21]
+ HWDATA[22] HWDATA[23] HWDATA[24] HWDATA[25] HWDATA[26] HWDATA[27] HWDATA[28] HWDATA[29]
+ HWDATA[2] HWDATA[30] HWDATA[31] HWDATA[3] HWDATA[4] HWDATA[5] HWDATA[6] HWDATA[7]
+ HWDATA[8] HWDATA[9] HWRITE IRQ[16] IRQ[17] IRQ[18] IRQ[19] IRQ[20] IRQ[21] IRQ[22]
+ IRQ[23] IRQ[24] IRQ[25] IRQ[26] IRQ[27] IRQ[28] IRQ[29] IRQ[30] IRQ[31] MSI_S2 MSI_S3
+ MSO_S2 MSO_S3 RsRx_S0 RsRx_S1 RsTx_S0 RsTx_S1 SCLK_S2 SCLK_S3 SSn_S2 SSn_S3 pwm_S6
+ pwm_S7 scl_i_S4 scl_i_S5 scl_o_S4 scl_o_S5 scl_oen_o_S4 scl_oen_o_S5 sda_i_S4 sda_i_S5
+ sda_o_S4 sda_o_S5 sda_oen_o_S4 sda_oen_o_S5 VPWR VGND
XANTENNA__13855__A1 _20673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21917__A2 _21916_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15821__A1_N _12293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18243__B1 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18869_ _18868_/X VGND VGND VPWR VPWR _18869_/Y sky130_fd_sc_hd__inv_2
XFILLER_228_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20900_ _20898_/Y _20894_/Y _20899_/X VGND VGND VPWR VPWR _20900_/X sky130_fd_sc_hd__o21a_4
X_21880_ _12807_/X _21879_/X _24262_/Q _21431_/X VGND VGND VPWR VPWR _21880_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_227_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20831_ _24036_/Q _24035_/Q _13640_/B VGND VGND VPWR VPWR _20831_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_208_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24992__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15830__A _11774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20762_ _20753_/X _20761_/X _15593_/A _20757_/X VGND VGND VPWR VPWR _20762_/X sky130_fd_sc_hd__a2bb2o_4
X_23550_ _23534_/CLK _23550_/D VGND VGND VPWR VPWR _19976_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_223_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21551__B _22119_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24921__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22501_ _17358_/A _22430_/X _12772_/A _22299_/X VGND VGND VPWR VPWR _22502_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23481_ _23497_/CLK _20162_/X VGND VGND VPWR VPWR _20161_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_168_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20693_ _13110_/A _13110_/B _13111_/B VGND VGND VPWR VPWR _20693_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_211_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22432_ _22431_/X VGND VGND VPWR VPWR _22432_/X sky130_fd_sc_hd__buf_2
X_25220_ _25113_/CLK _25220_/D HRESETn VGND VGND VPWR VPWR _14091_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_195_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16309__B1 _15946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22363_ _17730_/X _22342_/Y _22349_/Y _22356_/Y _22362_/Y VGND VGND VPWR VPWR _22363_/X
+ sky130_fd_sc_hd__a32o_4
X_25151_ _23926_/CLK _14378_/X HRESETn VGND VGND VPWR VPWR _20430_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21314_ _22712_/A _21313_/X VGND VGND VPWR VPWR _21314_/X sky130_fd_sc_hd__and2_4
X_24102_ _25471_/CLK _24102_/D HRESETn VGND VGND VPWR VPWR _24102_/Q sky130_fd_sc_hd__dfrtp_4
X_25082_ _25081_/CLK _25082_/D HRESETn VGND VGND VPWR VPWR _14615_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23055__B1 _12796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22294_ _22451_/A VGND VGND VPWR VPWR _22294_/X sky130_fd_sc_hd__buf_2
X_24033_ _24032_/CLK _20820_/X HRESETn VGND VGND VPWR VPWR _13125_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_163_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21245_ _21250_/A _21245_/B VGND VGND VPWR VPWR _21245_/X sky130_fd_sc_hd__or2_4
XANTENNA__14181__A _14181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21176_ _21176_/A VGND VGND VPWR VPWR _21955_/A sky130_fd_sc_hd__buf_2
XANTENNA__25027__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20127_ _20127_/A VGND VGND VPWR VPWR _21636_/B sky130_fd_sc_hd__inv_2
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12649__A2 _12626_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20058_ _20053_/X _18328_/X _13829_/A _13260_/B _20055_/X VGND VGND VPWR VPWR _23520_/D
+ sky130_fd_sc_hd__a32o_4
X_24935_ _23476_/CLK _15517_/X HRESETn VGND VGND VPWR VPWR _11673_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_218_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11900_ _19967_/A VGND VGND VPWR VPWR _19603_/A sky130_fd_sc_hd__buf_2
XANTENNA__13525__A _15908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12880_ _12861_/A _12880_/B _12880_/C VGND VGND VPWR VPWR _25393_/D sky130_fd_sc_hd__and3_4
X_24866_ _24866_/CLK _15749_/X HRESETn VGND VGND VPWR VPWR _24866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22838__A _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_128_0_HCLK clkbuf_7_64_0_HCLK/X VGND VGND VPWR VPWR _23644_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11829_/A _24227_/Q _11829_/Y _11830_/Y VGND VGND VPWR VPWR _11831_/X sky130_fd_sc_hd__o22a_4
X_23817_ _23873_/CLK _19214_/X VGND VGND VPWR VPWR _23817_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _24800_/CLK _24797_/D HRESETn VGND VGND VPWR VPWR _24797_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19734__B1 _19711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14550_/A _14550_/B VGND VGND VPWR VPWR _14550_/X sky130_fd_sc_hd__or2_4
XANTENNA__24662__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11759_/Y _11756_/X _11761_/X _11756_/X VGND VGND VPWR VPWR _25527_/D sky130_fd_sc_hd__a2bb2o_4
X_23748_ _24889_/CLK _23748_/D VGND VGND VPWR VPWR _19405_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _25308_/Q VGND VGND VPWR VPWR _13501_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _25114_/Q VGND VGND VPWR VPWR _14481_/Y sky130_fd_sc_hd__inv_2
XPHY_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11690_/Y _11684_/X _11691_/X _11692_/X VGND VGND VPWR VPWR _11693_/X sky130_fd_sc_hd__a2bb2o_4
X_23679_ _23559_/CLK _23679_/D VGND VGND VPWR VPWR _19609_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16219_/Y _16215_/X _15953_/X _16215_/X VGND VGND VPWR VPWR _24664_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _13193_/A _13432_/B _13431_/X VGND VGND VPWR VPWR _13432_/X sky130_fd_sc_hd__and3_4
X_25418_ _25409_/CLK _25418_/D HRESETn VGND VGND VPWR VPWR _25418_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22636__A3 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16151_ _16149_/Y _16150_/X _16059_/X _16150_/X VGND VGND VPWR VPWR _16151_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_139_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12585__B2 _24858_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13363_ _13363_/A _23387_/Q VGND VGND VPWR VPWR _13365_/B sky130_fd_sc_hd__or2_4
X_25349_ _25346_/CLK _25349_/D HRESETn VGND VGND VPWR VPWR _25349_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15102_ _15102_/A _15095_/X _15102_/C _15101_/X VGND VGND VPWR VPWR _15102_/X sky130_fd_sc_hd__or4_4
XFILLER_154_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12314_ _12304_/X _12314_/B _12310_/X _12314_/D VGND VGND VPWR VPWR _12328_/C sky130_fd_sc_hd__or4_4
X_16082_ _22816_/A VGND VGND VPWR VPWR _22505_/B sky130_fd_sc_hd__buf_2
X_13294_ _13363_/A _13294_/B VGND VGND VPWR VPWR _13294_/X sky130_fd_sc_hd__or2_4
X_15033_ _14942_/Y VGND VGND VPWR VPWR _15204_/B sky130_fd_sc_hd__buf_2
X_19910_ _19909_/Y _19905_/X _19820_/X _19905_/X VGND VGND VPWR VPWR _19910_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12245_ _24768_/Q VGND VGND VPWR VPWR _12245_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16721__D _21327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12176_ _12176_/A VGND VGND VPWR VPWR _12428_/C sky130_fd_sc_hd__buf_2
X_19841_ _19839_/Y _19835_/X _19813_/X _19840_/X VGND VGND VPWR VPWR _19841_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25305__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16984_ _24391_/Q VGND VGND VPWR VPWR _16984_/Y sky130_fd_sc_hd__inv_2
X_19772_ _21888_/B _19769_/X _16873_/X _19769_/X VGND VGND VPWR VPWR _23623_/D sky130_fd_sc_hd__a2bb2o_4
X_15935_ _15931_/X VGND VGND VPWR VPWR _15935_/X sky130_fd_sc_hd__buf_2
X_18723_ _18734_/A _18723_/B _18722_/X VGND VGND VPWR VPWR _24153_/D sky130_fd_sc_hd__and3_4
XANTENNA__15635__A2_N _15553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_24_0_HCLK clkbuf_7_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_49_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13435__A _13334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18654_ _18648_/X _18654_/B _18651_/X _18653_/X VGND VGND VPWR VPWR _18669_/B sky130_fd_sc_hd__or4_4
X_15866_ _12747_/Y _15862_/X _15564_/X _15865_/X VGND VGND VPWR VPWR _15866_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_87_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22748__A _24763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14817_ _23994_/Q VGND VGND VPWR VPWR _14817_/X sky130_fd_sc_hd__buf_2
X_17605_ _17561_/Y _17603_/X _17604_/X _17598_/Y VGND VGND VPWR VPWR _17606_/A sky130_fd_sc_hd__a211o_4
X_18585_ _18562_/A _18562_/B _18583_/B _18500_/X VGND VGND VPWR VPWR _18585_/X sky130_fd_sc_hd__a211o_4
X_15797_ _12297_/Y _15793_/X _15564_/X _15796_/X VGND VGND VPWR VPWR _24847_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17536_ _11690_/Y _17563_/A _11690_/Y _17563_/A VGND VGND VPWR VPWR _17536_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19122__A _18981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14748_ _14745_/X VGND VGND VPWR VPWR _14748_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24332__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17467_ _18910_/A _18336_/A _17481_/B VGND VGND VPWR VPWR _17467_/X sky130_fd_sc_hd__a21o_4
X_14679_ _13724_/X _14678_/X _13724_/X _14678_/X VGND VGND VPWR VPWR _14714_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16418_ _16418_/A VGND VGND VPWR VPWR _16418_/X sky130_fd_sc_hd__buf_2
X_19206_ _19205_/Y _19199_/X _19138_/X _19191_/A VGND VGND VPWR VPWR _23819_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22088__A1 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23285__B1 _24113_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17398_ _17398_/A VGND VGND VPWR VPWR _17398_/X sky130_fd_sc_hd__buf_2
X_19137_ _23843_/Q VGND VGND VPWR VPWR _19137_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13773__B1 _13459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16349_ _14380_/A VGND VGND VPWR VPWR _16349_/X sky130_fd_sc_hd__buf_2
XANTENNA__16481__A _24568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25538__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19068_ _19065_/Y _19062_/X _19067_/X _19062_/X VGND VGND VPWR VPWR _19068_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21099__A _22525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18019_ _18060_/A _18016_/X _18019_/C VGND VGND VPWR VPWR _18020_/C sky130_fd_sc_hd__and3_4
XANTENNA__15097__A _24604_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16504__A1_N _16503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21030_ _21030_/A VGND VGND VPWR VPWR _22730_/A sky130_fd_sc_hd__buf_2
XANTENNA__25191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21827__A _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25120__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18201__A _18095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22981_ _22908_/X _22980_/X _22495_/X _25541_/Q _22910_/X VGND VGND VPWR VPWR _22981_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24720_ _24744_/CLK _16066_/X HRESETn VGND VGND VPWR VPWR _24720_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_227_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21932_ _21936_/A _19998_/Y VGND VGND VPWR VPWR _21933_/C sky130_fd_sc_hd__or2_4
XFILLER_215_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24651_ _24654_/CLK _24651_/D HRESETn VGND VGND VPWR VPWR _21842_/A sky130_fd_sc_hd__dfrtp_4
X_21863_ _21127_/X VGND VGND VPWR VPWR _21863_/X sky130_fd_sc_hd__buf_2
XFILLER_24_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23602_ _24199_/CLK _23602_/D VGND VGND VPWR VPWR _23602_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15560__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20814_ _13125_/A _13125_/B _20805_/A VGND VGND VPWR VPWR _20814_/X sky130_fd_sc_hd__or3_4
X_21794_ _21657_/A _19866_/Y VGND VGND VPWR VPWR _21796_/B sky130_fd_sc_hd__or2_4
X_24582_ _24980_/CLK _24582_/D HRESETn VGND VGND VPWR VPWR _15110_/A sky130_fd_sc_hd__dfrtp_4
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23533_ _23411_/CLK _23533_/D VGND VGND VPWR VPWR _20024_/A sky130_fd_sc_hd__dfxtp_4
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24073__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20745_ _13121_/A _13121_/B VGND VGND VPWR VPWR _20749_/A sky130_fd_sc_hd__or2_4
XFILLER_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24002__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20676_ _20510_/B VGND VGND VPWR VPWR _20676_/Y sky130_fd_sc_hd__inv_2
X_23464_ _23464_/CLK _20207_/X VGND VGND VPWR VPWR _18033_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22393__A _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25203_ _25204_/CLK _25203_/D HRESETn VGND VGND VPWR VPWR _14203_/A sky130_fd_sc_hd__dfrtp_4
X_22415_ _22725_/A _22414_/Y VGND VGND VPWR VPWR _22427_/C sky130_fd_sc_hd__nor2_4
XFILLER_148_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23395_ _25272_/CLK _20381_/X VGND VGND VPWR VPWR _23395_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_137_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16391__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25134_ _25134_/CLK _14434_/X HRESETn VGND VGND VPWR VPWR _14433_/A sky130_fd_sc_hd__dfstp_4
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22346_ _21935_/A _22346_/B VGND VGND VPWR VPWR _22348_/B sky130_fd_sc_hd__or2_4
XFILLER_152_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16702__B1 _16522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13516__B1 SCLK_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22277_ _22274_/X _22276_/X _21306_/C _24826_/Q _21082_/X VGND VGND VPWR VPWR _22277_/X
+ sky130_fd_sc_hd__a32o_4
X_25065_ _25070_/CLK _25065_/D HRESETn VGND VGND VPWR VPWR _22044_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18640__A1_N _16576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12030_ _12029_/Y _12027_/X _25488_/Q _12027_/X VGND VGND VPWR VPWR _25489_/D sky130_fd_sc_hd__a2bb2o_4
X_21228_ _21024_/X VGND VGND VPWR VPWR _21235_/A sky130_fd_sc_hd__buf_2
X_24016_ _24049_/CLK _20747_/X HRESETn VGND VGND VPWR VPWR _13121_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_144_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15735__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21159_ _21159_/A VGND VGND VPWR VPWR _21159_/X sky130_fd_sc_hd__buf_2
X_13981_ _13990_/A _13978_/X _13980_/X VGND VGND VPWR VPWR _13981_/X sky130_fd_sc_hd__or3_4
XFILLER_93_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15720_ _15540_/X _15709_/X _15719_/X _24881_/Q _15707_/X VGND VGND VPWR VPWR _15720_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_86_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12932_ _12834_/A _12756_/X _12834_/C _12931_/X VGND VGND VPWR VPWR _12932_/X sky130_fd_sc_hd__or4_4
X_24918_ _24508_/CLK _15571_/X HRESETn VGND VGND VPWR VPWR _24918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24843__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15651_ _15651_/A VGND VGND VPWR VPWR _15651_/X sky130_fd_sc_hd__buf_2
XFILLER_206_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12863_ _12857_/A _12851_/X _12862_/X _12859_/B VGND VGND VPWR VPWR _12864_/A sky130_fd_sc_hd__a211o_4
X_24849_ _25341_/CLK _24849_/D HRESETn VGND VGND VPWR VPWR _24849_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16566__A _16566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22306__A2 _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _25081_/Q VGND VGND VPWR VPWR _14602_/Y sky130_fd_sc_hd__inv_2
XPHY_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _11814_/A VGND VGND VPWR VPWR _11814_/Y sky130_fd_sc_hd__inv_2
X_18370_ _18369_/Y _18357_/Y _18354_/A _18356_/X VGND VGND VPWR VPWR _24199_/D sky130_fd_sc_hd__o22a_4
XPHY_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15580_/Y _15576_/X _15581_/X _15576_/X VGND VGND VPWR VPWR _24914_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12255__B1 _12254_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12793_/Y VGND VGND VPWR VPWR _22667_/A sky130_fd_sc_hd__buf_2
XANTENNA__20088__A _20088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17318_/B VGND VGND VPWR VPWR _17322_/B sky130_fd_sc_hd__inv_2
XPHY_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _13999_/X VGND VGND VPWR VPWR _14534_/C sky130_fd_sc_hd__inv_2
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11741_/Y _11733_/X _11743_/X _11744_/X VGND VGND VPWR VPWR _11745_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_214_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17245_/Y _17246_/Y _17249_/X _17252_/D VGND VGND VPWR VPWR _17252_/X sky130_fd_sc_hd__or4_4
X_14464_ _14461_/Y _14463_/X _14400_/X _14463_/X VGND VGND VPWR VPWR _25121_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23267__B1 _12316_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _11676_/A _11676_/B VGND VGND VPWR VPWR _11700_/A sky130_fd_sc_hd__or2_4
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ _16190_/X VGND VGND VPWR VPWR _16203_/X sky130_fd_sc_hd__buf_2
X_13415_ _13314_/X _13415_/B _13414_/X VGND VGND VPWR VPWR _13416_/C sky130_fd_sc_hd__and3_4
X_17183_ _23078_/A VGND VGND VPWR VPWR _17183_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14395_ _14395_/A _14425_/B VGND VGND VPWR VPWR _14395_/X sky130_fd_sc_hd__or2_4
X_16134_ _16133_/Y _16129_/X _11743_/X _16129_/X VGND VGND VPWR VPWR _16134_/X sky130_fd_sc_hd__a2bb2o_4
X_13346_ _13220_/X _13346_/B VGND VGND VPWR VPWR _13346_/X sky130_fd_sc_hd__or2_4
XFILLER_154_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18608__A1_N _16578_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16065_ _15988_/X VGND VGND VPWR VPWR _16065_/X sky130_fd_sc_hd__buf_2
X_13277_ _13167_/A _19745_/A VGND VGND VPWR VPWR _13277_/X sky130_fd_sc_hd__or2_4
XFILLER_108_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22750__B _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15016_ _15009_/X _15011_/X _15016_/C _15015_/X VGND VGND VPWR VPWR _15017_/D sky130_fd_sc_hd__or4_4
X_12228_ _12228_/A _12228_/B _12224_/X _12227_/X VGND VGND VPWR VPWR _12228_/X sky130_fd_sc_hd__or4_4
XFILLER_170_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19824_ _19824_/A VGND VGND VPWR VPWR _19824_/X sky130_fd_sc_hd__buf_2
X_12159_ _12159_/A VGND VGND VPWR VPWR SSn_S3 sky130_fd_sc_hd__inv_2
XFILLER_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19755_ _19753_/Y _19754_/X _19708_/X _19754_/X VGND VGND VPWR VPWR _23629_/D sky130_fd_sc_hd__a2bb2o_4
X_16967_ _16073_/Y _17040_/A _16073_/Y _17040_/A VGND VGND VPWR VPWR _16967_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22545__A2 _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18706_ _18706_/A _18705_/X VGND VGND VPWR VPWR _18707_/C sky130_fd_sc_hd__or2_4
XFILLER_209_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15918_ _15773_/B _15918_/B VGND VGND VPWR VPWR _15918_/X sky130_fd_sc_hd__or2_4
XFILLER_37_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24584__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16898_ _24285_/Q VGND VGND VPWR VPWR _16898_/Y sky130_fd_sc_hd__inv_2
X_19686_ _19684_/Y _19685_/X _19540_/X _19685_/X VGND VGND VPWR VPWR _19686_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22478__A _21080_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15849_ _15958_/A VGND VGND VPWR VPWR _15850_/A sky130_fd_sc_hd__buf_2
X_18637_ _18637_/A _18637_/B _18634_/X _18637_/D VGND VGND VPWR VPWR _18637_/X sky130_fd_sc_hd__or4_4
XFILLER_224_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24513__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_111_0_HCLK clkbuf_7_55_0_HCLK/X VGND VGND VPWR VPWR _24903_/CLK sky130_fd_sc_hd__clkbuf_1
X_18568_ _18400_/Y _18567_/X VGND VGND VPWR VPWR _18568_/X sky130_fd_sc_hd__or2_4
XFILLER_220_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_174_0_HCLK clkbuf_7_87_0_HCLK/X VGND VGND VPWR VPWR _23831_/CLK sky130_fd_sc_hd__clkbuf_1
X_17519_ _24300_/Q VGND VGND VPWR VPWR _17519_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18499_ _18499_/A _18499_/B _18505_/A _18498_/X VGND VGND VPWR VPWR _18499_/X sky130_fd_sc_hd__or4_4
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20530_ _24074_/Q _20535_/B _20518_/X VGND VGND VPWR VPWR _20530_/X sky130_fd_sc_hd__a21o_4
XANTENNA__12549__B2 _12551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20461_ _20461_/A _20459_/Y VGND VGND VPWR VPWR _24086_/D sky130_fd_sc_hd__or2_4
XFILLER_165_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22200_ _22226_/A _22200_/B _22200_/C VGND VGND VPWR VPWR _22205_/B sky130_fd_sc_hd__and3_4
XANTENNA__25372__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23180_ _24440_/Q _23138_/X _23001_/X _23179_/X VGND VGND VPWR VPWR _23181_/C sky130_fd_sc_hd__a211o_4
XANTENNA__17488__B2 _17487_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20392_ _20391_/Y _20389_/X _19743_/X _20389_/X VGND VGND VPWR VPWR _23391_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15527__A2_N _15524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22131_ _22129_/X _22130_/X _21541_/X _12551_/A _21542_/X VGND VGND VPWR VPWR _22131_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22062_ _21250_/A VGND VGND VPWR VPWR _22365_/A sky130_fd_sc_hd__buf_2
XFILLER_245_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21013_ _21013_/A _21013_/B VGND VGND VPWR VPWR _21013_/X sky130_fd_sc_hd__and2_4
XFILLER_102_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16999__B1 _16035_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19937__B1 _19874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17770__A _23320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22964_ _22959_/Y _22963_/Y _22854_/X VGND VGND VPWR VPWR _22965_/D sky130_fd_sc_hd__o21a_4
XFILLER_244_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24703_ _24753_/CLK _24703_/D HRESETn VGND VGND VPWR VPWR _24703_/Q sky130_fd_sc_hd__dfrtp_4
X_21915_ _21911_/X _21914_/X _22212_/A VGND VGND VPWR VPWR _21915_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22819__C _22818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_70_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_70_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22895_ _23072_/A _22882_/Y _22895_/C _22895_/D VGND VGND VPWR VPWR _22895_/X sky130_fd_sc_hd__or4_4
XANTENNA__16386__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24634_ _24634_/CLK _24634_/D HRESETn VGND VGND VPWR VPWR _16303_/A sky130_fd_sc_hd__dfrtp_4
X_21846_ _21846_/A _14246_/A VGND VGND VPWR VPWR _21851_/A sky130_fd_sc_hd__or2_4
XFILLER_243_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15974__A1 _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15974__B2 _15925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12788__B2 _24797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24565_ _24540_/CLK _24565_/D HRESETn VGND VGND VPWR VPWR _24565_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21777_ _22380_/A _21777_/B _21777_/C VGND VGND VPWR VPWR _21777_/X sky130_fd_sc_hd__and3_4
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23516_ _23388_/CLK _23516_/D VGND VGND VPWR VPWR _13399_/B sky130_fd_sc_hd__dfxtp_4
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20728_ _20727_/Y _20723_/X _13117_/X VGND VGND VPWR VPWR _20728_/X sky130_fd_sc_hd__o21a_4
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24496_ _24427_/CLK _16676_/X HRESETn VGND VGND VPWR VPWR _24496_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23447_ _23808_/CLK _23447_/D VGND VGND VPWR VPWR _23447_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20659_ _20659_/A VGND VGND VPWR VPWR _20659_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ _13200_/A _20224_/A VGND VGND VPWR VPWR _13201_/C sky130_fd_sc_hd__or2_4
X_14180_ _14180_/A _12043_/Y _11668_/B _13765_/A VGND VGND VPWR VPWR _14181_/A sky130_fd_sc_hd__or4_4
XANTENNA__21275__A2 _21273_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23378_ _23378_/CLK _20425_/X VGND VGND VPWR VPWR _20424_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_136_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25042__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13131_ _13284_/A VGND VGND VPWR VPWR _13263_/A sky130_fd_sc_hd__buf_2
X_25117_ _25117_/CLK _25117_/D HRESETn VGND VGND VPWR VPWR _25117_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22329_ _22328_/X VGND VGND VPWR VPWR _22329_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13062_ _12340_/A _13062_/B VGND VGND VPWR VPWR _13064_/B sky130_fd_sc_hd__or2_4
X_25048_ _25050_/CLK _14849_/X HRESETn VGND VGND VPWR VPWR _14810_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20235__B1 _20061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12013_ _13513_/B _12013_/B _12013_/C _14278_/A VGND VGND VPWR VPWR _12014_/A sky130_fd_sc_hd__or4_4
XFILLER_151_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17870_ _16889_/Y _17873_/B VGND VGND VPWR VPWR _17874_/B sky130_fd_sc_hd__or2_4
XANTENNA__17100__B1 _17053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16821_ _16793_/A VGND VGND VPWR VPWR _16841_/A sky130_fd_sc_hd__buf_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16752_ _16751_/Y _16749_/X _16400_/X _16749_/X VGND VGND VPWR VPWR _24464_/D sky130_fd_sc_hd__a2bb2o_4
X_19540_ _11785_/A VGND VGND VPWR VPWR _19540_/X sky130_fd_sc_hd__buf_2
X_13964_ _14028_/A VGND VGND VPWR VPWR _13995_/A sky130_fd_sc_hd__buf_2
X_15703_ _11678_/X VGND VGND VPWR VPWR _15704_/A sky130_fd_sc_hd__buf_2
X_12915_ _12801_/X _12912_/X VGND VGND VPWR VPWR _12915_/X sky130_fd_sc_hd__or2_4
X_16683_ _16682_/Y _16680_/X _15741_/X _16680_/X VGND VGND VPWR VPWR _16683_/X sky130_fd_sc_hd__a2bb2o_4
X_19471_ _19469_/Y _19470_/X _11924_/X _19470_/X VGND VGND VPWR VPWR _19471_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25136__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13895_ _13892_/A _13935_/B _13943_/A _13894_/B VGND VGND VPWR VPWR _13895_/X sky130_fd_sc_hd__or4_4
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15634_ _15634_/A VGND VGND VPWR VPWR _21124_/A sky130_fd_sc_hd__inv_2
X_18422_ _24176_/Q VGND VGND VPWR VPWR _18467_/A sky130_fd_sc_hd__inv_2
XFILLER_64_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25199__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12846_ _12848_/B VGND VGND VPWR VPWR _12847_/B sky130_fd_sc_hd__inv_2
X_18353_ _18352_/Y _17476_/A _21979_/A _17480_/X VGND VGND VPWR VPWR _18353_/X sky130_fd_sc_hd__o22a_4
XFILLER_159_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15565_ _15563_/Y _15561_/X _15564_/X _15561_/X VGND VGND VPWR VPWR _15565_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_203_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16446__D _16446_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_247_0_HCLK clkbuf_8_247_0_HCLK/A VGND VGND VPWR VPWR _24967_/CLK sky130_fd_sc_hd__clkbuf_1
X_12777_ _25370_/Q _24787_/Q _12775_/Y _12776_/Y VGND VGND VPWR VPWR _12778_/D sky130_fd_sc_hd__o22a_4
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23977__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17304_ _17245_/Y _17246_/Y _17343_/B _17244_/X VGND VGND VPWR VPWR _17304_/X sky130_fd_sc_hd__or4_4
XFILLER_30_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14510_/X _14515_/X _25117_/Q _14506_/X VGND VGND VPWR VPWR _25105_/D sky130_fd_sc_hd__o22a_4
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _25535_/Q VGND VGND VPWR VPWR _11728_/Y sky130_fd_sc_hd__inv_2
X_18284_ _17711_/Y _18283_/X _18288_/A VGND VGND VPWR VPWR _18284_/X sky130_fd_sc_hd__or3_4
X_15496_ _15496_/A VGND VGND VPWR VPWR _15496_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12571__A2_N _24859_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17235_ _17292_/A VGND VGND VPWR VPWR _17236_/A sky130_fd_sc_hd__inv_2
XFILLER_202_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14447_ _14447_/A VGND VGND VPWR VPWR _14447_/Y sky130_fd_sc_hd__inv_2
X_11659_ _11659_/A VGND VGND VPWR VPWR _11660_/A sky130_fd_sc_hd__buf_2
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17166_ _17165_/Y VGND VGND VPWR VPWR _17366_/A sky130_fd_sc_hd__buf_2
XANTENNA__18667__B1 _16613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22463__A1 _22696_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14378_ _20462_/A _14371_/X _13829_/X _14373_/X VGND VGND VPWR VPWR _14378_/X sky130_fd_sc_hd__a2bb2o_4
X_16117_ _16115_/Y _16111_/X _15948_/X _16116_/X VGND VGND VPWR VPWR _24700_/D sky130_fd_sc_hd__a2bb2o_4
X_13329_ _13393_/A _13329_/B _13328_/X VGND VGND VPWR VPWR _13329_/X sky130_fd_sc_hd__and3_4
X_17097_ _17030_/D _17097_/B VGND VGND VPWR VPWR _17098_/B sky130_fd_sc_hd__or2_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16048_ _16047_/Y _16045_/X _15965_/X _16045_/X VGND VGND VPWR VPWR _16048_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24765__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19807_ _16854_/X VGND VGND VPWR VPWR _19807_/X sky130_fd_sc_hd__buf_2
XFILLER_85_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24338__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17999_ _17999_/A VGND VGND VPWR VPWR _18118_/A sky130_fd_sc_hd__buf_2
X_19738_ _19273_/A _18911_/B _19047_/C VGND VGND VPWR VPWR _19738_/X sky130_fd_sc_hd__or3_4
XFILLER_226_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19669_ _19668_/Y _19664_/X _19646_/X _19650_/Y VGND VGND VPWR VPWR _19669_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_57_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21700_ _21525_/A _21700_/B VGND VGND VPWR VPWR _21700_/X sky130_fd_sc_hd__and2_4
XFILLER_198_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13623__A _13622_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22680_ _11844_/Y _21956_/A _13556_/Y _22515_/A VGND VGND VPWR VPWR _22680_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21631_ _22380_/A _21631_/B _21631_/C VGND VGND VPWR VPWR _21631_/X sky130_fd_sc_hd__and3_4
XFILLER_100_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22151__B1 _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24350_ _24667_/CLK _17359_/X HRESETn VGND VGND VPWR VPWR _24350_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15708__A1 _15540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21562_ _14198_/Y _14182_/X _14224_/Y _14209_/X VGND VGND VPWR VPWR _21563_/A sky130_fd_sc_hd__o22a_4
XANTENNA__16905__B1 _16144_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23301_ _24610_/Q _23301_/B VGND VGND VPWR VPWR _23304_/B sky130_fd_sc_hd__or2_4
X_20513_ _24076_/Q _20512_/Y VGND VGND VPWR VPWR _20514_/C sky130_fd_sc_hd__and2_4
XFILLER_21_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21493_ _21484_/X _21493_/B _21493_/C VGND VGND VPWR VPWR _21493_/X sky130_fd_sc_hd__and3_4
X_24281_ _24275_/CLK _24281_/D HRESETn VGND VGND VPWR VPWR _17744_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_147_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20444_ _20444_/A _20444_/B VGND VGND VPWR VPWR _20444_/X sky130_fd_sc_hd__and2_4
X_23232_ _16647_/Y _23291_/B VGND VGND VPWR VPWR _23232_/X sky130_fd_sc_hd__and2_4
XFILLER_107_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20375_ _20369_/X VGND VGND VPWR VPWR _20375_/Y sky130_fd_sc_hd__inv_2
X_23163_ _23161_/X _23162_/X _22919_/X VGND VGND VPWR VPWR _23163_/X sky130_fd_sc_hd__or3_4
X_22114_ _12217_/Y _15780_/B _16925_/Y _21447_/X VGND VGND VPWR VPWR _22114_/X sky130_fd_sc_hd__o22a_4
X_23094_ _23094_/A _23093_/X VGND VGND VPWR VPWR _23094_/Y sky130_fd_sc_hd__nor2_4
XFILLER_122_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22045_ _14720_/A _19589_/Y _22042_/X _22044_/X VGND VGND VPWR VPWR _22045_/X sky130_fd_sc_hd__o22a_4
XFILLER_121_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19980__A _19962_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23996_ _24080_/CLK _23996_/D HRESETn VGND VGND VPWR VPWR _13839_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_216_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22947_ _12813_/Y _21446_/X _16938_/Y _22826_/X VGND VGND VPWR VPWR _22947_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22390__B1 _14710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12700_ _12697_/A _12697_/B VGND VGND VPWR VPWR _12701_/C sky130_fd_sc_hd__nand2_4
XFILLER_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13680_ _11806_/A _13692_/B _11843_/A _11820_/A VGND VGND VPWR VPWR _13680_/X sky130_fd_sc_hd__and4_4
XFILLER_71_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22878_ _22878_/A _22989_/B VGND VGND VPWR VPWR _22878_/X sky130_fd_sc_hd__and2_4
XFILLER_232_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12631_ _12633_/B VGND VGND VPWR VPWR _12632_/B sky130_fd_sc_hd__inv_2
X_24617_ _24618_/CLK _16347_/X HRESETn VGND VGND VPWR VPWR _24617_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21829_ _21714_/X _21751_/X _21790_/X _21828_/X VGND VGND VPWR VPWR HRDATA[3] sky130_fd_sc_hd__or4_4
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22142__B1 _23328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16844__A _24418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ _24997_/Q _15349_/Y VGND VGND VPWR VPWR _15350_/X sky130_fd_sc_hd__or2_4
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_0_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_12562_ _25418_/Q VGND VGND VPWR VPWR _12671_/A sky130_fd_sc_hd__inv_2
X_24548_ _24520_/CLK _16535_/X HRESETn VGND VGND VPWR VPWR _16534_/A sky130_fd_sc_hd__dfrtp_4
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22693__A1 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22693__B2 _22692_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_14_0_HCLK clkbuf_7_7_0_HCLK/X VGND VGND VPWR VPWR _23575_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14301_ _14295_/X _14299_/X _13466_/A _14300_/X VGND VGND VPWR VPWR _25177_/D sky130_fd_sc_hd__o22a_4
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ _15281_/A VGND VGND VPWR VPWR _15282_/B sky130_fd_sc_hd__inv_2
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12263_/A _12493_/B _12493_/C VGND VGND VPWR VPWR _25434_/D sky130_fd_sc_hd__and3_4
X_24479_ _24900_/CLK _24479_/D HRESETn VGND VGND VPWR VPWR _24479_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14364__A _14364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_77_0_HCLK clkbuf_8_77_0_HCLK/A VGND VGND VPWR VPWR _24753_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17020_ _24645_/Q VGND VGND VPWR VPWR _17020_/Y sky130_fd_sc_hd__inv_2
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _13927_/A _14232_/B _14232_/C _14231_/Y VGND VGND VPWR VPWR _14233_/B sky130_fd_sc_hd__and4_4
XFILLER_50_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15179__B _15311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22581__A _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14163_ _14159_/Y _14162_/Y _14154_/X VGND VGND VPWR VPWR _14163_/X sky130_fd_sc_hd__o21a_4
XFILLER_124_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13114_ _13114_/A _13113_/X VGND VGND VPWR VPWR _20704_/A sky130_fd_sc_hd__or2_4
XFILLER_98_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14094_ _14094_/A VGND VGND VPWR VPWR _14094_/Y sky130_fd_sc_hd__inv_2
X_18971_ _18970_/Y _18966_/X _18951_/X _18966_/X VGND VGND VPWR VPWR _18971_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15883__B1 _24800_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13045_ _12291_/X _13051_/B VGND VGND VPWR VPWR _13046_/B sky130_fd_sc_hd__or2_4
X_17922_ _24250_/Q VGND VGND VPWR VPWR _17926_/A sky130_fd_sc_hd__inv_2
XFILLER_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17853_ _16908_/Y _16889_/Y _16925_/Y _17853_/D VGND VGND VPWR VPWR _17862_/B sky130_fd_sc_hd__or4_4
XANTENNA__15635__B1 _15475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16804_ _16799_/A VGND VGND VPWR VPWR _16804_/X sky130_fd_sc_hd__buf_2
XANTENNA__15923__A _15783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24105__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14996_ _14995_/X _16743_/A _14995_/X _16743_/A VGND VGND VPWR VPWR _14996_/X sky130_fd_sc_hd__a2bb2o_4
X_17784_ _16945_/X _17775_/C _17783_/X _17780_/B VGND VGND VPWR VPWR _17784_/X sky130_fd_sc_hd__a211o_4
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19523_ _21215_/A VGND VGND VPWR VPWR _19523_/Y sky130_fd_sc_hd__inv_2
X_13947_ _13947_/A _13947_/B _13947_/C _13879_/X VGND VGND VPWR VPWR _13947_/X sky130_fd_sc_hd__or4_4
X_16735_ _16730_/A VGND VGND VPWR VPWR _16735_/X sky130_fd_sc_hd__buf_2
XFILLER_235_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16666_ _16665_/Y _16661_/X _16483_/X _16661_/X VGND VGND VPWR VPWR _16666_/X sky130_fd_sc_hd__a2bb2o_4
X_19454_ _18285_/B VGND VGND VPWR VPWR _19939_/B sky130_fd_sc_hd__buf_2
X_13878_ _13908_/A _13878_/B _13930_/A _13932_/C VGND VGND VPWR VPWR _13879_/C sky130_fd_sc_hd__or4_4
XFILLER_179_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22756__A _16679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16060__B1 _16059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15617_ _15615_/Y _15613_/X _15616_/X _15613_/X VGND VGND VPWR VPWR _15617_/X sky130_fd_sc_hd__a2bb2o_4
X_18405_ _16265_/Y _24158_/Q _16265_/Y _24158_/Q VGND VGND VPWR VPWR _18406_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12829_ _12879_/A _12759_/Y VGND VGND VPWR VPWR _12841_/C sky130_fd_sc_hd__or2_4
XFILLER_50_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16597_ HWDATA[9] VGND VGND VPWR VPWR _16597_/X sky130_fd_sc_hd__buf_2
X_19385_ _19384_/Y _19380_/X _19295_/X _19372_/A VGND VGND VPWR VPWR _19385_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_222_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12059__A _12058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15548_ _15540_/X _15544_/Y _15545_/X _23324_/A _15550_/A VGND VGND VPWR VPWR _15548_/X
+ sky130_fd_sc_hd__a32o_4
X_18336_ _18336_/A _17448_/A VGND VGND VPWR VPWR _20220_/B sky130_fd_sc_hd__or2_4
XFILLER_188_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11898__A _11897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18267_ _13783_/D _18256_/X _18257_/X _24224_/Q _18264_/X VGND VGND VPWR VPWR _18267_/X
+ sky130_fd_sc_hd__a32o_4
X_15479_ _24069_/Q _15478_/Y VGND VGND VPWR VPWR _24069_/D sky130_fd_sc_hd__nor2_4
XANTENNA__17288__C _17343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17218_ _16291_/Y _24367_/Q _22944_/A _17249_/D VGND VGND VPWR VPWR _17218_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22436__A1 _16144_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14374__B1 _13824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18198_ _17966_/A _18197_/X _24243_/Q _18024_/A VGND VGND VPWR VPWR _18198_/X sky130_fd_sc_hd__o22a_4
XFILLER_190_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17149_ _17039_/Y _17126_/B _17147_/B _17064_/X VGND VGND VPWR VPWR _17149_/X sky130_fd_sc_hd__a211o_4
XFILLER_7_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24946__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17312__B1 _17276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20160_ _22387_/B _20159_/X _20089_/X _20159_/X VGND VGND VPWR VPWR _23482_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15874__B1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20091_ _23505_/Q VGND VGND VPWR VPWR _22218_/B sky130_fd_sc_hd__inv_2
XFILLER_170_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15626__B1 _15466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23850_ _23774_/CLK _23850_/D VGND VGND VPWR VPWR _23850_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22801_ _22928_/A VGND VGND VPWR VPWR _22801_/X sky130_fd_sc_hd__buf_2
XFILLER_226_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23781_ _24252_/CLK _23781_/D VGND VGND VPWR VPWR _18138_/B sky130_fd_sc_hd__dfxtp_4
X_20993_ sda_oen_o_S4 _25099_/Q _20987_/A _14026_/X _20992_/Y VGND VGND VPWR VPWR
+ _23929_/D sky130_fd_sc_hd__a32o_4
XFILLER_38_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25520_ _24357_/CLK _11795_/X HRESETn VGND VGND VPWR VPWR _25520_/Q sky130_fd_sc_hd__dfrtp_4
X_22732_ _24429_/Q _22730_/X _22533_/X _22731_/X VGND VGND VPWR VPWR _22732_/X sky130_fd_sc_hd__a211o_4
XFILLER_214_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16051__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25451_ _24766_/CLK _12434_/X HRESETn VGND VGND VPWR VPWR _12187_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_41_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22663_ _16539_/A _22662_/X _22138_/C _11737_/A _21833_/X VGND VGND VPWR VPWR _22663_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_213_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22124__B1 _23962_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24402_ _24377_/CLK _24402_/D HRESETn VGND VGND VPWR VPWR _16978_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21614_ _21609_/X _21614_/B VGND VGND VPWR VPWR _21614_/X sky130_fd_sc_hd__or2_4
XFILLER_240_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25382_ _25382_/CLK _25382_/D HRESETn VGND VGND VPWR VPWR _22713_/A sky130_fd_sc_hd__dfrtp_4
X_22594_ _24796_/Q _22630_/B VGND VGND VPWR VPWR _22594_/X sky130_fd_sc_hd__or2_4
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17479__B _17448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_230_0_HCLK clkbuf_8_231_0_HCLK/A VGND VGND VPWR VPWR _24953_/CLK sky130_fd_sc_hd__clkbuf_1
X_24333_ _24958_/CLK _17416_/X HRESETn VGND VGND VPWR VPWR _20667_/A sky130_fd_sc_hd__dfrtp_4
X_21545_ _12211_/Y _21531_/X _16917_/A _21431_/X VGND VGND VPWR VPWR _21545_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17551__B1 _11772_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24264_ _24686_/CLK _17874_/X HRESETn VGND VGND VPWR VPWR _22190_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21476_ _21472_/X _21475_/X _18301_/X VGND VGND VPWR VPWR _21477_/C sky130_fd_sc_hd__o21a_4
XFILLER_153_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23215_ _23196_/X _23199_/X _23203_/Y _23214_/X VGND VGND VPWR VPWR HRDATA[27] sky130_fd_sc_hd__a211o_4
XFILLER_181_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20427_ _21253_/B _20422_/X _19852_/A _20409_/Y VGND VGND VPWR VPWR _20427_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24195_ _25471_/CLK _24195_/D HRESETn VGND VGND VPWR VPWR _24195_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24687__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23146_ _23035_/X _23144_/X _23145_/X _24846_/Q _23037_/X VGND VGND VPWR VPWR _23146_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_122_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20358_ _21940_/B _20355_/X _19610_/A _20355_/X VGND VGND VPWR VPWR _20358_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24616__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16717__A2_N _16655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20289_ _22358_/B _20288_/X _19964_/X _20288_/X VGND VGND VPWR VPWR _23433_/D sky130_fd_sc_hd__a2bb2o_4
X_23077_ _23251_/A _23074_/X _23076_/X VGND VGND VPWR VPWR _23077_/X sky130_fd_sc_hd__and3_4
XFILLER_103_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22028_ _22021_/A _22026_/X _22027_/X VGND VGND VPWR VPWR _22028_/X sky130_fd_sc_hd__and3_4
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15617__B1 _15616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14850_ _25047_/Q _14795_/B _25047_/Q _14795_/B VGND VGND VPWR VPWR _14850_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15743__A HWDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13801_ _11668_/A _13800_/X VGND VGND VPWR VPWR _14442_/A sky130_fd_sc_hd__or2_4
XANTENNA__16290__B1 _16004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14781_ _17983_/A VGND VGND VPWR VPWR _18052_/A sky130_fd_sc_hd__buf_2
X_11993_ _13492_/A _11992_/Y _13492_/A _11992_/Y VGND VGND VPWR VPWR _11993_/X sky130_fd_sc_hd__a2bb2o_4
X_23979_ _23986_/CLK _20637_/Y HRESETn VGND VGND VPWR VPWR _17388_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16520_ _16520_/A VGND VGND VPWR VPWR _16520_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13732_ _13731_/X VGND VGND VPWR VPWR _13732_/X sky130_fd_sc_hd__buf_2
XANTENNA__25475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20913__A1 _16670_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_40_0_HCLK clkbuf_6_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_81_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16451_ _15855_/B VGND VGND VPWR VPWR _16724_/A sky130_fd_sc_hd__buf_2
XANTENNA__25404__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13663_ _25296_/Q VGND VGND VPWR VPWR _13663_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15402_ _15281_/A VGND VGND VPWR VPWR _15402_/X sky130_fd_sc_hd__buf_2
XFILLER_25_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22295__B _22420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12614_ _12500_/Y _12614_/B VGND VGND VPWR VPWR _12615_/C sky130_fd_sc_hd__or2_4
X_19170_ _19170_/A VGND VGND VPWR VPWR _19170_/X sky130_fd_sc_hd__buf_2
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16382_ HWDATA[26] VGND VGND VPWR VPWR _16382_/X sky130_fd_sc_hd__buf_2
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13594_ _14628_/A _13592_/B _13593_/Y VGND VGND VPWR VPWR _13594_/X sky130_fd_sc_hd__o21a_4
XFILLER_169_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20096__A _20088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18121_ _18004_/X _18121_/B VGND VGND VPWR VPWR _18123_/B sky130_fd_sc_hd__or2_4
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15333_ _15333_/A _15333_/B VGND VGND VPWR VPWR _15338_/B sky130_fd_sc_hd__or2_4
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12545_ _12535_/X _12545_/B _12545_/C _12544_/X VGND VGND VPWR VPWR _12546_/D sky130_fd_sc_hd__or4_4
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18052_ _18052_/A VGND VGND VPWR VPWR _18099_/A sky130_fd_sc_hd__buf_2
X_15264_ _15245_/A _15266_/B _15263_/Y VGND VGND VPWR VPWR _25015_/D sky130_fd_sc_hd__o21a_4
X_12476_ _12257_/Y _12476_/B VGND VGND VPWR VPWR _12480_/B sky130_fd_sc_hd__or2_4
X_17003_ _16064_/Y _17039_/A _24744_/Q _17022_/A VGND VGND VPWR VPWR _17008_/B sky130_fd_sc_hd__a2bb2o_4
X_14215_ _14215_/A VGND VGND VPWR VPWR _14215_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23200__A _16650_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15195_ _15189_/A _15188_/X _15194_/X _15190_/Y VGND VGND VPWR VPWR _15195_/X sky130_fd_sc_hd__a211o_4
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14146_ _14118_/X _14145_/X _14428_/A _14125_/X VGND VGND VPWR VPWR _14146_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__24357__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14077_ _14005_/B _14070_/X _14058_/X _14005_/A _14073_/X VGND VGND VPWR VPWR _25229_/D
+ sky130_fd_sc_hd__a32o_4
X_18954_ _18953_/Y _18947_/X _17440_/X _18947_/A VGND VGND VPWR VPWR _23907_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13028_ _13028_/A _13024_/Y _13028_/C VGND VGND VPWR VPWR _13028_/X sky130_fd_sc_hd__or3_4
X_17905_ _21997_/A _17904_/X _21997_/A _17904_/X VGND VGND VPWR VPWR _24257_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18885_ _18885_/A VGND VGND VPWR VPWR _18885_/X sky130_fd_sc_hd__buf_2
XFILLER_67_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18270__A1 _13783_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17836_ _17757_/Y _17833_/X VGND VGND VPWR VPWR _17836_/X sky130_fd_sc_hd__or2_4
XANTENNA__19125__A _18985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_122_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_122_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17767_ _17555_/X _17766_/X VGND VGND VPWR VPWR _17768_/D sky130_fd_sc_hd__or2_4
XFILLER_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14979_ _14946_/X _14958_/X _14969_/X _14979_/D VGND VGND VPWR VPWR _14979_/X sky130_fd_sc_hd__or4_4
XANTENNA__21157__B2 _14422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18558__C1 _18489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23992__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19506_ _22236_/B _19503_/X _11906_/X _19503_/X VGND VGND VPWR VPWR _23713_/D sky130_fd_sc_hd__a2bb2o_4
X_16718_ _16365_/A VGND VGND VPWR VPWR _16719_/A sky130_fd_sc_hd__inv_2
XFILLER_34_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17698_ _17665_/D VGND VGND VPWR VPWR _17698_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22486__A _21864_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21390__A _22196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19437_ _17992_/B VGND VGND VPWR VPWR _19437_/Y sky130_fd_sc_hd__inv_2
X_16649_ _16647_/Y _16643_/X _16464_/X _16648_/X VGND VGND VPWR VPWR _16649_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13_0_HCLK_A clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19368_ _19364_/Y _19367_/X _19301_/X _19367_/X VGND VGND VPWR VPWR _23762_/D sky130_fd_sc_hd__a2bb2o_4
X_18319_ _18285_/B _18318_/X _18282_/A _18318_/X VGND VGND VPWR VPWR _18319_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19299_ _19299_/A VGND VGND VPWR VPWR _19299_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17533__B1 _11732_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21330_ _21338_/A VGND VGND VPWR VPWR _22891_/A sky130_fd_sc_hd__buf_2
XANTENNA__22409__A1 _21501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22409__B2 _22408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_60_0_HCLK clkbuf_7_30_0_HCLK/X VGND VGND VPWR VPWR _25091_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_117_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21261_ _22069_/A _21259_/X _21261_/C VGND VGND VPWR VPWR _21261_/X sky130_fd_sc_hd__and3_4
XANTENNA__23082__A1 _12759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19286__B1 _19194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24780__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23000_ _15084_/A _23177_/B VGND VGND VPWR VPWR _23000_/X sky130_fd_sc_hd__or2_4
X_20212_ _18139_/B VGND VGND VPWR VPWR _20212_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21192_ _21205_/A _21192_/B VGND VGND VPWR VPWR _21192_/X sky130_fd_sc_hd__or2_4
XFILLER_89_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24098__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20143_ _20137_/Y VGND VGND VPWR VPWR _20143_/X sky130_fd_sc_hd__buf_2
XFILLER_143_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19038__B1 _18965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24027__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20074_ _23511_/Q VGND VGND VPWR VPWR _20074_/Y sky130_fd_sc_hd__inv_2
X_24951_ _24953_/CLK _15476_/X HRESETn VGND VGND VPWR VPWR _24951_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21565__A _15662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23902_ _23884_/CLK _23902_/D VGND VGND VPWR VPWR _18114_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_245_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24882_ _24874_/CLK _15718_/X HRESETn VGND VGND VPWR VPWR _12515_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23833_ _24089_/CLK _23833_/D VGND VGND VPWR VPWR _23833_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15282__B _15282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14179__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13083__A _13085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23764_ _23767_/CLK _23764_/D VGND VGND VPWR VPWR _23764_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _12143_/X _12147_/A VGND VGND VPWR VPWR _24107_/D sky130_fd_sc_hd__and2_4
XPHY_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25503_ _23691_/CLK _25503_/D HRESETn VGND VGND VPWR VPWR _19874_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_5_27_0_HCLK clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_54_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22715_ _24869_/Q _21863_/X _21118_/X _22714_/X VGND VGND VPWR VPWR _22715_/X sky130_fd_sc_hd__a211o_4
XFILLER_198_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23695_ _23406_/CLK _23695_/D VGND VGND VPWR VPWR _23695_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25434_ _25444_/CLK _25434_/D HRESETn VGND VGND VPWR VPWR _12268_/A sky130_fd_sc_hd__dfrtp_4
X_22646_ _17756_/Y _21447_/X _12418_/B _21448_/X VGND VGND VPWR VPWR _22646_/X sky130_fd_sc_hd__o22a_4
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22648__B2 _22647_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25365_ _25387_/CLK _12999_/Y HRESETn VGND VGND VPWR VPWR _25365_/Q sky130_fd_sc_hd__dfrtp_4
X_22577_ _22539_/X _22577_/B _22577_/C _22577_/D VGND VGND VPWR VPWR HRDATA[10] sky130_fd_sc_hd__or4_4
XFILLER_194_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24868__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12330_ _25340_/Q VGND VGND VPWR VPWR _12330_/Y sky130_fd_sc_hd__inv_2
X_24316_ _24310_/CLK _17618_/X HRESETn VGND VGND VPWR VPWR _17564_/A sky130_fd_sc_hd__dfrtp_4
X_21528_ _24787_/Q _21528_/B VGND VGND VPWR VPWR _21528_/X sky130_fd_sc_hd__or2_4
X_25296_ _24233_/CLK _25296_/D HRESETn VGND VGND VPWR VPWR _25296_/Q sky130_fd_sc_hd__dfrtp_4
X_12261_ _12261_/A _12261_/B VGND VGND VPWR VPWR _12261_/X sky130_fd_sc_hd__or2_4
X_24247_ _23774_/CLK _18064_/X HRESETn VGND VGND VPWR VPWR _24247_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19277__B1 _19144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21459_ _21817_/A _20281_/Y VGND VGND VPWR VPWR _21459_/X sky130_fd_sc_hd__or2_4
XFILLER_135_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14000_ _13978_/X VGND VGND VPWR VPWR _14000_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24450__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12192_ _24756_/Q VGND VGND VPWR VPWR _12192_/Y sky130_fd_sc_hd__inv_2
X_24178_ _24675_/CLK _18532_/Y HRESETn VGND VGND VPWR VPWR _24178_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15457__B _14212_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23129_ _23129_/A VGND VGND VPWR VPWR _23169_/A sky130_fd_sc_hd__buf_2
XFILLER_1_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19029__B1 _19006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15951_ HWDATA[18] VGND VGND VPWR VPWR _15951_/X sky130_fd_sc_hd__buf_2
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16569__A _16569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14902_ _14902_/A VGND VGND VPWR VPWR _15056_/D sky130_fd_sc_hd__inv_2
X_15882_ _15879_/X _15880_/X _15735_/X _24801_/Q _15881_/X VGND VGND VPWR VPWR _15882_/X
+ sky130_fd_sc_hd__a32o_4
X_18670_ _18638_/X _18670_/B VGND VGND VPWR VPWR _18705_/B sky130_fd_sc_hd__or2_4
X_17621_ _17615_/B VGND VGND VPWR VPWR _17621_/Y sky130_fd_sc_hd__inv_2
X_14833_ _25052_/Q _14811_/X _25052_/Q _14811_/X VGND VGND VPWR VPWR _14833_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21139__B2 _21348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14764_ _14764_/A VGND VGND VPWR VPWR _14764_/X sky130_fd_sc_hd__buf_2
X_17552_ _11763_/Y _24297_/Q _11777_/Y _24294_/Q VGND VGND VPWR VPWR _17553_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19201__B1 _19200_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11976_ _11976_/A VGND VGND VPWR VPWR _11976_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16015__B1 _11691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13715_ _13670_/X _13714_/Y _13708_/X _13700_/X _11816_/A VGND VGND VPWR VPWR _25284_/D
+ sky130_fd_sc_hd__a32o_4
X_16503_ _24560_/Q VGND VGND VPWR VPWR _16503_/Y sky130_fd_sc_hd__inv_2
X_17483_ _17453_/X _17482_/A _17455_/Y _17482_/Y VGND VGND VPWR VPWR _17483_/X sky130_fd_sc_hd__o22a_4
X_14695_ _20157_/C _14673_/A _13723_/A _14741_/A VGND VGND VPWR VPWR _14695_/X sky130_fd_sc_hd__o22a_4
XFILLER_232_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19222_ _19220_/Y _19216_/X _19221_/X _19216_/X VGND VGND VPWR VPWR _19222_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_232_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13646_ _24042_/Q _20857_/B _24044_/Q _24043_/Q VGND VGND VPWR VPWR _13647_/B sky130_fd_sc_hd__or4_4
X_16434_ HWDATA[2] VGND VGND VPWR VPWR _19063_/A sky130_fd_sc_hd__buf_2
XFILLER_232_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16365_ _16365_/A VGND VGND VPWR VPWR _16366_/B sky130_fd_sc_hd__buf_2
X_19153_ _18126_/B VGND VGND VPWR VPWR _19153_/Y sky130_fd_sc_hd__inv_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13577_ _15904_/B _13577_/B VGND VGND VPWR VPWR _15694_/A sky130_fd_sc_hd__and2_4
XFILLER_9_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22753__B _22638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15316_ _15315_/X VGND VGND VPWR VPWR _15316_/Y sky130_fd_sc_hd__inv_2
X_18104_ _18104_/A _19376_/A VGND VGND VPWR VPWR _18104_/X sky130_fd_sc_hd__or2_4
X_12528_ _12526_/A _24879_/Q _12644_/A _12527_/Y VGND VGND VPWR VPWR _12528_/X sky130_fd_sc_hd__o22a_4
X_16296_ _16294_/Y _16292_/X _16295_/X _16292_/X VGND VGND VPWR VPWR _24637_/D sky130_fd_sc_hd__a2bb2o_4
X_19084_ _21760_/B _19079_/X _16878_/X _19079_/X VGND VGND VPWR VPWR _19084_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24538__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_47_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15247_ _15247_/A VGND VGND VPWR VPWR _15248_/B sky130_fd_sc_hd__inv_2
X_18035_ _18220_/A _18035_/B _18034_/X VGND VGND VPWR VPWR _18043_/B sky130_fd_sc_hd__or3_4
XFILLER_117_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12459_ _12197_/Y _12257_/Y _12217_/Y _12475_/B VGND VGND VPWR VPWR _12459_/X sky130_fd_sc_hd__or4_4
XFILLER_160_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15178_ _15177_/X VGND VGND VPWR VPWR _25036_/D sky130_fd_sc_hd__inv_2
XFILLER_207_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24191__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14129_ _14128_/X VGND VGND VPWR VPWR _14129_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13168__A _13168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19986_ _19986_/A VGND VGND VPWR VPWR _21185_/B sky130_fd_sc_hd__inv_2
X_18937_ _18936_/Y _18934_/X _17418_/X _18934_/X VGND VGND VPWR VPWR _18937_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25397__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18868_ _18825_/Y _18724_/X _18846_/X _18867_/X VGND VGND VPWR VPWR _18868_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25326__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17819_ _16938_/Y _17814_/B _17783_/X _17816_/B VGND VGND VPWR VPWR _17819_/X sky130_fd_sc_hd__a211o_4
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18799_ _24135_/Q _18798_/Y VGND VGND VPWR VPWR _18801_/B sky130_fd_sc_hd__or2_4
XFILLER_227_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20830_ _20830_/A VGND VGND VPWR VPWR _20830_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20761_ _20759_/Y _20755_/Y _20760_/X VGND VGND VPWR VPWR _20761_/X sky130_fd_sc_hd__o21a_4
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22500_ _12208_/X _22499_/X _16915_/A _21056_/X VGND VGND VPWR VPWR _22500_/X sky130_fd_sc_hd__a2bb2o_4
X_23480_ _23490_/CLK _23480_/D VGND VGND VPWR VPWR _20163_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_196_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20692_ _20692_/A VGND VGND VPWR VPWR _24003_/D sky130_fd_sc_hd__inv_2
XFILLER_195_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22431_ _23172_/A VGND VGND VPWR VPWR _22431_/X sky130_fd_sc_hd__buf_2
XFILLER_176_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24961__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25150_ _23926_/CLK _14381_/X HRESETn VGND VGND VPWR VPWR _20467_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22362_ _17725_/A _22361_/X _17730_/X VGND VGND VPWR VPWR _22362_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21853__A2 _12086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24279__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24101_ _25109_/CLK _20970_/Y HRESETn VGND VGND VPWR VPWR _24101_/Q sky130_fd_sc_hd__dfrtp_4
X_21313_ _21305_/B _21310_/X _21312_/X _24717_/Q _22523_/B VGND VGND VPWR VPWR _21313_/X
+ sky130_fd_sc_hd__a32o_4
X_25081_ _25081_/CLK _25081_/D HRESETn VGND VGND VPWR VPWR _25081_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24208__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22293_ _21748_/A _22293_/B VGND VGND VPWR VPWR _22293_/Y sky130_fd_sc_hd__nor2_4
XFILLER_190_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24032_ _24032_/CLK _20816_/X HRESETn VGND VGND VPWR VPWR _13125_/A sky130_fd_sc_hd__dfrtp_4
X_21244_ _21239_/A VGND VGND VPWR VPWR _21250_/A sky130_fd_sc_hd__buf_2
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_4_0_HCLK clkbuf_5_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21175_ _21175_/A _21175_/B _21175_/C VGND VGND VPWR VPWR _21224_/C sky130_fd_sc_hd__and3_4
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16493__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20126_ _21778_/B _20121_/X _20102_/X _20121_/X VGND VGND VPWR VPWR _23494_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16389__A _24603_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20057_ _20053_/X _18328_/X _13826_/A _13214_/B _20055_/X VGND VGND VPWR VPWR _20057_/X
+ sky130_fd_sc_hd__a32o_4
X_24934_ _25510_/CLK _24934_/D HRESETn VGND VGND VPWR VPWR _15518_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11857__A1 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19431__B1 _19408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25067__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24865_ _24834_/CLK _24865_/D HRESETn VGND VGND VPWR VPWR _12511_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _24227_/Q VGND VGND VPWR VPWR _11830_/Y sky130_fd_sc_hd__inv_2
X_23816_ _23873_/CLK _23816_/D VGND VGND VPWR VPWR _23816_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24796_ _24886_/CLK _15888_/X HRESETn VGND VGND VPWR VPWR _24796_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23015__A _22946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11760_/X VGND VGND VPWR VPWR _11761_/X sky130_fd_sc_hd__buf_2
X_23747_ _23747_/CLK _19409_/X VGND VGND VPWR VPWR _23747_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ _20828_/X _20958_/X _16639_/A _20874_/X VGND VGND VPWR VPWR _20959_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13498_/Y _13494_/X _11786_/X _13499_/X VGND VGND VPWR VPWR _25309_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14477_/Y _14475_/X _14479_/X _14475_/X VGND VGND VPWR VPWR _14480_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11683_/X VGND VGND VPWR VPWR _11692_/X sky130_fd_sc_hd__buf_2
X_23678_ _23678_/CLK _23678_/D VGND VGND VPWR VPWR _19612_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22854__A _23328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _13431_/A _13431_/B VGND VGND VPWR VPWR _13431_/X sky130_fd_sc_hd__or2_4
X_25417_ _25409_/CLK _12674_/X HRESETn VGND VGND VPWR VPWR _12508_/A sky130_fd_sc_hd__dfrtp_4
X_22629_ _22629_/A _22629_/B _22628_/X VGND VGND VPWR VPWR _22650_/C sky130_fd_sc_hd__and3_4
XFILLER_186_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16150_ _16124_/A VGND VGND VPWR VPWR _16150_/X sky130_fd_sc_hd__buf_2
X_13362_ _13394_/A _13362_/B _13362_/C VGND VGND VPWR VPWR _13370_/B sky130_fd_sc_hd__or3_4
X_25348_ _25346_/CLK _25348_/D HRESETn VGND VGND VPWR VPWR _12340_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21844__A2 _21325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24631__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15101_ _24983_/Q _24587_/Q _15294_/C _15100_/Y VGND VGND VPWR VPWR _15101_/X sky130_fd_sc_hd__o22a_4
X_12313_ _25342_/Q _24827_/Q _13072_/A _12312_/Y VGND VGND VPWR VPWR _12314_/D sky130_fd_sc_hd__o22a_4
XFILLER_6_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16081_ _23316_/A VGND VGND VPWR VPWR _16081_/Y sky130_fd_sc_hd__inv_2
X_13293_ _13293_/A _13293_/B _13292_/X VGND VGND VPWR VPWR _13302_/B sky130_fd_sc_hd__or3_4
X_25279_ _23528_/CLK _13752_/X HRESETn VGND VGND VPWR VPWR _25279_/Q sky130_fd_sc_hd__dfrtp_4
X_15032_ _15245_/A _24453_/Q _15245_/A _24453_/Q VGND VGND VPWR VPWR _15035_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12244_ _12266_/C _24752_/Q _12264_/A _12243_/Y VGND VGND VPWR VPWR _12244_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12604__B _12569_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19840_ _19835_/A VGND VGND VPWR VPWR _19840_/X sky130_fd_sc_hd__buf_2
X_12175_ _12175_/A VGND VGND VPWR VPWR _12176_/A sky130_fd_sc_hd__inv_2
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16484__B1 _16483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18498__B _18774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19771_ _19771_/A VGND VGND VPWR VPWR _21888_/B sky130_fd_sc_hd__inv_2
X_16983_ _24718_/Q _24375_/Q _16069_/Y _16982_/Y VGND VGND VPWR VPWR _16983_/X sky130_fd_sc_hd__o22a_4
X_18722_ _18698_/A _18719_/X VGND VGND VPWR VPWR _18722_/X sky130_fd_sc_hd__or2_4
XFILLER_237_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25490__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15934_ _12243_/Y _15932_/X _15560_/X _15932_/X VGND VGND VPWR VPWR _24776_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19422__B1 _19351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21711__A1_N _12252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18653_ _16582_/Y _18769_/A _16582_/Y _18769_/A VGND VGND VPWR VPWR _18653_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15865_ _15861_/X VGND VGND VPWR VPWR _15865_/X sky130_fd_sc_hd__buf_2
X_17604_ _17625_/A VGND VGND VPWR VPWR _17604_/X sky130_fd_sc_hd__buf_2
XFILLER_236_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14816_ _25201_/Q _14805_/X _14806_/X _14815_/Y VGND VGND VPWR VPWR _25056_/D sky130_fd_sc_hd__o22a_4
X_18584_ _18579_/B _18583_/X _18593_/C VGND VGND VPWR VPWR _18584_/X sky130_fd_sc_hd__and3_4
X_15796_ _15792_/X VGND VGND VPWR VPWR _15796_/X sky130_fd_sc_hd__buf_2
X_17535_ _11737_/Y _17659_/A _11737_/Y _17659_/A VGND VGND VPWR VPWR _17535_/X sky130_fd_sc_hd__a2bb2o_4
X_11959_ _18900_/A _11956_/X _11948_/B _11853_/X VGND VGND VPWR VPWR _11962_/A sky130_fd_sc_hd__o22a_4
X_14747_ _14678_/X _14739_/X VGND VGND VPWR VPWR _14747_/X sky130_fd_sc_hd__and2_4
XANTENNA__13470__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18019__A _18060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_10_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_10_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_14678_ _21902_/A VGND VGND VPWR VPWR _14678_/X sky130_fd_sc_hd__buf_2
X_17466_ _24208_/Q _19208_/B VGND VGND VPWR VPWR _17481_/B sky130_fd_sc_hd__and2_4
XFILLER_220_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24719__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19205_ _23819_/Q VGND VGND VPWR VPWR _19205_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13629_ _13627_/X _13629_/B VGND VGND VPWR VPWR _25301_/D sky130_fd_sc_hd__or2_4
X_16417_ _24591_/Q VGND VGND VPWR VPWR _16417_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23285__A1 _22552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17397_ _17399_/B VGND VGND VPWR VPWR _17398_/A sky130_fd_sc_hd__inv_2
XANTENNA__23285__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19136_ _19135_/Y _19133_/X _19067_/X _19133_/X VGND VGND VPWR VPWR _19136_/X sky130_fd_sc_hd__a2bb2o_4
X_16348_ _24616_/Q VGND VGND VPWR VPWR _16348_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24372__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16279_ _16278_/X VGND VGND VPWR VPWR _16279_/X sky130_fd_sc_hd__buf_2
X_19067_ _19360_/A VGND VGND VPWR VPWR _19067_/X sky130_fd_sc_hd__buf_2
XANTENNA__24301__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18018_ _18097_/A _18018_/B VGND VGND VPWR VPWR _18019_/C sky130_fd_sc_hd__or2_4
XFILLER_133_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21599__B2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17593__A _17625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_134_0_HCLK clkbuf_7_67_0_HCLK/X VGND VGND VPWR VPWR _23456_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_102_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_197_0_HCLK clkbuf_7_98_0_HCLK/X VGND VGND VPWR VPWR _24900_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_99_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15817__A3 _15746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25507__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19969_ _19969_/A VGND VGND VPWR VPWR _19969_/Y sky130_fd_sc_hd__inv_2
X_22980_ _22980_/A _22909_/B VGND VGND VPWR VPWR _22980_/X sky130_fd_sc_hd__or2_4
XANTENNA__16227__B1 _16226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21931_ _22015_/A VGND VGND VPWR VPWR _21936_/A sky130_fd_sc_hd__buf_2
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21843__A _16527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16043__A1_N _16042_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22658__B _22658_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24650_ _24650_/CLK _24650_/D HRESETn VGND VGND VPWR VPWR _24650_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_243_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15841__A _15670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14789__B1 _25057_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21862_ _24584_/Q _23088_/B VGND VGND VPWR VPWR _21866_/B sky130_fd_sc_hd__or2_4
X_23601_ _24199_/CLK _23601_/D VGND VGND VPWR VPWR _19837_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20813_ _13125_/A VGND VGND VPWR VPWR _20813_/Y sky130_fd_sc_hd__inv_2
X_24581_ _24591_/CLK _24581_/D HRESETn VGND VGND VPWR VPWR _15120_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21793_ _21656_/A _21791_/X _21792_/X VGND VGND VPWR VPWR _21793_/X sky130_fd_sc_hd__and3_4
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22720__B1 _11732_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23532_ _23411_/CLK _20028_/X VGND VGND VPWR VPWR _23532_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20744_ _13121_/A VGND VGND VPWR VPWR _20744_/Y sky130_fd_sc_hd__inv_2
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23463_ _23464_/CLK _23463_/D VGND VGND VPWR VPWR _18070_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_168_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17768__A _16913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23276__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20675_ _20495_/C _20675_/B _20674_/X VGND VGND VPWR VPWR _20675_/X sky130_fd_sc_hd__and3_4
XFILLER_149_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16688__A1_N _16687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23276__B2 _22838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25202_ _25043_/CLK _14206_/X HRESETn VGND VGND VPWR VPWR _20678_/A sky130_fd_sc_hd__dfrtp_4
X_22414_ _21077_/X _22411_/X _22946_/A _22413_/X VGND VGND VPWR VPWR _22414_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23394_ _25272_/CLK _23394_/D VGND VGND VPWR VPWR _21216_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_136_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25133_ _25134_/CLK _14436_/X HRESETn VGND VGND VPWR VPWR _25133_/Q sky130_fd_sc_hd__dfstp_4
X_22345_ _21933_/A _22345_/B _22344_/X VGND VGND VPWR VPWR _22345_/X sky130_fd_sc_hd__and3_4
XANTENNA__24042__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13516__A1 _13503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_30_0_HCLK clkbuf_7_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_30_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_25064_ _23526_/CLK _25064_/D HRESETn VGND VGND VPWR VPWR _25064_/Q sky130_fd_sc_hd__dfrtp_4
X_22276_ _22276_/A _22275_/X VGND VGND VPWR VPWR _22276_/X sky130_fd_sc_hd__or2_4
XFILLER_128_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_93_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_24015_ _24049_/CLK _24015_/D HRESETn VGND VGND VPWR VPWR _13120_/A sky130_fd_sc_hd__dfrtp_4
X_21227_ _22794_/A VGND VGND VPWR VPWR _21227_/X sky130_fd_sc_hd__buf_2
XFILLER_151_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25248__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21158_ _25244_/Q VGND VGND VPWR VPWR _21158_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23993__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20109_ _16880_/A VGND VGND VPWR VPWR _20109_/X sky130_fd_sc_hd__buf_2
X_13980_ _13980_/A _25240_/Q _13979_/X VGND VGND VPWR VPWR _13980_/X sky130_fd_sc_hd__or3_4
XANTENNA__19404__B1 _19357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21089_ _21015_/B _21089_/B VGND VGND VPWR VPWR _21089_/X sky130_fd_sc_hd__and2_4
XFILLER_219_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16218__B1 _15951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22849__A _22130_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12931_ _12762_/Y _12948_/A _12781_/Y _12947_/B VGND VGND VPWR VPWR _12931_/X sky130_fd_sc_hd__or4_4
X_24917_ _24508_/CLK _24917_/D HRESETn VGND VGND VPWR VPWR _15572_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12862_ _12887_/A VGND VGND VPWR VPWR _12862_/X sky130_fd_sc_hd__buf_2
X_15650_ _15649_/Y VGND VGND VPWR VPWR _15651_/A sky130_fd_sc_hd__buf_2
XFILLER_74_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24848_ _25341_/CLK _24848_/D HRESETn VGND VGND VPWR VPWR _24848_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _11805_/X _11813_/B _11809_/X _11813_/D VGND VGND VPWR VPWR _11813_/X sky130_fd_sc_hd__or4_4
X_14601_ _25083_/Q _14588_/X _13758_/X _14549_/B VGND VGND VPWR VPWR _14601_/X sky130_fd_sc_hd__o22a_4
XPHY_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ HWDATA[21] VGND VGND VPWR VPWR _15581_/X sky130_fd_sc_hd__buf_2
XFILLER_27_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12793_ _12793_/A VGND VGND VPWR VPWR _12793_/Y sky130_fd_sc_hd__inv_2
X_24779_ _25380_/CLK _24779_/D HRESETn VGND VGND VPWR VPWR _23307_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_221_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24883__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _13995_/X _14032_/Y _14532_/C VGND VGND VPWR VPWR _14532_/X sky130_fd_sc_hd__or3_4
X_17320_ _17338_/A _17314_/X _17320_/C VGND VGND VPWR VPWR _17320_/X sky130_fd_sc_hd__and3_4
XPHY_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11766_/A VGND VGND VPWR VPWR _11744_/X sky130_fd_sc_hd__buf_2
XFILLER_202_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24812__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14468_/A VGND VGND VPWR VPWR _14463_/X sky130_fd_sc_hd__buf_2
X_17251_ _17179_/Y _17200_/Y _17251_/C _17314_/C VGND VGND VPWR VPWR _17252_/D sky130_fd_sc_hd__or4_4
XFILLER_159_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _16446_/D VGND VGND VPWR VPWR _11676_/B sky130_fd_sc_hd__buf_2
XFILLER_230_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23267__B2 _22846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _13227_/X _13414_/B VGND VGND VPWR VPWR _13414_/X sky130_fd_sc_hd__or2_4
X_16202_ _23074_/A VGND VGND VPWR VPWR _16202_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17182_ _24620_/Q _24349_/Q _16339_/Y _17243_/B VGND VGND VPWR VPWR _17188_/B sky130_fd_sc_hd__o22a_4
X_14394_ _25145_/Q VGND VGND VPWR VPWR _14394_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16133_ _22638_/A VGND VGND VPWR VPWR _16133_/Y sky130_fd_sc_hd__inv_2
X_13345_ _13345_/A _13341_/X _13344_/X VGND VGND VPWR VPWR _13345_/X sky130_fd_sc_hd__or3_4
XFILLER_182_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16064_ _24720_/Q VGND VGND VPWR VPWR _16064_/Y sky130_fd_sc_hd__inv_2
X_13276_ _13231_/X _13273_/X _13275_/X VGND VGND VPWR VPWR _13276_/X sky130_fd_sc_hd__and3_4
XFILLER_155_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15015_ _25021_/Q _24459_/Q _15204_/A _15014_/Y VGND VGND VPWR VPWR _15015_/X sky130_fd_sc_hd__o22a_4
X_12227_ _12226_/X _24762_/Q _12273_/B _24762_/Q VGND VGND VPWR VPWR _12227_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15926__A _15925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16457__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17216__A2_N _21856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_207_0_HCLK clkbuf_8_206_0_HCLK/A VGND VGND VPWR VPWR _24555_/CLK sky130_fd_sc_hd__clkbuf_1
X_19823_ _19805_/Y VGND VGND VPWR VPWR _19823_/X sky130_fd_sc_hd__buf_2
XANTENNA__21450__B1 _21449_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12158_ _20971_/B _12157_/X SCLK_S3 _20971_/B VGND VGND VPWR VPWR _12158_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19754_ _19740_/A VGND VGND VPWR VPWR _19754_/X sky130_fd_sc_hd__buf_2
X_12089_ _12089_/A VGND VGND VPWR VPWR _12102_/A sky130_fd_sc_hd__inv_2
X_16966_ _24737_/Q _17032_/A _24743_/Q _16965_/Y VGND VGND VPWR VPWR _16966_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18705_ _18774_/A _18705_/B VGND VGND VPWR VPWR _18705_/X sky130_fd_sc_hd__and2_4
X_15917_ _15642_/X _15829_/X _15838_/X _21015_/B _15916_/X VGND VGND VPWR VPWR _24782_/D
+ sky130_fd_sc_hd__a32o_4
X_19685_ _19672_/Y VGND VGND VPWR VPWR _19685_/X sky130_fd_sc_hd__buf_2
X_16897_ _24279_/Q VGND VGND VPWR VPWR _17817_/A sky130_fd_sc_hd__inv_2
XFILLER_49_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15661__A _15661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18636_ _16615_/A _24128_/Q _16615_/Y _18819_/A VGND VGND VPWR VPWR _18637_/D sky130_fd_sc_hd__o22a_4
XFILLER_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15848_ _22816_/A VGND VGND VPWR VPWR _15958_/A sky130_fd_sc_hd__buf_2
XFILLER_91_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18567_ _18567_/A _18567_/B VGND VGND VPWR VPWR _18567_/X sky130_fd_sc_hd__or2_4
X_15779_ _15778_/X VGND VGND VPWR VPWR _15780_/B sky130_fd_sc_hd__buf_2
XFILLER_33_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17518_ _17516_/A _24112_/Q _17516_/Y _17517_/Y VGND VGND VPWR VPWR _17518_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24553__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18498_ _16441_/X _18774_/A VGND VGND VPWR VPWR _18498_/X sky130_fd_sc_hd__and2_4
XANTENNA__22494__A _22494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17449_ _18910_/B VGND VGND VPWR VPWR _18326_/B sky130_fd_sc_hd__inv_2
XFILLER_177_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23258__B2 _22290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16492__A _16492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20460_ _23999_/Q _20448_/X _20453_/X _20459_/Y VGND VGND VPWR VPWR _20460_/X sky130_fd_sc_hd__a211o_4
XFILLER_146_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19119_ _19133_/A VGND VGND VPWR VPWR _19119_/X sky130_fd_sc_hd__buf_2
XFILLER_118_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20391_ _13206_/B VGND VGND VPWR VPWR _20391_/Y sky130_fd_sc_hd__inv_2
X_22130_ _22130_/A _22130_/B VGND VGND VPWR VPWR _22130_/X sky130_fd_sc_hd__or2_4
XANTENNA__20492__A1 _20517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_17_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_161_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22061_ _22385_/A _19768_/Y VGND VGND VPWR VPWR _22061_/X sky130_fd_sc_hd__or2_4
XFILLER_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21557__B _21721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18212__A _18052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14740__A _14739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14429__A1_N _14428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21012_ _21012_/A _21012_/B VGND VGND VPWR VPWR _21012_/X sky130_fd_sc_hd__and2_4
XFILLER_245_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25341__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13356__A _13388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22963_ _22962_/X VGND VGND VPWR VPWR _22963_/Y sky130_fd_sc_hd__inv_2
XFILLER_244_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21914_ _21896_/X _21914_/B _21913_/X VGND VGND VPWR VPWR _21914_/X sky130_fd_sc_hd__and3_4
X_24702_ _24696_/CLK _16112_/X HRESETn VGND VGND VPWR VPWR _22980_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22894_ _23005_/A _22890_/X _22894_/C VGND VGND VPWR VPWR _22895_/D sky130_fd_sc_hd__and3_4
XANTENNA__16620__B1 _16361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24633_ _24629_/CLK _16307_/X HRESETn VGND VGND VPWR VPWR _24633_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21845_ _21845_/A _21842_/X _21845_/C VGND VGND VPWR VPWR _21845_/X sky130_fd_sc_hd__and3_4
XANTENNA__13803__B _17410_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14187__A _20628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_230_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24564_ _24540_/CLK _24564_/D HRESETn VGND VGND VPWR VPWR _16492_/A sky130_fd_sc_hd__dfrtp_4
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24294__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21776_ _21771_/A _20043_/Y VGND VGND VPWR VPWR _21777_/C sky130_fd_sc_hd__or2_4
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17176__B2 _17175_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23515_ _23388_/CLK _20064_/X VGND VGND VPWR VPWR _13431_/B sky130_fd_sc_hd__dfxtp_4
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20727_ _20727_/A VGND VGND VPWR VPWR _20727_/Y sky130_fd_sc_hd__inv_2
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24223__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24495_ _24427_/CLK _16678_/X HRESETn VGND VGND VPWR VPWR _24495_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_211_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23446_ _23808_/CLK _23446_/D VGND VGND VPWR VPWR _20252_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_11_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20812__A1_N _20690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20658_ _14222_/Y _20638_/X _20629_/A _20657_/X VGND VGND VPWR VPWR _20659_/A sky130_fd_sc_hd__a211o_4
XFILLER_149_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23377_ _23859_/CLK _20427_/X VGND VGND VPWR VPWR _23377_/Q sky130_fd_sc_hd__dfxtp_4
X_20589_ _18882_/B _20589_/B _20572_/X VGND VGND VPWR VPWR _20589_/X sky130_fd_sc_hd__and3_4
XFILLER_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13130_ _25334_/Q _13128_/X _13129_/Y VGND VGND VPWR VPWR _13130_/X sky130_fd_sc_hd__o21a_4
X_25116_ _25146_/CLK _14476_/X HRESETn VGND VGND VPWR VPWR _25116_/Q sky130_fd_sc_hd__dfrtp_4
X_22328_ _14174_/Y _14182_/A _14242_/Y _14245_/A VGND VGND VPWR VPWR _22328_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21748__A _21748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13061_ _13063_/B VGND VGND VPWR VPWR _13062_/B sky130_fd_sc_hd__inv_2
X_25047_ _25050_/CLK _25047_/D HRESETn VGND VGND VPWR VPWR _25047_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15746__A HWDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22259_ _22255_/A _22259_/B VGND VGND VPWR VPWR _22260_/C sky130_fd_sc_hd__or2_4
XFILLER_79_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18122__A _18014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12012_ _12012_/A _12004_/X _12012_/C _12012_/D VGND VGND VPWR VPWR _12013_/B sky130_fd_sc_hd__or4_4
XFILLER_151_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16439__B1 _16361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25082__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16820_ _16820_/A VGND VGND VPWR VPWR _16820_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25011__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_180_0_HCLK clkbuf_7_90_0_HCLK/X VGND VGND VPWR VPWR _25117_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_120_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_37_0_HCLK clkbuf_8_37_0_HCLK/A VGND VGND VPWR VPWR _25070_/CLK sky130_fd_sc_hd__clkbuf_1
X_16751_ _24464_/Q VGND VGND VPWR VPWR _16751_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13963_ _25242_/Q VGND VGND VPWR VPWR _14028_/A sky130_fd_sc_hd__inv_2
XFILLER_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17939__B1 _18020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21735__A1 _21556_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15702_ HWDATA[31] VGND VGND VPWR VPWR _15702_/X sky130_fd_sc_hd__buf_2
XFILLER_219_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12914_ _12800_/A _12914_/B VGND VGND VPWR VPWR _12914_/X sky130_fd_sc_hd__or2_4
X_19470_ _19457_/Y VGND VGND VPWR VPWR _19470_/X sky130_fd_sc_hd__buf_2
X_13894_ _13934_/B _13894_/B _13935_/A _13943_/D VGND VGND VPWR VPWR _13958_/B sky130_fd_sc_hd__and4_4
X_16682_ _16682_/A VGND VGND VPWR VPWR _16682_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18421_ _24649_/Q _18420_/A _16261_/Y _18420_/Y VGND VGND VPWR VPWR _18424_/C sky130_fd_sc_hd__o22a_4
X_12845_ _12769_/Y _12857_/A _12845_/C _12857_/B VGND VGND VPWR VPWR _12848_/B sky130_fd_sc_hd__or4_4
X_15633_ _15632_/Y _15628_/X _14479_/X _15628_/X VGND VGND VPWR VPWR _15633_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18352_ _21979_/A VGND VGND VPWR VPWR _18352_/Y sky130_fd_sc_hd__inv_2
X_12776_ _24787_/Q VGND VGND VPWR VPWR _12776_/Y sky130_fd_sc_hd__inv_2
X_15564_ HWDATA[27] VGND VGND VPWR VPWR _15564_/X sky130_fd_sc_hd__buf_2
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17341_/A VGND VGND VPWR VPWR _17338_/A sky130_fd_sc_hd__buf_2
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11725_/Y _11723_/X _11726_/X _11723_/X VGND VGND VPWR VPWR _25536_/D sky130_fd_sc_hd__a2bb2o_4
X_14515_ _25105_/Q _14499_/X _25104_/Q _14494_/X VGND VGND VPWR VPWR _14515_/X sky130_fd_sc_hd__o22a_4
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15493_/Y _15494_/X HADDR[19] _15494_/X VGND VGND VPWR VPWR _24944_/D sky130_fd_sc_hd__a2bb2o_4
X_18283_ _17704_/X VGND VGND VPWR VPWR _18283_/X sky130_fd_sc_hd__buf_2
XFILLER_159_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16914__B2 _16913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17234_ _17298_/A VGND VGND VPWR VPWR _17234_/Y sky130_fd_sc_hd__inv_2
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _24067_/Q VGND VGND VPWR VPWR _11659_/A sky130_fd_sc_hd__inv_2
X_14446_ _14445_/Y _14443_/X _14403_/X _14443_/X VGND VGND VPWR VPWR _25128_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_156_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14544__B _13577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _20430_/A VGND VGND VPWR VPWR _20462_/A sky130_fd_sc_hd__inv_2
X_17165_ _24347_/Q VGND VGND VPWR VPWR _17165_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23946__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16678__B1 _16320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13328_ _13200_/A _20231_/A VGND VGND VPWR VPWR _13328_/X sky130_fd_sc_hd__or2_4
X_16116_ _16111_/A VGND VGND VPWR VPWR _16116_/X sky130_fd_sc_hd__buf_2
XFILLER_115_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17096_ _17095_/X VGND VGND VPWR VPWR _24393_/D sky130_fd_sc_hd__inv_2
X_13259_ _13334_/A _18917_/A VGND VGND VPWR VPWR _13259_/X sky130_fd_sc_hd__or2_4
X_16047_ _24726_/Q VGND VGND VPWR VPWR _16047_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12164__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19092__B2 _19074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19806_ _19805_/Y VGND VGND VPWR VPWR _19806_/X sky130_fd_sc_hd__buf_2
XFILLER_229_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17998_ _18095_/A VGND VGND VPWR VPWR _18085_/A sky130_fd_sc_hd__buf_2
XANTENNA__16850__B1 _16849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21393__A _22197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19737_ _23634_/Q VGND VGND VPWR VPWR _19737_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16949_ _16929_/X _16934_/X _16949_/C _16948_/X VGND VGND VPWR VPWR _16950_/B sky130_fd_sc_hd__or4_4
XFILLER_37_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21726__B2 _21351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19668_ _13435_/B VGND VGND VPWR VPWR _19668_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24734__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_8_0_HCLK clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__16602__B1 _16601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18619_ _24144_/Q VGND VGND VPWR VPWR _18760_/A sky130_fd_sc_hd__inv_2
X_19599_ _19598_/Y VGND VGND VPWR VPWR _19599_/X sky130_fd_sc_hd__buf_2
XFILLER_212_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21630_ _21771_/A _21630_/B VGND VGND VPWR VPWR _21631_/C sky130_fd_sc_hd__or2_4
XFILLER_52_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22151__B2 _23171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21561_ _21561_/A VGND VGND VPWR VPWR _21564_/C sky130_fd_sc_hd__inv_2
XFILLER_221_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23300_ _22708_/A _23297_/X _23299_/X VGND VGND VPWR VPWR _23305_/C sky130_fd_sc_hd__and3_4
X_20512_ _20488_/B VGND VGND VPWR VPWR _20512_/Y sky130_fd_sc_hd__inv_2
X_24280_ _24275_/CLK _17809_/Y HRESETn VGND VGND VPWR VPWR _24280_/Q sky130_fd_sc_hd__dfrtp_4
X_21492_ _21487_/A _21492_/B VGND VGND VPWR VPWR _21493_/C sky130_fd_sc_hd__or2_4
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23231_ _23229_/X _23231_/B _22140_/A VGND VGND VPWR VPWR _23231_/X sky130_fd_sc_hd__or3_4
X_20443_ _20441_/Y VGND VGND VPWR VPWR _20444_/B sky130_fd_sc_hd__buf_2
XFILLER_181_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22671__B _21047_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16669__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23162_ _17255_/A _22916_/X _25394_/Q _22917_/X VGND VGND VPWR VPWR _23162_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25522__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20374_ _20374_/A VGND VGND VPWR VPWR _20374_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22113_ _22110_/X _22112_/X _21111_/A VGND VGND VPWR VPWR _22113_/Y sky130_fd_sc_hd__a21oi_4
X_23093_ _12195_/Y _22718_/X _22719_/X _12309_/Y _22846_/X VGND VGND VPWR VPWR _23093_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__25142__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21414__B1 _14672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22044_ _22044_/A _19594_/Y _22043_/X VGND VGND VPWR VPWR _22044_/X sky130_fd_sc_hd__and3_4
XFILLER_161_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17781__A _16913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_253_0_HCLK clkbuf_7_126_0_HCLK/X VGND VGND VPWR VPWR _24959_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_236_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23995_ _24146_/CLK _23995_/D HRESETn VGND VGND VPWR VPWR _23995_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16397__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21717__B2 _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22946_ _22946_/A _22943_/X _22945_/X VGND VGND VPWR VPWR _22965_/B sky130_fd_sc_hd__and3_4
XFILLER_216_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24475__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22390__A1 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22877_ _16672_/Y _22921_/B VGND VGND VPWR VPWR _22877_/X sky130_fd_sc_hd__and2_4
XANTENNA__24404__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12630_ _12681_/A _12630_/B VGND VGND VPWR VPWR _12633_/B sky130_fd_sc_hd__or2_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21828_ _21821_/Y _21827_/X _22041_/A VGND VGND VPWR VPWR _21828_/X sky130_fd_sc_hd__o21a_4
X_24616_ _24662_/CLK _16351_/X HRESETn VGND VGND VPWR VPWR _24616_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12561_ _12608_/A _24878_/Q _12608_/A _24878_/Q VGND VGND VPWR VPWR _12561_/X sky130_fd_sc_hd__a2bb2o_4
X_24547_ _24133_/CLK _16537_/X HRESETn VGND VGND VPWR VPWR _24547_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16947__A2_N _22190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21759_ _21609_/X _21759_/B VGND VGND VPWR VPWR _21759_/X sky130_fd_sc_hd__or2_4
XFILLER_196_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14300_ _14294_/A VGND VGND VPWR VPWR _14300_/X sky130_fd_sc_hd__buf_2
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17021__A _17020_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15280_ _15311_/B VGND VGND VPWR VPWR _15281_/A sky130_fd_sc_hd__buf_2
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12492_ _12492_/A _12456_/X VGND VGND VPWR VPWR _12493_/C sky130_fd_sc_hd__nand2_4
X_24478_ _24976_/CLK _16722_/X HRESETn VGND VGND VPWR VPWR _15285_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ _14231_/A VGND VGND VPWR VPWR _14231_/Y sky130_fd_sc_hd__inv_2
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23429_ _23534_/CLK _23429_/D VGND VGND VPWR VPWR _20297_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14162_ _14162_/A _14161_/X VGND VGND VPWR VPWR _14162_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21653__B1 _13772_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21478__A _17709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13113_ _13113_/A _13113_/B VGND VGND VPWR VPWR _13113_/X sky130_fd_sc_hd__or2_4
XFILLER_124_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14093_ _14092_/X VGND VGND VPWR VPWR _14093_/Y sky130_fd_sc_hd__inv_2
X_18970_ _18970_/A VGND VGND VPWR VPWR _18970_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14380__A _14380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_63_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13044_ _12302_/Y _13048_/B _13043_/Y VGND VGND VPWR VPWR _25354_/D sky130_fd_sc_hd__o21a_4
X_17921_ _24251_/Q VGND VGND VPWR VPWR _17921_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17852_ _17748_/Y _17852_/B VGND VGND VPWR VPWR _17853_/D sky130_fd_sc_hd__or2_4
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23158__B1 _25546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16803_ _24440_/Q VGND VGND VPWR VPWR _16803_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16832__B1 _15746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15635__B2 _15553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17783_ _17791_/A VGND VGND VPWR VPWR _17783_/X sky130_fd_sc_hd__buf_2
X_14995_ _14995_/A VGND VGND VPWR VPWR _14995_/X sky130_fd_sc_hd__buf_2
X_19522_ _19522_/A _14181_/A VGND VGND VPWR VPWR _21215_/A sky130_fd_sc_hd__or2_4
XFILLER_235_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16734_ _15010_/Y _16730_/X _16467_/X _16730_/X VGND VGND VPWR VPWR _24473_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13946_ _24975_/Q _13927_/B VGND VGND VPWR VPWR _13947_/B sky130_fd_sc_hd__or2_4
XFILLER_234_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19453_ _23730_/Q VGND VGND VPWR VPWR _22350_/B sky130_fd_sc_hd__inv_2
XFILLER_35_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16665_ _24500_/Q VGND VGND VPWR VPWR _16665_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20392__B1 _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24145__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13877_ _24975_/Q VGND VGND VPWR VPWR _13924_/A sky130_fd_sc_hd__buf_2
XFILLER_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15938__A2 _15928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18404_ _22996_/A _18468_/A _23206_/A _18505_/A VGND VGND VPWR VPWR _18404_/X sky130_fd_sc_hd__a2bb2o_4
X_15616_ _14400_/A VGND VGND VPWR VPWR _15616_/X sky130_fd_sc_hd__buf_2
XFILLER_62_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12828_ _12828_/A VGND VGND VPWR VPWR _12857_/A sky130_fd_sc_hd__inv_2
X_19384_ _18200_/B VGND VGND VPWR VPWR _19384_/Y sky130_fd_sc_hd__inv_2
X_16596_ _24524_/Q VGND VGND VPWR VPWR _16596_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23330__B1 _21339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18335_ _20220_/A VGND VGND VPWR VPWR _19716_/C sky130_fd_sc_hd__buf_2
X_15547_ _16637_/A _15773_/A VGND VGND VPWR VPWR _15550_/A sky130_fd_sc_hd__or2_4
X_12759_ _25392_/Q VGND VGND VPWR VPWR _12759_/Y sky130_fd_sc_hd__inv_2
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18266_ _23346_/A _18265_/Y _16778_/X _18265_/Y VGND VGND VPWR VPWR _24225_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_202_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15478_ _24068_/Q VGND VGND VPWR VPWR _15478_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17217_ _24361_/Q VGND VGND VPWR VPWR _17249_/D sky130_fd_sc_hd__inv_2
X_14429_ _14428_/Y _14426_/X _14403_/X _14426_/X VGND VGND VPWR VPWR _25136_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15571__B1 _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18197_ _15691_/A _18181_/X _18196_/X _24244_/Q _18022_/A VGND VGND VPWR VPWR _18197_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_156_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22436__A2 _21833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12075__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17148_ _17127_/X _17148_/B _17148_/C VGND VGND VPWR VPWR _24378_/D sky130_fd_sc_hd__and3_4
XFILLER_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17079_ _16973_/Y _17075_/X VGND VGND VPWR VPWR _17080_/C sky130_fd_sc_hd__nand2_4
XFILLER_143_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20090_ _22375_/B _20088_/X _20089_/X _20088_/X VGND VGND VPWR VPWR _23506_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24986__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24915__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16823__B1 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23108__A _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22800_ _16404_/A _22800_/B VGND VGND VPWR VPWR _22800_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_20_0_HCLK clkbuf_8_21_0_HCLK/A VGND VGND VPWR VPWR _23427_/CLK sky130_fd_sc_hd__clkbuf_1
X_23780_ _24252_/CLK _23780_/D VGND VGND VPWR VPWR _18170_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_226_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20992_ _20992_/A _20990_/Y VGND VGND VPWR VPWR _20992_/Y sky130_fd_sc_hd__nor2_4
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_83_0_HCLK clkbuf_8_83_0_HCLK/A VGND VGND VPWR VPWR _25380_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_225_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22731_ _24461_/Q _22534_/X _22535_/X VGND VGND VPWR VPWR _22731_/X sky130_fd_sc_hd__o21a_4
XFILLER_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15929__A2 _15928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15036__A1_N _25014_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22666__B _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25450_ _25450_/CLK _12437_/X HRESETn VGND VGND VPWR VPWR _12234_/A sky130_fd_sc_hd__dfrtp_4
X_22662_ _22662_/A _22661_/X VGND VGND VPWR VPWR _22662_/X sky130_fd_sc_hd__or2_4
XFILLER_197_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24401_ _23427_/CLK _24401_/D HRESETn VGND VGND VPWR VPWR _24401_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_201_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23321__B1 _25399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21613_ _21608_/X _21612_/X _14707_/X VGND VGND VPWR VPWR _21613_/X sky130_fd_sc_hd__o21a_4
X_25381_ _25390_/CLK _12924_/X HRESETn VGND VGND VPWR VPWR _12793_/A sky130_fd_sc_hd__dfrtp_4
X_22593_ _22629_/A _22590_/X _22592_/X VGND VGND VPWR VPWR _22614_/C sky130_fd_sc_hd__and3_4
Xclkbuf_2_3_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24332_ _24980_/CLK _24332_/D HRESETn VGND VGND VPWR VPWR _24332_/Q sky130_fd_sc_hd__dfrtp_4
X_21544_ _21532_/X _21536_/Y _22712_/A _21543_/X VGND VGND VPWR VPWR _21544_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24263_ _24263_/CLK _24263_/D HRESETn VGND VGND VPWR VPWR _16925_/A sky130_fd_sc_hd__dfrtp_4
X_21475_ _21475_/A _21475_/B _21474_/X VGND VGND VPWR VPWR _21475_/X sky130_fd_sc_hd__and3_4
XFILLER_194_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15562__B1 _15560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23214_ _23182_/A _23205_/Y _23214_/C _23214_/D VGND VGND VPWR VPWR _23214_/X sky130_fd_sc_hd__or4_4
XFILLER_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20426_ _23377_/Q VGND VGND VPWR VPWR _21253_/B sky130_fd_sc_hd__inv_2
XFILLER_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24194_ _25471_/CLK _18384_/X HRESETn VGND VGND VPWR VPWR _24194_/Q sky130_fd_sc_hd__dfrtp_4
X_23145_ _22146_/X VGND VGND VPWR VPWR _23145_/X sky130_fd_sc_hd__buf_2
X_20357_ _20357_/A VGND VGND VPWR VPWR _21940_/B sky130_fd_sc_hd__inv_2
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23076_ _24539_/Q _22730_/X _15663_/X _23075_/X VGND VGND VPWR VPWR _23076_/X sky130_fd_sc_hd__a211o_4
X_20288_ _20287_/Y VGND VGND VPWR VPWR _20288_/X sky130_fd_sc_hd__buf_2
XANTENNA__14230__A1_N _14229_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22027_ _22016_/A _22027_/B VGND VGND VPWR VPWR _22027_/X sky130_fd_sc_hd__or2_4
XANTENNA__14860__A1_N _14817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24656__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16814__B1 _16483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13800_ _12084_/A _13800_/B VGND VGND VPWR VPWR _13800_/X sky130_fd_sc_hd__or2_4
XFILLER_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17016__A _17343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11992_ _11992_/A VGND VGND VPWR VPWR _11992_/Y sky130_fd_sc_hd__inv_2
X_14780_ _14628_/A VGND VGND VPWR VPWR _17983_/A sky130_fd_sc_hd__inv_2
X_23978_ _23976_/CLK _23978_/D HRESETn VGND VGND VPWR VPWR _20630_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_28_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13731_ _14755_/A _13726_/X _14775_/A _14764_/A VGND VGND VPWR VPWR _13731_/X sky130_fd_sc_hd__or4_4
XFILLER_232_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22929_ _24566_/Q _22885_/X _22802_/X VGND VGND VPWR VPWR _22929_/X sky130_fd_sc_hd__o21a_4
XFILLER_217_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20913__A2 _20846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16450_ _24578_/Q VGND VGND VPWR VPWR _16450_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13662_ _13630_/A _25297_/Q _25298_/Q VGND VGND VPWR VPWR _25297_/D sky130_fd_sc_hd__a21o_4
XFILLER_189_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15401_ _15294_/D _15385_/X VGND VGND VPWR VPWR _15401_/Y sky130_fd_sc_hd__nand2_4
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12613_ _12613_/A _12613_/B VGND VGND VPWR VPWR _12615_/B sky130_fd_sc_hd__or2_4
X_13593_ _13593_/A VGND VGND VPWR VPWR _13593_/Y sky130_fd_sc_hd__inv_2
X_16381_ _16387_/A VGND VGND VPWR VPWR _16381_/X sky130_fd_sc_hd__buf_2
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18120_ _18085_/A _18118_/X _18120_/C VGND VGND VPWR VPWR _18120_/X sky130_fd_sc_hd__and3_4
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12544_ _25419_/Q _24873_/Q _12664_/A _12543_/Y VGND VGND VPWR VPWR _12544_/X sky130_fd_sc_hd__o22a_4
X_15332_ _15130_/Y _15339_/A VGND VGND VPWR VPWR _15333_/B sky130_fd_sc_hd__or2_4
XFILLER_212_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12607__B _12606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18051_ _18124_/A _18047_/X _18050_/X VGND VGND VPWR VPWR _18062_/B sky130_fd_sc_hd__or3_4
X_12475_ _12217_/Y _12475_/B VGND VGND VPWR VPWR _12476_/B sky130_fd_sc_hd__or2_4
X_15263_ _15245_/A _15266_/B _15169_/X VGND VGND VPWR VPWR _15263_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_144_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17002_ _24401_/Q VGND VGND VPWR VPWR _17022_/A sky130_fd_sc_hd__inv_2
X_14214_ _14207_/Y _14213_/X _13824_/X _14213_/X VGND VGND VPWR VPWR _14214_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11709__A3 HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15194_ _14982_/A VGND VGND VPWR VPWR _15194_/X sky130_fd_sc_hd__buf_2
XFILLER_126_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14145_ _14103_/C _14088_/X _14103_/C _14088_/X VGND VGND VPWR VPWR _14145_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14076_ _14005_/A _14070_/X _14067_/X _14007_/D _14073_/X VGND VGND VPWR VPWR _14076_/X
+ sky130_fd_sc_hd__a32o_4
X_18953_ _18953_/A VGND VGND VPWR VPWR _18953_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21936__A _21936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13027_ _12986_/X _13005_/D _12349_/Y VGND VGND VPWR VPWR _13028_/C sky130_fd_sc_hd__o21a_4
X_17904_ _17906_/B _17901_/Y _17901_/A _17903_/X VGND VGND VPWR VPWR _17904_/X sky130_fd_sc_hd__o22a_4
X_18884_ _18884_/A VGND VGND VPWR VPWR _18885_/A sky130_fd_sc_hd__inv_2
XFILLER_67_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24397__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16805__B1 _15719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17835_ _17757_/A _17835_/B VGND VGND VPWR VPWR _17837_/B sky130_fd_sc_hd__or2_4
XANTENNA__24326__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17766_ _16898_/Y _17786_/B VGND VGND VPWR VPWR _17766_/X sky130_fd_sc_hd__or2_4
X_14978_ _14978_/A _14973_/X _14974_/X _14977_/X VGND VGND VPWR VPWR _14979_/D sky130_fd_sc_hd__or4_4
XANTENNA__21157__A2 _21348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22767__A _24764_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19505_ _23713_/Q VGND VGND VPWR VPWR _22236_/B sky130_fd_sc_hd__inv_2
X_16717_ _16715_/Y _16655_/A _16716_/X _16655_/A VGND VGND VPWR VPWR _24479_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_212_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13929_ _13928_/X VGND VGND VPWR VPWR _13929_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20365__B1 _19620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17697_ _17697_/A _17696_/Y _17688_/C VGND VGND VPWR VPWR _17697_/X sky130_fd_sc_hd__and3_4
XANTENNA__16765__A _16765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19436_ _19432_/Y _19435_/X _19414_/X _19435_/X VGND VGND VPWR VPWR _23738_/D sky130_fd_sc_hd__a2bb2o_4
X_16648_ _16655_/A VGND VGND VPWR VPWR _16648_/X sky130_fd_sc_hd__buf_2
XANTENNA__22106__B2 _21351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20287__A _20286_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20380__A3 _20061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19367_ _19372_/A VGND VGND VPWR VPWR _19367_/X sky130_fd_sc_hd__buf_2
X_16579_ _16547_/A VGND VGND VPWR VPWR _16598_/A sky130_fd_sc_hd__buf_2
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18980__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23961__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18318_ _18301_/A _18303_/B _18298_/B VGND VGND VPWR VPWR _18318_/X sky130_fd_sc_hd__o21a_4
XANTENNA__11702__A _11701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21865__B1 _21730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19298_ _19341_/A _19002_/B _19320_/C VGND VGND VPWR VPWR _19299_/A sky130_fd_sc_hd__or3_4
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18249_ _11833_/Y _18245_/X _16601_/X _18245_/X VGND VGND VPWR VPWR _24234_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21260_ _21884_/A _21260_/B VGND VGND VPWR VPWR _21261_/C sky130_fd_sc_hd__or2_4
XFILLER_117_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20211_ _20210_/Y _20206_/X _19728_/X _20206_/X VGND VGND VPWR VPWR _20211_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21191_ _21204_/A _21188_/X _21190_/X VGND VGND VPWR VPWR _21191_/X sky130_fd_sc_hd__and3_4
XFILLER_237_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20142_ _23488_/Q VGND VGND VPWR VPWR _20142_/Y sky130_fd_sc_hd__inv_2
X_20073_ _20071_/Y _20067_/X _19813_/X _20072_/X VGND VGND VPWR VPWR _20073_/X sky130_fd_sc_hd__a2bb2o_4
X_24950_ _24973_/CLK _24950_/D HRESETn VGND VGND VPWR VPWR _24950_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23901_ _23875_/CLK _18969_/X VGND VGND VPWR VPWR _23901_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24067__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24881_ _24834_/CLK _15720_/X HRESETn VGND VGND VPWR VPWR _24881_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23832_ _23846_/CLK _23832_/D VGND VGND VPWR VPWR _19169_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_122_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14179__B _14179_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23763_ _23767_/CLK _23763_/D VGND VGND VPWR VPWR _19362_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20975_ _12137_/X _12147_/A VGND VGND VPWR VPWR _24106_/D sky130_fd_sc_hd__and2_4
XFILLER_199_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20356__B1 _19606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25502_ _24209_/CLK _25502_/D HRESETn VGND VGND VPWR VPWR _18901_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_214_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22714_ _22714_/A _21124_/B _21864_/C VGND VGND VPWR VPWR _22714_/X sky130_fd_sc_hd__and3_4
XPHY_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23694_ _23437_/CLK _23694_/D VGND VGND VPWR VPWR _23694_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20371__A3 _11760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22645_ _22645_/A VGND VGND VPWR VPWR _22645_/Y sky130_fd_sc_hd__inv_2
X_25433_ _25444_/CLK _25433_/D HRESETn VGND VGND VPWR VPWR _21078_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25364_ _25346_/CLK _25364_/D HRESETn VGND VGND VPWR VPWR _12315_/A sky130_fd_sc_hd__dfrtp_4
X_22576_ _22575_/X VGND VGND VPWR VPWR _22577_/D sky130_fd_sc_hd__inv_2
XFILLER_166_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21320__A2 _21315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21527_ _21533_/A VGND VGND VPWR VPWR _21528_/B sky130_fd_sc_hd__buf_2
X_24315_ _24315_/CLK _17620_/X HRESETn VGND VGND VPWR VPWR _24315_/Q sky130_fd_sc_hd__dfrtp_4
X_25295_ _25091_/CLK _13688_/Y HRESETn VGND VGND VPWR VPWR _11820_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12260_ _12228_/X _12260_/B _12250_/X _12259_/X VGND VGND VPWR VPWR _12261_/B sky130_fd_sc_hd__or4_4
X_24246_ _23774_/CLK _18102_/X HRESETn VGND VGND VPWR VPWR _24246_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21458_ _22262_/A VGND VGND VPWR VPWR _21817_/A sky130_fd_sc_hd__buf_2
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20409_ _20408_/X VGND VGND VPWR VPWR _20409_/Y sky130_fd_sc_hd__inv_2
X_12191_ _12191_/A VGND VGND VPWR VPWR _12191_/X sky130_fd_sc_hd__buf_2
X_24177_ _24667_/CLK _24177_/D HRESETn VGND VGND VPWR VPWR _18407_/A sky130_fd_sc_hd__dfrtp_4
X_21389_ _21385_/X _21389_/B VGND VGND VPWR VPWR _21389_/X sky130_fd_sc_hd__or2_4
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24837__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23128_ _23128_/A VGND VGND VPWR VPWR _23182_/A sky130_fd_sc_hd__buf_2
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15754__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15950_ _12202_/Y _15944_/X _15948_/X _15949_/X VGND VGND VPWR VPWR _15950_/X sky130_fd_sc_hd__a2bb2o_4
X_23059_ _22786_/X _23057_/X _22789_/X _23058_/X VGND VGND VPWR VPWR _23060_/B sky130_fd_sc_hd__o22a_4
XFILLER_1_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24490__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14901_ _14898_/X _14899_/Y _14886_/A _14900_/Y VGND VGND VPWR VPWR _14901_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15881_ _15881_/A VGND VGND VPWR VPWR _15881_/X sky130_fd_sc_hd__buf_2
X_17620_ _17620_/A _17616_/X _17619_/Y VGND VGND VPWR VPWR _17620_/X sky130_fd_sc_hd__and3_4
XFILLER_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13274__A _13199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14832_ _14820_/X _14831_/Y _14812_/C _14820_/X VGND VGND VPWR VPWR _25053_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21139__A2 _14209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17551_ _17561_/A _17541_/Y _11772_/Y _24295_/Q VGND VGND VPWR VPWR _17551_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14763_ _14762_/X VGND VGND VPWR VPWR _14763_/Y sky130_fd_sc_hd__inv_2
X_11975_ _25495_/Q VGND VGND VPWR VPWR _11975_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16502_ _16500_/Y _16496_/X _16229_/X _16501_/X VGND VGND VPWR VPWR _16502_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_232_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13714_ _13670_/A _13669_/X VGND VGND VPWR VPWR _13714_/Y sky130_fd_sc_hd__nand2_4
XFILLER_204_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17482_ _17482_/A VGND VGND VPWR VPWR _17482_/Y sky130_fd_sc_hd__inv_2
X_14694_ _22213_/A VGND VGND VPWR VPWR _21901_/A sky130_fd_sc_hd__buf_2
XFILLER_204_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19221_ _18965_/A VGND VGND VPWR VPWR _19221_/X sky130_fd_sc_hd__buf_2
X_16433_ _16432_/Y _16430_/X _16353_/X _16430_/X VGND VGND VPWR VPWR _24583_/D sky130_fd_sc_hd__a2bb2o_4
X_13645_ _24041_/Q _13644_/X VGND VGND VPWR VPWR _20857_/B sky130_fd_sc_hd__or2_4
X_19152_ _19151_/Y _19149_/X _19057_/X _19149_/X VGND VGND VPWR VPWR _19152_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16364_ _16364_/A _14365_/B _14365_/C _14365_/D VGND VGND VPWR VPWR _16365_/A sky130_fd_sc_hd__or4_4
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13576_ _14764_/A VGND VGND VPWR VPWR _13577_/B sky130_fd_sc_hd__inv_2
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18103_ _18103_/A _18103_/B VGND VGND VPWR VPWR _18105_/B sky130_fd_sc_hd__or2_4
X_15315_ _15315_/A _15326_/A _15323_/A _15303_/X VGND VGND VPWR VPWR _15315_/X sky130_fd_sc_hd__or4_4
XFILLER_157_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12527_ _24879_/Q VGND VGND VPWR VPWR _12527_/Y sky130_fd_sc_hd__inv_2
X_19083_ _23862_/Q VGND VGND VPWR VPWR _21760_/B sky130_fd_sc_hd__inv_2
XFILLER_173_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16295_ HWDATA[25] VGND VGND VPWR VPWR _16295_/X sky130_fd_sc_hd__buf_2
XANTENNA__18305__A _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18034_ _17981_/A _18034_/B _18033_/X VGND VGND VPWR VPWR _18034_/X sky130_fd_sc_hd__and3_4
X_15246_ _15251_/A _15254_/A _15246_/C _15254_/B VGND VGND VPWR VPWR _15247_/A sky130_fd_sc_hd__or4_4
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12458_ _12266_/C _12458_/B VGND VGND VPWR VPWR _12475_/B sky130_fd_sc_hd__or2_4
X_12389_ _12413_/A _12387_/X _12388_/X VGND VGND VPWR VPWR _12389_/X sky130_fd_sc_hd__and3_4
X_15177_ _15168_/B _15168_/C _15169_/X _15173_/Y VGND VGND VPWR VPWR _15177_/X sky130_fd_sc_hd__a211o_4
XFILLER_141_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24578__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14128_ _14106_/A _14106_/B _14106_/A _14106_/B VGND VGND VPWR VPWR _14128_/X sky130_fd_sc_hd__a2bb2o_4
X_19985_ _19983_/Y _19980_/X _19984_/X _19980_/X VGND VGND VPWR VPWR _19985_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24507__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14059_ _14059_/A _14020_/Y VGND VGND VPWR VPWR _14060_/B sky130_fd_sc_hd__or2_4
X_18936_ _13208_/B VGND VGND VPWR VPWR _18936_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22575__B2 _22574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18867_ _18851_/X _18856_/X _18861_/X _18867_/D VGND VGND VPWR VPWR _18867_/X sky130_fd_sc_hd__or4_4
XANTENNA__24160__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13184__A _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17818_ _17818_/A _17818_/B _17818_/C VGND VGND VPWR VPWR _24279_/D sky130_fd_sc_hd__and3_4
X_18798_ _18798_/A VGND VGND VPWR VPWR _18798_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14265__B1 _13798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17749_ _21059_/A VGND VGND VPWR VPWR _17750_/D sky130_fd_sc_hd__inv_2
XFILLER_70_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16495__A _16453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20760_ _13107_/C _20754_/X VGND VGND VPWR VPWR _20760_/X sky130_fd_sc_hd__or2_4
XANTENNA__25366__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19419_ _19426_/A VGND VGND VPWR VPWR _19419_/X sky130_fd_sc_hd__buf_2
XFILLER_223_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20691_ _21124_/A _20687_/X _13110_/B _20690_/X VGND VGND VPWR VPWR _20692_/A sky130_fd_sc_hd__o22a_4
XANTENNA__15765__B1 _24858_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_157_0_HCLK clkbuf_7_78_0_HCLK/X VGND VGND VPWR VPWR _24325_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_195_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22944__B _22821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22430_ _22429_/X VGND VGND VPWR VPWR _22430_/X sky130_fd_sc_hd__buf_2
XFILLER_149_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23121__A _22730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22361_ _17709_/A _22357_/X _22358_/X _22359_/X _22360_/X VGND VGND VPWR VPWR _22361_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15517__B1 HADDR[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24100_ _25164_/CLK _14320_/Y HRESETn VGND VGND VPWR VPWR _14339_/A sky130_fd_sc_hd__dfrtp_4
X_21312_ _21311_/X VGND VGND VPWR VPWR _21312_/X sky130_fd_sc_hd__buf_2
XFILLER_248_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25080_ _25081_/CLK _25080_/D HRESETn VGND VGND VPWR VPWR _21964_/A sky130_fd_sc_hd__dfrtp_4
X_22292_ _22287_/X _22289_/X _22290_/X _22291_/X VGND VGND VPWR VPWR _22293_/B sky130_fd_sc_hd__o22a_4
X_24031_ _24508_/CLK _24031_/D HRESETn VGND VGND VPWR VPWR _13125_/B sky130_fd_sc_hd__dfrtp_4
X_21243_ _21262_/A _21243_/B VGND VGND VPWR VPWR _21243_/X sky130_fd_sc_hd__or2_4
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24930__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21174_ _16438_/Y _15662_/A _16365_/A _21173_/X VGND VGND VPWR VPWR _21175_/C sky130_fd_sc_hd__a211o_4
XFILLER_116_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17773__B _17602_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24248__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20125_ _20125_/A VGND VGND VPWR VPWR _21778_/B sky130_fd_sc_hd__inv_2
XFILLER_89_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_22_0_HCLK_A clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20056_ _20053_/X _18328_/X _11760_/X _13178_/B _20055_/X VGND VGND VPWR VPWR _20056_/X
+ sky130_fd_sc_hd__a32o_4
X_24933_ _25070_/CLK _24933_/D HRESETn VGND VGND VPWR VPWR _11674_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24864_ _25409_/CLK _24864_/D HRESETn VGND VGND VPWR VPWR _24864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22318__B2 _21351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23815_ _23873_/CLK _19219_/X VGND VGND VPWR VPWR _19218_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24795_ _24795_/CLK _15890_/X HRESETn VGND VGND VPWR VPWR _22553_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19195__B1 _19194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ HWDATA[7] VGND VGND VPWR VPWR _11760_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_53_0_HCLK clkbuf_7_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _20956_/Y _20957_/Y _13655_/B VGND VGND VPWR VPWR _20958_/X sky130_fd_sc_hd__o21a_4
X_23746_ _23785_/CLK _23746_/D VGND VGND VPWR VPWR _17956_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25036__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ HWDATA[23] VGND VGND VPWR VPWR _11691_/X sky130_fd_sc_hd__buf_2
XANTENNA__15756__B1 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _20889_/A _20888_/A VGND VGND VPWR VPWR _20889_/X sky130_fd_sc_hd__or2_4
X_23677_ _24317_/CLK _23677_/D VGND VGND VPWR VPWR _23677_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _13252_/A _23915_/Q VGND VGND VPWR VPWR _13432_/B sky130_fd_sc_hd__or2_4
X_25416_ _25409_/CLK _25416_/D HRESETn VGND VGND VPWR VPWR _12676_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_158_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22628_ _16589_/A _21098_/X _21738_/X _22627_/X VGND VGND VPWR VPWR _22628_/X sky130_fd_sc_hd__a211o_4
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _13393_/A _13361_/B _13360_/X VGND VGND VPWR VPWR _13362_/C sky130_fd_sc_hd__and3_4
XFILLER_166_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22559_ _21127_/X VGND VGND VPWR VPWR _22559_/X sky130_fd_sc_hd__buf_2
X_25347_ _25346_/CLK _25347_/D HRESETn VGND VGND VPWR VPWR _12335_/A sky130_fd_sc_hd__dfrtp_4
X_15100_ _24587_/Q VGND VGND VPWR VPWR _15100_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12312_ _24827_/Q VGND VGND VPWR VPWR _12312_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13292_ _13393_/A _13292_/B _13291_/X VGND VGND VPWR VPWR _13292_/X sky130_fd_sc_hd__and3_4
X_16080_ _11699_/A _21587_/A _15920_/X _24713_/Q _16079_/X VGND VGND VPWR VPWR _16080_/X
+ sky130_fd_sc_hd__a32o_4
X_25278_ _23528_/CLK _13755_/X HRESETn VGND VGND VPWR VPWR _14683_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12243_ _23216_/A VGND VGND VPWR VPWR _12243_/Y sky130_fd_sc_hd__inv_2
X_15031_ _15059_/A VGND VGND VPWR VPWR _15245_/A sky130_fd_sc_hd__buf_2
X_24229_ _23398_/CLK _24229_/D HRESETn VGND VGND VPWR VPWR _24229_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15187__C _15242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24671__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12742__B1 _12741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21486__A _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12174_ _12166_/X _12168_/X _12171_/X _12173_/X VGND VGND VPWR VPWR _12174_/X sky130_fd_sc_hd__or4_4
XFILLER_122_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24600__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15484__A _24070_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19770_ _19768_/Y _19764_/X _16869_/X _19769_/X VGND VGND VPWR VPWR _23624_/D sky130_fd_sc_hd__a2bb2o_4
X_16982_ _24375_/Q VGND VGND VPWR VPWR _16982_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18721_ _24153_/Q _18720_/Y VGND VGND VPWR VPWR _18723_/B sky130_fd_sc_hd__or2_4
X_15933_ _12205_/Y _15932_/X _15557_/X _15932_/X VGND VGND VPWR VPWR _15933_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18652_ _18689_/A VGND VGND VPWR VPWR _18769_/A sky130_fd_sc_hd__buf_2
X_15864_ _12808_/Y _15862_/X _15560_/X _15862_/X VGND VGND VPWR VPWR _24813_/D sky130_fd_sc_hd__a2bb2o_4
X_17603_ _17585_/A _17584_/X _17494_/Y _17602_/X VGND VGND VPWR VPWR _17603_/X sky130_fd_sc_hd__or4_4
X_14815_ _14801_/C _14815_/B VGND VGND VPWR VPWR _14815_/Y sky130_fd_sc_hd__nor2_4
XFILLER_92_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18583_ _24163_/Q _18583_/B VGND VGND VPWR VPWR _18583_/X sky130_fd_sc_hd__or2_4
X_15795_ _12352_/Y _15793_/X _15560_/X _15793_/X VGND VGND VPWR VPWR _24848_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_236_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17534_ _17528_/X _17531_/X _17532_/X _17533_/X VGND VGND VPWR VPWR _17554_/A sky130_fd_sc_hd__or4_4
XANTENNA__13732__A _13731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14746_ _14744_/X _14745_/X _14741_/X VGND VGND VPWR VPWR _25063_/D sky130_fd_sc_hd__o21a_4
XFILLER_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11958_ _17479_/C VGND VGND VPWR VPWR _18900_/A sky130_fd_sc_hd__buf_2
XFILLER_45_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17465_ _19208_/B VGND VGND VPWR VPWR _18336_/A sky130_fd_sc_hd__inv_2
XFILLER_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15747__B1 _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14677_ _22056_/A VGND VGND VPWR VPWR _21902_/A sky130_fd_sc_hd__buf_2
X_11889_ _11849_/B _11873_/X VGND VGND VPWR VPWR _11889_/Y sky130_fd_sc_hd__nor2_4
X_19204_ _19202_/Y _19199_/X _19203_/X _19199_/X VGND VGND VPWR VPWR _23820_/D sky130_fd_sc_hd__a2bb2o_4
X_16416_ _16415_/Y _16411_/X _16236_/X _16411_/X VGND VGND VPWR VPWR _24592_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13628_ _12013_/B _13509_/X _13513_/B VGND VGND VPWR VPWR _13629_/B sky130_fd_sc_hd__o21a_4
X_17396_ _17396_/A _17396_/B VGND VGND VPWR VPWR _17399_/B sky130_fd_sc_hd__or2_4
X_19135_ _23844_/Q VGND VGND VPWR VPWR _19135_/Y sky130_fd_sc_hd__inv_2
X_16347_ _16346_/Y _16344_/X _16062_/X _16344_/X VGND VGND VPWR VPWR _16347_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15659__A _15666_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13559_ _13559_/A VGND VGND VPWR VPWR _13559_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24759__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19066_ HWDATA[1] VGND VGND VPWR VPWR _19360_/A sky130_fd_sc_hd__buf_2
XFILLER_157_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16278_ _16318_/A VGND VGND VPWR VPWR _16278_/X sky130_fd_sc_hd__buf_2
X_18017_ _18017_/A VGND VGND VPWR VPWR _18097_/A sky130_fd_sc_hd__buf_2
X_15229_ _15229_/A _15229_/B VGND VGND VPWR VPWR _15230_/C sky130_fd_sc_hd__or2_4
XFILLER_173_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19110__B1 _19063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21396__A _22197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24341__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19968_ _22247_/B _19963_/X _19967_/X _19963_/X VGND VGND VPWR VPWR _23553_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18919_ _18917_/Y _18913_/X _17421_/X _18918_/X VGND VGND VPWR VPWR _23920_/D sky130_fd_sc_hd__a2bb2o_4
X_19899_ _19898_/X VGND VGND VPWR VPWR _19900_/A sky130_fd_sc_hd__inv_2
XFILLER_67_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21930_ _21920_/A VGND VGND VPWR VPWR _22015_/A sky130_fd_sc_hd__buf_2
XANTENNA__21843__B _21843_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21861_ _21323_/A VGND VGND VPWR VPWR _23088_/B sky130_fd_sc_hd__buf_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14789__A1 _13579_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14789__B2 _14611_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20812_ _20690_/X _20811_/Y _15559_/A _20735_/X VGND VGND VPWR VPWR _24031_/D sky130_fd_sc_hd__a2bb2o_4
X_23600_ _23528_/CLK _19841_/X VGND VGND VPWR VPWR _23600_/Q sky130_fd_sc_hd__dfxtp_4
X_21792_ _21487_/A _21792_/B VGND VGND VPWR VPWR _21792_/X sky130_fd_sc_hd__or2_4
X_24580_ _24591_/CLK _24580_/D HRESETn VGND VGND VPWR VPWR _24580_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22720__A1 _16128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22720__B2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20743_ _20731_/X _20742_/Y _24905_/Q _20736_/X VGND VGND VPWR VPWR _24015_/D sky130_fd_sc_hd__a2bb2o_4
X_23531_ _24302_/CLK _20030_/X VGND VGND VPWR VPWR _20029_/A sky130_fd_sc_hd__dfxtp_4
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23462_ _23464_/CLK _20211_/X VGND VGND VPWR VPWR _18107_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_211_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20674_ _20678_/A _20515_/B VGND VGND VPWR VPWR _20674_/X sky130_fd_sc_hd__or2_4
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22413_ _22279_/X _22412_/X _21306_/C _24723_/Q _22282_/X VGND VGND VPWR VPWR _22413_/X
+ sky130_fd_sc_hd__a32o_4
X_25201_ _25056_/CLK _14214_/X HRESETn VGND VGND VPWR VPWR _25201_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23393_ _23932_/CLK _23393_/D VGND VGND VPWR VPWR _23393_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23229__A2_N _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22344_ _21926_/A _22344_/B VGND VGND VPWR VPWR _22344_/X sky130_fd_sc_hd__or2_4
X_25132_ _25117_/CLK _14438_/X HRESETn VGND VGND VPWR VPWR _25132_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_136_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24429__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25063_ _23494_/CLK _25063_/D HRESETn VGND VGND VPWR VPWR _14705_/A sky130_fd_sc_hd__dfrtp_4
X_22275_ _21441_/X VGND VGND VPWR VPWR _22275_/X sky130_fd_sc_hd__buf_2
XFILLER_191_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24014_ _24049_/CLK _20740_/X HRESETn VGND VGND VPWR VPWR _20738_/A sky130_fd_sc_hd__dfrtp_4
X_21226_ _22829_/A VGND VGND VPWR VPWR _22794_/A sky130_fd_sc_hd__buf_2
XFILLER_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21157_ _21156_/Y _21348_/A _14876_/Y _14422_/A VGND VGND VPWR VPWR _21157_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24011__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20108_ _23500_/Q VGND VGND VPWR VPWR _21397_/B sky130_fd_sc_hd__inv_2
X_21088_ _21088_/A _22420_/B VGND VGND VPWR VPWR _21096_/B sky130_fd_sc_hd__or2_4
XFILLER_59_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12930_ _12807_/X _12929_/X VGND VGND VPWR VPWR _12947_/B sky130_fd_sc_hd__or2_4
X_20039_ _20034_/A VGND VGND VPWR VPWR _20039_/X sky130_fd_sc_hd__buf_2
X_24916_ _24508_/CLK _24916_/D HRESETn VGND VGND VPWR VPWR _15574_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_219_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25288__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ _12861_/A _12861_/B _12860_/X VGND VGND VPWR VPWR _12861_/X sky130_fd_sc_hd__and3_4
X_24847_ _25341_/CLK _24847_/D HRESETn VGND VGND VPWR VPWR _24847_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15977__B1 _15976_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19168__B1 _19122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14600_ _14550_/B _14599_/X _14546_/X _14591_/X _25084_/Q VGND VGND VPWR VPWR _14600_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11810_/Y _11808_/A _25296_/Q _22735_/A VGND VGND VPWR VPWR _11813_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _24914_/Q VGND VGND VPWR VPWR _15580_/Y sky130_fd_sc_hd__inv_2
XPHY_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12782_/X _12792_/B _12788_/X _12792_/D VGND VGND VPWR VPWR _12792_/X sky130_fd_sc_hd__or4_4
X_24778_ _25380_/CLK _24778_/D HRESETn VGND VGND VPWR VPWR _23275_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22865__A _21127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22711__A1 _24730_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14524_/Y _14061_/Y _20453_/C VGND VGND VPWR VPWR _14531_/X sky130_fd_sc_hd__o21a_4
XFILLER_214_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _16236_/A VGND VGND VPWR VPWR _11743_/X sky130_fd_sc_hd__buf_2
X_23729_ _23406_/CLK _19461_/X VGND VGND VPWR VPWR _19460_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__15729__B1 _15581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _24357_/Q VGND VGND VPWR VPWR _17314_/C sky130_fd_sc_hd__inv_2
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14462_/A _14442_/B VGND VGND VPWR VPWR _14468_/A sky130_fd_sc_hd__nor2_4
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11674_/A _13765_/A _15640_/B _15640_/C VGND VGND VPWR VPWR _16446_/D sky130_fd_sc_hd__or4_4
XANTENNA__14401__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23267__A2 _22718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_140_0_HCLK clkbuf_7_70_0_HCLK/X VGND VGND VPWR VPWR _23873_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15744__A3 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ _16200_/Y _16198_/X _11685_/X _16198_/X VGND VGND VPWR VPWR _16201_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_230_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _13445_/A _19756_/A VGND VGND VPWR VPWR _13415_/B sky130_fd_sc_hd__or2_4
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17181_ _24349_/Q VGND VGND VPWR VPWR _17243_/B sky130_fd_sc_hd__inv_2
X_14393_ _14391_/Y _14372_/X _14392_/X _14372_/X VGND VGND VPWR VPWR _14393_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14383__A _14083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24852__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16132_ _16131_/Y _16129_/X _11739_/X _16129_/X VGND VGND VPWR VPWR _24694_/D sky130_fd_sc_hd__a2bb2o_4
X_13344_ _13268_/X _13344_/B _13343_/X VGND VGND VPWR VPWR _13344_/X sky130_fd_sc_hd__and3_4
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16063_ _16061_/Y _16058_/X _16062_/X _16058_/X VGND VGND VPWR VPWR _24721_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13275_ _13312_/A _13275_/B VGND VGND VPWR VPWR _13275_/X sky130_fd_sc_hd__or2_4
X_15014_ _24459_/Q VGND VGND VPWR VPWR _15014_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12226_ _12273_/B VGND VGND VPWR VPWR _12226_/X sky130_fd_sc_hd__buf_2
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12157_ _12111_/Y _12156_/Y SCLK_S3 _12155_/X VGND VGND VPWR VPWR _12157_/X sky130_fd_sc_hd__o22a_4
X_19822_ _23605_/Q VGND VGND VPWR VPWR _21605_/B sky130_fd_sc_hd__inv_2
XFILLER_123_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12088_ _13483_/A _12086_/X _12058_/C _12087_/X VGND VGND VPWR VPWR _12089_/A sky130_fd_sc_hd__or4_4
X_16965_ _16965_/A VGND VGND VPWR VPWR _16965_/Y sky130_fd_sc_hd__inv_2
X_19753_ _19753_/A VGND VGND VPWR VPWR _19753_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15916_ _15771_/B _15918_/B VGND VGND VPWR VPWR _15916_/X sky130_fd_sc_hd__or2_4
X_18704_ _18734_/A _18704_/B _18704_/C VGND VGND VPWR VPWR _18704_/X sky130_fd_sc_hd__and3_4
XFILLER_77_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15942__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19684_ _13372_/B VGND VGND VPWR VPWR _19684_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19414__A _19006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16896_ _22564_/A _16895_/X _16098_/Y _24284_/Q VGND VGND VPWR VPWR _16901_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18635_ _24128_/Q VGND VGND VPWR VPWR _18819_/A sky130_fd_sc_hd__inv_2
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15847_ _21579_/B VGND VGND VPWR VPWR _22816_/A sky130_fd_sc_hd__buf_2
XFILLER_237_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19159__B1 _19067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18566_ _18409_/Y _18566_/B VGND VGND VPWR VPWR _18567_/B sky130_fd_sc_hd__or2_4
X_15778_ _13454_/A _13453_/A _11660_/A _15984_/D VGND VGND VPWR VPWR _15778_/X sky130_fd_sc_hd__or4_4
XFILLER_80_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18906__B1 HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17517_ _24112_/Q VGND VGND VPWR VPWR _17517_/Y sky130_fd_sc_hd__inv_2
X_14729_ _14729_/A VGND VGND VPWR VPWR _22048_/A sky130_fd_sc_hd__inv_2
XFILLER_220_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18497_ _18497_/A _18497_/B _18497_/C VGND VGND VPWR VPWR _24187_/D sky130_fd_sc_hd__and3_4
XFILLER_177_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22494__B _22654_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17448_ _17448_/A VGND VGND VPWR VPWR _18910_/B sky130_fd_sc_hd__buf_2
XFILLER_220_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23258__A2 _21597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17379_ _17203_/X _17344_/B VGND VGND VPWR VPWR _17379_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24593__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19118_ _19117_/X VGND VGND VPWR VPWR _19133_/A sky130_fd_sc_hd__inv_2
XFILLER_229_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20390_ _20386_/Y _20389_/X _18250_/X _20389_/X VGND VGND VPWR VPWR _23392_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24522__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19049_ _19054_/A VGND VGND VPWR VPWR _19049_/X sky130_fd_sc_hd__buf_2
XFILLER_173_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22501__A1_N _17358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22060_ _21627_/A VGND VGND VPWR VPWR _22373_/A sky130_fd_sc_hd__buf_2
XFILLER_161_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21011_ sda_oen_o_S5 _24950_/Q _21006_/A _15422_/A _21010_/Y VGND VGND VPWR VPWR
+ _21011_/X sky130_fd_sc_hd__a32o_4
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23194__A1 _22552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15852__A _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23194__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25381__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22962_ _22761_/X _22960_/X _22691_/X _22961_/X VGND VGND VPWR VPWR _22962_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22941__A1 _16569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24701_ _24696_/CLK _24701_/D HRESETn VGND VGND VPWR VPWR _24701_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21913_ _21913_/A _20074_/Y VGND VGND VPWR VPWR _21913_/X sky130_fd_sc_hd__or2_4
XANTENNA__11693__B1 _11691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25310__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15959__B1 _24763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22893_ _14908_/A _22807_/X _21737_/X _22892_/X VGND VGND VPWR VPWR _22894_/C sky130_fd_sc_hd__a211o_4
XANTENNA__14468__A _14468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24632_ _24629_/CLK _24632_/D HRESETn VGND VGND VPWR VPWR _22944_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_243_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16620__B2 _16541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21844_ _16610_/A _21325_/X _23001_/A _21843_/X VGND VGND VPWR VPWR _21845_/C sky130_fd_sc_hd__a211o_4
XFILLER_231_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15974__A3 _15830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14187__B _14187_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21775_ _21775_/A _21775_/B VGND VGND VPWR VPWR _21777_/B sky130_fd_sc_hd__or2_4
X_24563_ _24540_/CLK _16497_/X HRESETn VGND VGND VPWR VPWR _16494_/A sky130_fd_sc_hd__dfrtp_4
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20726_ _20725_/X VGND VGND VPWR VPWR _20726_/Y sky130_fd_sc_hd__inv_2
X_23514_ _24199_/CLK _20068_/X VGND VGND VPWR VPWR _23514_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24494_ _24051_/CLK _24494_/D HRESETn VGND VGND VPWR VPWR _16679_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_23_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15726__A3 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_213_0_HCLK clkbuf_7_106_0_HCLK/X VGND VGND VPWR VPWR _24060_/CLK sky130_fd_sc_hd__clkbuf_1
X_20657_ _17394_/B _20657_/B _20661_/C VGND VGND VPWR VPWR _20657_/X sky130_fd_sc_hd__and3_4
X_23445_ _23499_/CLK _20256_/X VGND VGND VPWR VPWR _20254_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21710__A1_N _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23376_ _25346_/CLK HSEL VGND VGND VPWR VPWR _23339_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_139_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12231__A2_N _24761_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20588_ _23947_/Q _18881_/B VGND VGND VPWR VPWR _20589_/B sky130_fd_sc_hd__nand2_4
XANTENNA__24263__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25115_ _24326_/CLK _14480_/X HRESETn VGND VGND VPWR VPWR _14477_/A sky130_fd_sc_hd__dfrtp_4
X_22327_ _15456_/Y _22327_/B VGND VGND VPWR VPWR _22327_/Y sky130_fd_sc_hd__nor2_4
XFILLER_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13060_ _12985_/B _13059_/X VGND VGND VPWR VPWR _13063_/B sky130_fd_sc_hd__or2_4
X_22258_ _22261_/A _22258_/B VGND VGND VPWR VPWR _22258_/X sky130_fd_sc_hd__or2_4
X_25046_ _25050_/CLK _14855_/X HRESETn VGND VGND VPWR VPWR _14809_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_151_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12011_ _12009_/Y _12010_/X _12009_/Y _12010_/X VGND VGND VPWR VPWR _12012_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21209_ _21209_/A _21209_/B VGND VGND VPWR VPWR _21210_/C sky130_fd_sc_hd__or2_4
XFILLER_133_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17019__A _24403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22189_ _22189_/A VGND VGND VPWR VPWR _22194_/A sky130_fd_sc_hd__buf_2
XANTENNA__12451__A _12418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16750_ _16748_/Y _16745_/X _16397_/X _16749_/X VGND VGND VPWR VPWR _16750_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15762__A _11774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13962_ _13962_/A _13961_/X VGND VGND VPWR VPWR _13962_/X sky130_fd_sc_hd__or2_4
XFILLER_171_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21735__A2 _21728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15701_ _15700_/X VGND VGND VPWR VPWR _15701_/X sky130_fd_sc_hd__buf_2
XFILLER_58_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12913_ _12912_/X VGND VGND VPWR VPWR _12914_/B sky130_fd_sc_hd__inv_2
XANTENNA__25051__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16681_ _16679_/Y _16680_/X _15739_/X _16680_/X VGND VGND VPWR VPWR _24494_/D sky130_fd_sc_hd__a2bb2o_4
X_13893_ _13935_/B VGND VGND VPWR VPWR _13943_/D sky130_fd_sc_hd__inv_2
X_18420_ _18420_/A VGND VGND VPWR VPWR _18420_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15632_ _24894_/Q VGND VGND VPWR VPWR _15632_/Y sky130_fd_sc_hd__inv_2
X_12844_ _12617_/B _12851_/A VGND VGND VPWR VPWR _12857_/B sky130_fd_sc_hd__or2_4
XFILLER_203_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18351_ _18350_/Y _17476_/X _18350_/A _17480_/X VGND VGND VPWR VPWR _18365_/A sky130_fd_sc_hd__o22a_4
XFILLER_221_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15563_ _15563_/A VGND VGND VPWR VPWR _15563_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12775_ _25370_/Q VGND VGND VPWR VPWR _12775_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_23_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17301_/X VGND VGND VPWR VPWR _24363_/D sky130_fd_sc_hd__inv_2
XANTENNA__22160__A2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14514_ _14510_/X _14513_/X _25118_/Q _14506_/X VGND VGND VPWR VPWR _25106_/D sky130_fd_sc_hd__o22a_4
XFILLER_42_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ HWDATA[16] VGND VGND VPWR VPWR _11726_/X sky130_fd_sc_hd__buf_2
X_18282_ _18282_/A VGND VGND VPWR VPWR _18285_/B sky130_fd_sc_hd__buf_2
XFILLER_159_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15489_/A VGND VGND VPWR VPWR _15494_/X sky130_fd_sc_hd__buf_2
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16914__A2 _16913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17233_ _24367_/Q VGND VGND VPWR VPWR _17255_/A sky130_fd_sc_hd__inv_2
X_14445_ _20539_/A VGND VGND VPWR VPWR _14445_/Y sky130_fd_sc_hd__inv_2
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _15636_/B VGND VGND VPWR VPWR _14178_/B sky130_fd_sc_hd__buf_2
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17164_ _16275_/Y _17261_/A _16275_/Y _17261_/A VGND VGND VPWR VPWR _17164_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16127__B1 _11730_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _14375_/Y _14371_/X _13826_/X _14373_/X VGND VGND VPWR VPWR _14376_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17416__A1_N _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16115_ _22909_/A VGND VGND VPWR VPWR _16115_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13327_ _13391_/A _23814_/Q VGND VGND VPWR VPWR _13329_/B sky130_fd_sc_hd__or2_4
X_17095_ _17004_/Y _17090_/B _17064_/X _17091_/Y VGND VGND VPWR VPWR _17095_/X sky130_fd_sc_hd__a211o_4
XFILLER_182_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16046_ _16044_/Y _16045_/X _11748_/X _16045_/X VGND VGND VPWR VPWR _24727_/D sky130_fd_sc_hd__a2bb2o_4
X_13258_ _13365_/A _13256_/X _13257_/X VGND VGND VPWR VPWR _13262_/B sky130_fd_sc_hd__and3_4
XANTENNA__23986__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12209_ _22476_/A VGND VGND VPWR VPWR _12209_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13189_ _13189_/A VGND VGND VPWR VPWR _13285_/A sky130_fd_sc_hd__buf_2
XFILLER_69_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19805_ _19805_/A VGND VGND VPWR VPWR _19805_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17997_ _17947_/A _17997_/B _17996_/X VGND VGND VPWR VPWR _17997_/X sky130_fd_sc_hd__and3_4
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19144__A _19006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16948_ _16943_/X _16944_/X _16948_/C _16947_/X VGND VGND VPWR VPWR _16948_/X sky130_fd_sc_hd__or4_4
X_19736_ _19735_/Y _19731_/X _19646_/X _19723_/A VGND VGND VPWR VPWR _19736_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21726__A2 _14182_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_105_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_211_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16879_ _16876_/Y _16877_/X _16878_/X _16877_/X VGND VGND VPWR VPWR _24408_/D sky130_fd_sc_hd__a2bb2o_4
X_19667_ _19666_/Y _19664_/X _19543_/X _19664_/X VGND VGND VPWR VPWR _19667_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11705__A _22807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18618_ _18608_/X _18618_/B _18618_/C _18618_/D VGND VGND VPWR VPWR _18638_/B sky130_fd_sc_hd__or4_4
X_19598_ _19598_/A VGND VGND VPWR VPWR _19598_/Y sky130_fd_sc_hd__inv_2
XFILLER_241_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18549_ _18465_/Y _18524_/X _18500_/X _18547_/B VGND VGND VPWR VPWR _18549_/X sky130_fd_sc_hd__a211o_4
XFILLER_212_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24774__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21560_ _21559_/Y _21159_/X _14863_/Y _21365_/X VGND VGND VPWR VPWR _21561_/A sky130_fd_sc_hd__o22a_4
XFILLER_21_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24703__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15708__A3 _15702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20511_ _24077_/Q _20510_/X _14271_/X VGND VGND VPWR VPWR _20514_/B sky130_fd_sc_hd__o21a_4
XANTENNA__22439__B1 _12306_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21491_ _21654_/A _19472_/Y VGND VGND VPWR VPWR _21493_/B sky130_fd_sc_hd__or2_4
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19304__B1 _19279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23230_ _17231_/X _22485_/X _12828_/A _22444_/X VGND VGND VPWR VPWR _23231_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20442_ _20603_/A _20441_/Y VGND VGND VPWR VPWR _20461_/A sky130_fd_sc_hd__and2_4
XFILLER_146_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21849__A _14182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14965__A2_N _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23161_ _12278_/A _22984_/X _24284_/Q _22914_/X VGND VGND VPWR VPWR _23161_/X sky130_fd_sc_hd__a2bb2o_4
X_20373_ _20372_/X _20368_/X _13826_/A _23400_/Q _20370_/X VGND VGND VPWR VPWR _20373_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15847__A _21579_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_43_0_HCLK clkbuf_8_43_0_HCLK/A VGND VGND VPWR VPWR _24209_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_109_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21568__B _21568_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22112_ _12781_/Y _21019_/X _20847_/Y _22111_/X VGND VGND VPWR VPWR _22112_/X sky130_fd_sc_hd__o22a_4
X_23092_ _22824_/X _23083_/Y _23087_/Y _23091_/X VGND VGND VPWR VPWR _23092_/X sky130_fd_sc_hd__a211o_4
XFILLER_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22043_ _22043_/A _19592_/Y VGND VGND VPWR VPWR _22043_/X sky130_fd_sc_hd__or2_4
XFILLER_133_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23994_ _23972_/CLK _23994_/D HRESETn VGND VGND VPWR VPWR _23994_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21717__A2 _14212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22945_ _24736_/Q _21061_/X _21062_/X _22944_/X VGND VGND VPWR VPWR _22945_/X sky130_fd_sc_hd__a211o_4
XFILLER_216_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22876_ _22874_/X _22875_/X _22876_/C VGND VGND VPWR VPWR _22876_/X sky130_fd_sc_hd__or3_4
XANTENNA__22127__C1 _22101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24615_ _24662_/CLK _16354_/X HRESETn VGND VGND VPWR VPWR _24615_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21827_ _22393_/A _21827_/B _21827_/C VGND VGND VPWR VPWR _21827_/X sky130_fd_sc_hd__and3_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15834__A1_N _12332_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _12560_/A VGND VGND VPWR VPWR _12608_/A sky130_fd_sc_hd__inv_2
X_24546_ _24080_/CLK _24546_/D HRESETn VGND VGND VPWR VPWR _24546_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12091__B1 _11753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21758_ _21754_/X _21757_/X _14707_/X VGND VGND VPWR VPWR _21758_/X sky130_fd_sc_hd__o21a_4
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24444__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20709_ _20709_/A VGND VGND VPWR VPWR _20709_/Y sky130_fd_sc_hd__inv_2
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12480_/A _12491_/B _12490_/Y VGND VGND VPWR VPWR _25435_/D sky130_fd_sc_hd__and3_4
X_24477_ _24477_/CLK _16727_/X HRESETn VGND VGND VPWR VPWR _24477_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21689_ _21668_/X _21688_/X _21501_/X VGND VGND VPWR VPWR _21689_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_196_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _14229_/Y _14225_/X _13798_/X _14213_/A VGND VGND VPWR VPWR _14230_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23428_ _23427_/CLK _20301_/X VGND VGND VPWR VPWR _20299_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16109__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21653__A1 _21641_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14161_ _14161_/A VGND VGND VPWR VPWR _14161_/X sky130_fd_sc_hd__buf_2
X_23359_ VGND VGND VPWR VPWR _23359_/HI sda_o_S5 sky130_fd_sc_hd__conb_1
XFILLER_124_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22850__B1 _12547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13112_ _13112_/A VGND VGND VPWR VPWR _13113_/B sky130_fd_sc_hd__inv_2
XFILLER_125_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14092_ _14092_/A _14092_/B _25223_/Q VGND VGND VPWR VPWR _14092_/X sky130_fd_sc_hd__or3_4
XFILLER_180_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12185__A2_N _21088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13043_ _12302_/Y _13048_/B _13019_/X VGND VGND VPWR VPWR _13043_/Y sky130_fd_sc_hd__a21oi_4
X_17920_ _17914_/Y _13528_/X _17917_/Y _17914_/A _17919_/X VGND VGND VPWR VPWR _24253_/D
+ sky130_fd_sc_hd__a32o_4
X_25029_ _25028_/CLK _15211_/X HRESETn VGND VGND VPWR VPWR _14898_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17851_ _17753_/D _17850_/X VGND VGND VPWR VPWR _17852_/B sky130_fd_sc_hd__or2_4
XFILLER_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21494__A _21463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16802_ _14900_/Y _16799_/X _16467_/X _16799_/X VGND VGND VPWR VPWR _24441_/D sky130_fd_sc_hd__a2bb2o_4
X_17782_ _17790_/A _17782_/B _17782_/C VGND VGND VPWR VPWR _17782_/X sky130_fd_sc_hd__and3_4
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14994_ _14976_/X _16781_/A _14976_/X _16781_/A VGND VGND VPWR VPWR _14997_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21169__B1 _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22102__B _21849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16733_ _16732_/Y _16730_/X _16464_/X _16730_/X VGND VGND VPWR VPWR _16733_/X sky130_fd_sc_hd__a2bb2o_4
X_19521_ _23706_/Q VGND VGND VPWR VPWR _19521_/Y sky130_fd_sc_hd__inv_2
X_13945_ _13914_/X VGND VGND VPWR VPWR _13947_/A sky130_fd_sc_hd__inv_2
XFILLER_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19452_ _19451_/Y _19447_/X _19408_/X _19447_/A VGND VGND VPWR VPWR _19452_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16664_ _16663_/Y _16661_/X _16391_/X _16661_/X VGND VGND VPWR VPWR _24501_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13876_ _13876_/A VGND VGND VPWR VPWR _14232_/C sky130_fd_sc_hd__buf_2
XFILLER_234_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15938__A3 HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15615_ _24900_/Q VGND VGND VPWR VPWR _15615_/Y sky130_fd_sc_hd__inv_2
X_18403_ _24185_/Q VGND VGND VPWR VPWR _18505_/A sky130_fd_sc_hd__inv_2
X_12827_ _12967_/A VGND VGND VPWR VPWR _12861_/A sky130_fd_sc_hd__buf_2
X_19383_ _19382_/Y _19380_/X _19360_/X _19380_/X VGND VGND VPWR VPWR _23756_/D sky130_fd_sc_hd__a2bb2o_4
X_16595_ _16594_/Y _16592_/X _16420_/X _16592_/X VGND VGND VPWR VPWR _24525_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_222_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23330__A1 _24578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18334_ _18910_/B _17485_/A _19094_/B _18326_/B VGND VGND VPWR VPWR _24209_/D sky130_fd_sc_hd__o22a_4
X_15546_ _11678_/X VGND VGND VPWR VPWR _16637_/A sky130_fd_sc_hd__buf_2
X_12758_ _12755_/A _24793_/Q _12756_/X _12757_/Y VGND VGND VPWR VPWR _12765_/B sky130_fd_sc_hd__o22a_4
XFILLER_15_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24185__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11709_ _11699_/X _11707_/X HWDATA[21] _25541_/Q _11708_/X VGND VGND VPWR VPWR _25541_/D
+ sky130_fd_sc_hd__a32o_4
X_18265_ _18264_/X VGND VGND VPWR VPWR _18265_/Y sky130_fd_sc_hd__inv_2
X_15477_ _24950_/Q _15433_/X _15430_/X VGND VGND VPWR VPWR _24950_/D sky130_fd_sc_hd__a21bo_4
XANTENNA__24114__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12689_ _12689_/A _12592_/Y VGND VGND VPWR VPWR _12716_/B sky130_fd_sc_hd__or2_4
XFILLER_202_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17216_ _16348_/Y _21856_/A _24640_/Q _17215_/Y VGND VGND VPWR VPWR _17221_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_175_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14428_ _14428_/A VGND VGND VPWR VPWR _14428_/Y sky130_fd_sc_hd__inv_2
X_18196_ _18132_/A _18196_/B _18196_/C VGND VGND VPWR VPWR _18196_/X sky130_fd_sc_hd__and3_4
XANTENNA__22436__A3 _22432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17147_ _16991_/A _17147_/B VGND VGND VPWR VPWR _17148_/B sky130_fd_sc_hd__or2_4
X_14359_ _25155_/Q _14338_/B _25154_/Q _14345_/A VGND VGND VPWR VPWR _14359_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_2_0_HCLK clkbuf_8_3_0_HCLK/A VGND VGND VPWR VPWR _23859_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_144_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17078_ _17026_/A _17076_/X _17077_/Y VGND VGND VPWR VPWR _17078_/X sky130_fd_sc_hd__o21a_4
X_16029_ _24733_/Q VGND VGND VPWR VPWR _16029_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19719_ _19715_/Y _19718_/X _19652_/X _19718_/X VGND VGND VPWR VPWR _19719_/X sky130_fd_sc_hd__a2bb2o_4
X_20991_ _23930_/Q _23931_/Q _20990_/Y VGND VGND VPWR VPWR _20991_/X sky130_fd_sc_hd__o21a_4
XFILLER_226_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22730_ _22730_/A VGND VGND VPWR VPWR _22730_/X sky130_fd_sc_hd__buf_2
XFILLER_53_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21580__B1 _21582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15929__A3 _15710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23124__A _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22661_ _22145_/B VGND VGND VPWR VPWR _22661_/X sky130_fd_sc_hd__buf_2
XFILLER_53_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18218__A _18014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24400_ _24390_/CLK _24400_/D HRESETn VGND VGND VPWR VPWR _16965_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21612_ _21757_/A _21610_/X _21612_/C VGND VGND VPWR VPWR _21612_/X sky130_fd_sc_hd__and3_4
XFILLER_179_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25380_ _25380_/CLK _12926_/Y HRESETn VGND VGND VPWR VPWR _25380_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12073__B1 _11786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22592_ _16591_/A _21098_/X _21738_/X _22591_/X VGND VGND VPWR VPWR _22592_/X sky130_fd_sc_hd__a211o_4
XFILLER_194_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24331_ _24980_/CLK _24331_/D HRESETn VGND VGND VPWR VPWR _24331_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21543_ _22279_/A _21540_/X _21541_/X _24718_/Q _21542_/X VGND VGND VPWR VPWR _21543_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25405__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21474_ _21665_/A _21474_/B VGND VGND VPWR VPWR _21474_/X sky130_fd_sc_hd__or2_4
X_24262_ _24263_/CLK _17879_/Y HRESETn VGND VGND VPWR VPWR _24262_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21579__A _15005_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20425_ _21396_/B _20422_/X _19827_/A _20422_/X VGND VGND VPWR VPWR _20425_/X sky130_fd_sc_hd__a2bb2o_4
X_23213_ _23213_/A _23210_/X _23213_/C VGND VGND VPWR VPWR _23214_/D sky130_fd_sc_hd__and3_4
X_24193_ _25471_/CLK _18387_/X HRESETn VGND VGND VPWR VPWR _24193_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20356_ _22033_/B _20350_/X _19606_/A _20355_/X VGND VGND VPWR VPWR _23407_/D sky130_fd_sc_hd__a2bb2o_4
X_23144_ _23144_/A _22897_/X VGND VGND VPWR VPWR _23144_/X sky130_fd_sc_hd__or2_4
XANTENNA__16511__B1 _16420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23075_ _24571_/Q _23075_/B _23075_/C VGND VGND VPWR VPWR _23075_/X sky130_fd_sc_hd__and3_4
X_20287_ _20286_/X VGND VGND VPWR VPWR _20287_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22026_ _21670_/X _22026_/B VGND VGND VPWR VPWR _22026_/X sky130_fd_sc_hd__or2_4
XFILLER_248_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11991_ _24093_/Q _11977_/X _11990_/Y VGND VGND VPWR VPWR _11992_/A sky130_fd_sc_hd__o21a_4
X_23977_ _23976_/CLK _20627_/Y HRESETn VGND VGND VPWR VPWR _23977_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24696__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12300__B2 _24820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13730_ _13730_/A _13729_/Y VGND VGND VPWR VPWR _14775_/A sky130_fd_sc_hd__or2_4
XFILLER_17_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22928_ _22928_/A VGND VGND VPWR VPWR _22928_/X sky130_fd_sc_hd__buf_2
XFILLER_205_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24625__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23034__A _23011_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13661_ _25298_/Q _13510_/X _13660_/Y VGND VGND VPWR VPWR _25298_/D sky130_fd_sc_hd__o21a_4
XFILLER_232_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22859_ _22474_/X _22857_/X _22858_/X _24838_/Q _22478_/X VGND VGND VPWR VPWR _22859_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_231_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15400_ _15379_/A _15400_/B _15399_/Y VGND VGND VPWR VPWR _24983_/D sky130_fd_sc_hd__and3_4
XFILLER_231_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12612_ _12614_/B VGND VGND VPWR VPWR _12613_/B sky130_fd_sc_hd__inv_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16380_ _24606_/Q VGND VGND VPWR VPWR _16380_/Y sky130_fd_sc_hd__inv_2
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13592_ _14628_/A _13592_/B VGND VGND VPWR VPWR _13593_/A sky130_fd_sc_hd__and2_4
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15331_ _15331_/A _15331_/B _15137_/Y _15301_/A VGND VGND VPWR VPWR _15339_/A sky130_fd_sc_hd__or4_4
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12543_ _24873_/Q VGND VGND VPWR VPWR _12543_/Y sky130_fd_sc_hd__inv_2
X_24529_ _24558_/CLK _24529_/D HRESETn VGND VGND VPWR VPWR _24529_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18050_ _18123_/A _18050_/B _18050_/C VGND VGND VPWR VPWR _18050_/X sky130_fd_sc_hd__and3_4
X_15262_ _15265_/A _15269_/B VGND VGND VPWR VPWR _15266_/B sky130_fd_sc_hd__or2_4
XFILLER_200_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12474_ _12474_/A VGND VGND VPWR VPWR _12474_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16750__B1 _16397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17001_ _16016_/Y _24395_/Q _24726_/Q _17038_/D VGND VGND VPWR VPWR _17008_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14213_ _14213_/A VGND VGND VPWR VPWR _14213_/X sky130_fd_sc_hd__buf_2
XFILLER_138_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12367__B2 _24823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15193_ _15165_/A _15191_/X _15192_/X VGND VGND VPWR VPWR _25033_/D sky130_fd_sc_hd__and3_4
XANTENNA__25484__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12904__A _12838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14144_ _14135_/X _14143_/Y _25137_/Q _14135_/X VGND VGND VPWR VPWR _14144_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16502__B1 _16229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24922__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14075_ _24001_/Q _14067_/A _14062_/X _14008_/A _14073_/X VGND VGND VPWR VPWR _14075_/X
+ sky130_fd_sc_hd__a32o_4
X_18952_ _18950_/Y _18947_/X _18951_/X _18947_/X VGND VGND VPWR VPWR _18952_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_180_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13026_ _12970_/X _13017_/X _13025_/X VGND VGND VPWR VPWR _25358_/D sky130_fd_sc_hd__and3_4
X_17903_ _17893_/Y _17906_/A VGND VGND VPWR VPWR _17903_/X sky130_fd_sc_hd__and2_4
XFILLER_79_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18883_ _23949_/Q _20593_/A VGND VGND VPWR VPWR _18884_/A sky130_fd_sc_hd__or2_4
XFILLER_121_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17834_ _17833_/X VGND VGND VPWR VPWR _17835_/B sky130_fd_sc_hd__inv_2
XFILLER_239_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18270__A3 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18653__A1_N _16582_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14977_ _15265_/A _14885_/A _14976_/X _16847_/A VGND VGND VPWR VPWR _14977_/X sky130_fd_sc_hd__a2bb2o_4
X_17765_ _17743_/Y _17764_/X VGND VGND VPWR VPWR _17786_/B sky130_fd_sc_hd__or2_4
XANTENNA__19755__B1 _19708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19504_ _22351_/B _19503_/X _11902_/X _19503_/X VGND VGND VPWR VPWR _23714_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13928_ _13914_/X _13928_/B _13923_/D _13879_/X VGND VGND VPWR VPWR _13928_/X sky130_fd_sc_hd__or4_4
X_16716_ _16361_/A VGND VGND VPWR VPWR _16716_/X sky130_fd_sc_hd__buf_2
XFILLER_81_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17696_ _17521_/Y _17696_/B VGND VGND VPWR VPWR _17696_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24366__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16647_ _24507_/Q VGND VGND VPWR VPWR _16647_/Y sky130_fd_sc_hd__inv_2
X_19435_ _19447_/A VGND VGND VPWR VPWR _19435_/X sky130_fd_sc_hd__buf_2
XFILLER_222_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13859_ _13841_/X _13858_/X _25191_/Q _13856_/X VGND VGND VPWR VPWR _13859_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22106__A2 _21349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23303__A1 _16796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16578_ _16578_/A VGND VGND VPWR VPWR _16578_/Y sky130_fd_sc_hd__inv_2
X_19366_ _19365_/X VGND VGND VPWR VPWR _19372_/A sky130_fd_sc_hd__buf_2
X_15529_ _16446_/C _15524_/X HADDR[5] _15524_/X VGND VGND VPWR VPWR _15529_/X sky130_fd_sc_hd__a2bb2o_4
X_18317_ _18296_/X _18316_/Y _18298_/B _18315_/X VGND VGND VPWR VPWR _18317_/X sky130_fd_sc_hd__o22a_4
XFILLER_148_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21865__A1 _24418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19297_ _17951_/B VGND VGND VPWR VPWR _19297_/Y sky130_fd_sc_hd__inv_2
X_18248_ _18238_/X _18240_/X _16597_/X _22517_/A _18241_/X VGND VGND VPWR VPWR _18248_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_148_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18179_ _17968_/X _18177_/X _18179_/C VGND VGND VPWR VPWR _18179_/X sky130_fd_sc_hd__and3_4
XFILLER_191_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20210_ _18107_/B VGND VGND VPWR VPWR _20210_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16931__A2_N _17744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23930__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21190_ _21209_/A _21190_/B VGND VGND VPWR VPWR _21190_/X sky130_fd_sc_hd__or2_4
XANTENNA__25154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20141_ _20140_/Y _20138_/X _20092_/X _20138_/X VGND VGND VPWR VPWR _20141_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_117_0_HCLK clkbuf_7_58_0_HCLK/X VGND VGND VPWR VPWR _24872_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18246__B1 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20072_ _20067_/A VGND VGND VPWR VPWR _20072_/X sky130_fd_sc_hd__buf_2
XANTENNA__23119__A _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23900_ _23884_/CLK _18971_/X VGND VGND VPWR VPWR _18970_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_218_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24880_ _24834_/CLK _24880_/D HRESETn VGND VGND VPWR VPWR _24880_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18261__A3 _16267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23831_ _23831_/CLK _23831_/D VGND VGND VPWR VPWR _23831_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21862__A _24584_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23762_ _24089_/CLK _23762_/D VGND VGND VPWR VPWR _17949_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20974_ _12119_/B _12147_/A VGND VGND VPWR VPWR _20974_/X sky130_fd_sc_hd__and2_4
XFILLER_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25501_ _24209_/CLK _25501_/D HRESETn VGND VGND VPWR VPWR _11945_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22713_ _22713_/A _21235_/A VGND VGND VPWR VPWR _22713_/X sky130_fd_sc_hd__or2_4
XFILLER_241_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23693_ _23427_/CLK _19563_/X VGND VGND VPWR VPWR _19561_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_14_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24036__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13380__A _13254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25432_ _25428_/CLK _25432_/D HRESETn VGND VGND VPWR VPWR _12613_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22644_ _21055_/X _22639_/X _21832_/X _22643_/Y VGND VGND VPWR VPWR _22645_/A sky130_fd_sc_hd__a211o_4
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25363_ _25346_/CLK _13007_/Y HRESETn VGND VGND VPWR VPWR _25363_/Q sky130_fd_sc_hd__dfrtp_4
X_22575_ _22557_/Y _22563_/Y _22571_/Y _21445_/X _22574_/X VGND VGND VPWR VPWR _22575_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_166_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24314_ _24315_/CLK _24314_/D HRESETn VGND VGND VPWR VPWR _17563_/A sky130_fd_sc_hd__dfrtp_4
X_21526_ _21423_/A VGND VGND VPWR VPWR _22716_/A sky130_fd_sc_hd__buf_2
XFILLER_167_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25294_ _25091_/CLK _13691_/X HRESETn VGND VGND VPWR VPWR _11843_/A sky130_fd_sc_hd__dfrtp_4
X_24245_ _23767_/CLK _18134_/X HRESETn VGND VGND VPWR VPWR _24245_/Q sky130_fd_sc_hd__dfrtp_4
X_21457_ _21654_/A _19496_/Y VGND VGND VPWR VPWR _21457_/X sky130_fd_sc_hd__or2_4
XFILLER_135_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12190_ _25441_/Q VGND VGND VPWR VPWR _12191_/A sky130_fd_sc_hd__inv_2
X_20408_ _19072_/C _13741_/D _19803_/X VGND VGND VPWR VPWR _20408_/X sky130_fd_sc_hd__or3_4
X_21388_ _14668_/X _19778_/Y VGND VGND VPWR VPWR _21388_/X sky130_fd_sc_hd__or2_4
X_24176_ _24667_/CLK _24176_/D HRESETn VGND VGND VPWR VPWR _24176_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15525__A2_N _15519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_13_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_26_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_190_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23127_ _23235_/A _23127_/B VGND VGND VPWR VPWR _23127_/Y sky130_fd_sc_hd__nor2_4
XFILLER_162_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20339_ _21798_/B _20334_/X _19613_/A _20334_/X VGND VGND VPWR VPWR _23413_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_76_0_HCLK clkbuf_7_77_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_76_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18237__B1 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23058_ _15574_/Y _22989_/B VGND VGND VPWR VPWR _23058_/X sky130_fd_sc_hd__and2_4
XANTENNA__23230__B1 _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24877__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14900_ _24441_/Q VGND VGND VPWR VPWR _14900_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22009_ _21924_/A VGND VGND VPWR VPWR _22014_/A sky130_fd_sc_hd__buf_2
X_15880_ _15850_/A VGND VGND VPWR VPWR _15880_/X sky130_fd_sc_hd__buf_2
XFILLER_103_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22868__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24806__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14831_ _14805_/X _14829_/X _25198_/Q _14830_/X VGND VGND VPWR VPWR _14831_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_56_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21772__A _22380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14274__A1 _23442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17550_ _17587_/A _24113_/Q _17587_/A _24113_/Q VGND VGND VPWR VPWR _17550_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15770__A _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14762_ _14765_/A _14758_/B _14762_/C VGND VGND VPWR VPWR _14762_/X sky130_fd_sc_hd__or3_4
XFILLER_57_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11974_ _11932_/B _11963_/X _11973_/Y VGND VGND VPWR VPWR _25496_/D sky130_fd_sc_hd__o21a_4
XANTENNA__21544__B1 _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16501_ _16521_/A VGND VGND VPWR VPWR _16501_/X sky130_fd_sc_hd__buf_2
XFILLER_204_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13713_ _13672_/B _13712_/Y _13708_/X _13700_/X _11803_/A VGND VGND VPWR VPWR _25285_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_44_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17481_ _17460_/A _17481_/B VGND VGND VPWR VPWR _17482_/A sky130_fd_sc_hd__and2_4
X_14693_ _25064_/Q VGND VGND VPWR VPWR _22213_/A sky130_fd_sc_hd__inv_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16432_ _16432_/A VGND VGND VPWR VPWR _16432_/Y sky130_fd_sc_hd__inv_2
X_19220_ _23814_/Q VGND VGND VPWR VPWR _19220_/Y sky130_fd_sc_hd__inv_2
X_13644_ _13644_/A _13644_/B VGND VGND VPWR VPWR _13644_/X sky130_fd_sc_hd__or2_4
XFILLER_71_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19151_ _23839_/Q VGND VGND VPWR VPWR _19151_/Y sky130_fd_sc_hd__inv_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16363_ _16363_/A VGND VGND VPWR VPWR _16363_/Y sky130_fd_sc_hd__inv_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _13575_/A _13575_/B _13575_/C _13574_/X VGND VGND VPWR VPWR _14764_/A sky130_fd_sc_hd__or4_4
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18102_ _17966_/X _18101_/X _24246_/Q _18024_/X VGND VGND VPWR VPWR _18102_/X sky130_fd_sc_hd__o22a_4
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ _15314_/A VGND VGND VPWR VPWR _15314_/Y sky130_fd_sc_hd__inv_2
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12526_ _12526_/A VGND VGND VPWR VPWR _12644_/A sky130_fd_sc_hd__inv_2
X_19082_ _21894_/B _19079_/X _16873_/X _19079_/X VGND VGND VPWR VPWR _19082_/X sky130_fd_sc_hd__a2bb2o_4
X_16294_ _24637_/Q VGND VGND VPWR VPWR _16294_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18033_ _17979_/X _18033_/B VGND VGND VPWR VPWR _18033_/X sky130_fd_sc_hd__or2_4
X_15245_ _15245_/A _15265_/A _15261_/A _15261_/B VGND VGND VPWR VPWR _15254_/B sky130_fd_sc_hd__or4_4
XFILLER_185_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12457_ _12270_/D _12456_/X VGND VGND VPWR VPWR _12458_/B sky130_fd_sc_hd__or2_4
XANTENNA__15648__C _16446_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15176_ _15165_/A _15174_/X _15176_/C VGND VGND VPWR VPWR _15176_/X sky130_fd_sc_hd__and3_4
XFILLER_114_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12388_ _12204_/Y _12385_/X VGND VGND VPWR VPWR _12388_/X sky130_fd_sc_hd__or2_4
XFILLER_141_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14127_ _14114_/X _14126_/Y _14092_/A _14114_/X VGND VGND VPWR VPWR _14127_/X sky130_fd_sc_hd__a2bb2o_4
X_19984_ _19984_/A VGND VGND VPWR VPWR _19984_/X sky130_fd_sc_hd__buf_2
XFILLER_113_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14058_ _14067_/A VGND VGND VPWR VPWR _14058_/X sky130_fd_sc_hd__buf_2
X_18935_ _18931_/Y _18934_/X _17415_/X _18934_/X VGND VGND VPWR VPWR _23914_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13009_ _13008_/X VGND VGND VPWR VPWR _13009_/Y sky130_fd_sc_hd__inv_2
X_18866_ _18862_/X _18866_/B _18864_/X _18865_/X VGND VGND VPWR VPWR _18867_/D sky130_fd_sc_hd__or4_4
XFILLER_94_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21783__B1 _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24547__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21682__A _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17817_ _17817_/A _17817_/B VGND VGND VPWR VPWR _17818_/C sky130_fd_sc_hd__or2_4
X_18797_ _18797_/A _18797_/B VGND VGND VPWR VPWR _18798_/A sky130_fd_sc_hd__or2_4
X_17748_ _24262_/Q VGND VGND VPWR VPWR _17748_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21535__B1 _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17679_ _17670_/A _17670_/B VGND VGND VPWR VPWR _17680_/C sky130_fd_sc_hd__nand2_4
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19418_ _18037_/B VGND VGND VPWR VPWR _19418_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20690_ _20780_/A VGND VGND VPWR VPWR _20690_/X sky130_fd_sc_hd__buf_2
XANTENNA__23288__B1 _24288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21838__A1 _20517_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22944__C _22817_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19349_ _19347_/Y _19343_/X _19282_/X _19348_/X VGND VGND VPWR VPWR _19349_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22360_ _21935_/A _19876_/Y _21207_/A VGND VGND VPWR VPWR _22360_/X sky130_fd_sc_hd__o21a_4
XFILLER_248_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25335__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16714__B1 _16358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21311_ _21297_/Y VGND VGND VPWR VPWR _21311_/X sky130_fd_sc_hd__buf_2
XFILLER_164_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22291_ _22291_/A _22417_/B VGND VGND VPWR VPWR _22291_/X sky130_fd_sc_hd__and2_4
XFILLER_248_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16016__A _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21242_ _22196_/A VGND VGND VPWR VPWR _21627_/A sky130_fd_sc_hd__buf_2
X_24030_ _24060_/CLK _20808_/Y HRESETn VGND VGND VPWR VPWR _24030_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21173_ _21323_/A _21170_/X _21172_/X VGND VGND VPWR VPWR _21173_/X sky130_fd_sc_hd__and3_4
XFILLER_144_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20124_ _20123_/Y _20121_/X _20099_/X _20121_/X VGND VGND VPWR VPWR _23495_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24970__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20055_ _20055_/A VGND VGND VPWR VPWR _20055_/X sky130_fd_sc_hd__buf_2
X_24932_ _25070_/CLK _15525_/X HRESETn VGND VGND VPWR VPWR _21133_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24288__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21774__B1 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24863_ _25409_/CLK _24863_/D HRESETn VGND VGND VPWR VPWR _24863_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24217__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22318__A2 _21349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23814_ _23873_/CLK _19222_/X VGND VGND VPWR VPWR _23814_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24794_ _24795_/CLK _15891_/X HRESETn VGND VGND VPWR VPWR _22482_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _23785_/CLK _23745_/D VGND VGND VPWR VPWR _19416_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_226_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _20953_/X VGND VGND VPWR VPWR _20957_/Y sky130_fd_sc_hd__inv_2
XPHY_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23279__B1 _24885_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11690_/A VGND VGND VPWR VPWR _11690_/Y sky130_fd_sc_hd__inv_2
X_23676_ _24317_/CLK _23676_/D VGND VGND VPWR VPWR _19619_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_214_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _20888_/A VGND VGND VPWR VPWR _20888_/Y sky130_fd_sc_hd__inv_2
XPHY_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25415_ _25403_/CLK _12679_/Y HRESETn VGND VGND VPWR VPWR _25415_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22627_ _24559_/Q _22432_/X _22536_/X VGND VGND VPWR VPWR _22627_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23312__A _22716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17310__A _17249_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13360_ _13200_/A _13360_/B VGND VGND VPWR VPWR _13360_/X sky130_fd_sc_hd__or2_4
X_25346_ _25346_/CLK _25346_/D HRESETn VGND VGND VPWR VPWR _12280_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25076__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22558_ _22558_/A _21441_/X VGND VGND VPWR VPWR _22558_/X sky130_fd_sc_hd__or2_4
XFILLER_220_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16705__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12311_ _25342_/Q VGND VGND VPWR VPWR _13072_/A sky130_fd_sc_hd__inv_2
X_21509_ _21178_/X VGND VGND VPWR VPWR _21510_/A sky130_fd_sc_hd__buf_2
XFILLER_127_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25005__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13291_ _13200_/A _23455_/Q VGND VGND VPWR VPWR _13291_/X sky130_fd_sc_hd__or2_4
X_25277_ _23528_/CLK _13756_/X HRESETn VGND VGND VPWR VPWR _13736_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22489_ _21311_/X VGND VGND VPWR VPWR _22489_/X sky130_fd_sc_hd__buf_2
XFILLER_10_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15030_ _14921_/X _24465_/Q _14921_/X _24465_/Q VGND VGND VPWR VPWR _15035_/B sky130_fd_sc_hd__a2bb2o_4
X_12242_ _25437_/Q VGND VGND VPWR VPWR _12266_/C sky130_fd_sc_hd__inv_2
X_24228_ _24233_/CLK _18259_/X HRESETn VGND VGND VPWR VPWR _11841_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21767__A _22381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12742__B2 _24801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12173_ _12172_/Y _23101_/A _12172_/Y _23101_/A VGND VGND VPWR VPWR _12173_/X sky130_fd_sc_hd__a2bb2o_4
X_24159_ _24159_/CLK _24159_/D HRESETn VGND VGND VPWR VPWR _18595_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16981_ _24725_/Q _24382_/Q _16049_/Y _17035_/A VGND VGND VPWR VPWR _16981_/X sky130_fd_sc_hd__o22a_4
XFILLER_123_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19958__B1 _19874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18720_ _18719_/X VGND VGND VPWR VPWR _18720_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13285__A _13285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_100_0_HCLK clkbuf_7_50_0_HCLK/X VGND VGND VPWR VPWR _25521_/CLK sky130_fd_sc_hd__clkbuf_1
X_15932_ _15931_/X VGND VGND VPWR VPWR _15932_/X sky130_fd_sc_hd__buf_2
XFILLER_237_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24640__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_163_0_HCLK clkbuf_7_81_0_HCLK/X VGND VGND VPWR VPWR _23890_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_49_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_6_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15863_ _12770_/Y _15862_/X _15557_/X _15862_/X VGND VGND VPWR VPWR _24814_/D sky130_fd_sc_hd__a2bb2o_4
X_18651_ _16576_/Y _24143_/Q _16566_/A _18613_/X VGND VGND VPWR VPWR _18651_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_236_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14814_ _14814_/A _14814_/B _14814_/C VGND VGND VPWR VPWR _14815_/B sky130_fd_sc_hd__and3_4
X_17602_ _17614_/A _17602_/B VGND VGND VPWR VPWR _17602_/X sky130_fd_sc_hd__and2_4
XANTENNA__12258__B1 _12252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15794_ _12316_/Y _15793_/X _15557_/X _15793_/X VGND VGND VPWR VPWR _24849_/D sky130_fd_sc_hd__a2bb2o_4
X_18582_ _18563_/B VGND VGND VPWR VPWR _18583_/B sky130_fd_sc_hd__inv_2
X_14745_ _14671_/X _14739_/X VGND VGND VPWR VPWR _14745_/X sky130_fd_sc_hd__and2_4
X_17533_ _11732_/Y _17568_/A _11732_/Y _17568_/A VGND VGND VPWR VPWR _17533_/X sky130_fd_sc_hd__a2bb2o_4
X_11957_ _24324_/Q VGND VGND VPWR VPWR _17479_/C sky130_fd_sc_hd__inv_2
XFILLER_33_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17464_ _20220_/A VGND VGND VPWR VPWR _18910_/A sky130_fd_sc_hd__inv_2
X_14676_ _25061_/Q VGND VGND VPWR VPWR _22056_/A sky130_fd_sc_hd__buf_2
XFILLER_233_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11888_ _11848_/B _11883_/Y VGND VGND VPWR VPWR _11888_/X sky130_fd_sc_hd__and2_4
XFILLER_149_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20846__A _20846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16415_ _16415_/A VGND VGND VPWR VPWR _16415_/Y sky130_fd_sc_hd__inv_2
X_19203_ _19360_/A VGND VGND VPWR VPWR _19203_/X sky130_fd_sc_hd__buf_2
X_13627_ _13512_/Y VGND VGND VPWR VPWR _13627_/X sky130_fd_sc_hd__buf_2
XANTENNA__16963__A1_N _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17395_ _23986_/Q _17394_/X VGND VGND VPWR VPWR _17396_/B sky130_fd_sc_hd__or2_4
XANTENNA__23285__A3 _22135_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16346_ _24617_/Q VGND VGND VPWR VPWR _16346_/Y sky130_fd_sc_hd__inv_2
X_19134_ _19132_/Y _19133_/X _19063_/X _19133_/X VGND VGND VPWR VPWR _19134_/X sky130_fd_sc_hd__a2bb2o_4
X_13558_ _13556_/A _14563_/C _13556_/Y _14570_/A VGND VGND VPWR VPWR _13565_/B sky130_fd_sc_hd__o22a_4
XFILLER_158_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12509_ _12509_/A VGND VGND VPWR VPWR _12664_/C sky130_fd_sc_hd__buf_2
X_19065_ _23868_/Q VGND VGND VPWR VPWR _19065_/Y sky130_fd_sc_hd__inv_2
X_16277_ _16277_/A VGND VGND VPWR VPWR _16318_/A sky130_fd_sc_hd__buf_2
X_13489_ _11976_/Y _13485_/X _11761_/X _13488_/X VGND VGND VPWR VPWR _25314_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15228_ _15228_/A _15228_/B VGND VGND VPWR VPWR _15230_/B sky130_fd_sc_hd__or2_4
X_18016_ _18016_/A _23833_/Q VGND VGND VPWR VPWR _18016_/X sky130_fd_sc_hd__or2_4
XANTENNA__15380__C1 _15334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24799__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15159_ _15242_/B VGND VGND VPWR VPWR _15311_/B sky130_fd_sc_hd__buf_2
XANTENNA__24728__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19967_ _19967_/A VGND VGND VPWR VPWR _19967_/X sky130_fd_sc_hd__buf_2
XFILLER_102_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18918_ _18925_/A VGND VGND VPWR VPWR _18918_/X sky130_fd_sc_hd__buf_2
X_19898_ _13745_/A _13737_/X _20136_/A _19898_/D VGND VGND VPWR VPWR _19898_/X sky130_fd_sc_hd__or4_4
XANTENNA__24381__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18849_ _16527_/A _18787_/A _16520_/A _18788_/B VGND VGND VPWR VPWR _18849_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21843__C _21741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24310__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12249__B1 _12248_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21860_ _16719_/A VGND VGND VPWR VPWR _23091_/A sky130_fd_sc_hd__buf_2
XFILLER_215_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20811_ _13125_/B _20805_/A _20810_/X VGND VGND VPWR VPWR _20811_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_24_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21791_ _21654_/A _21791_/B VGND VGND VPWR VPWR _21791_/X sky130_fd_sc_hd__or2_4
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22720__A2 _22718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23530_ _24199_/CLK _20035_/X VGND VGND VPWR VPWR _20031_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__19610__A _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20742_ _13120_/A _13120_/B _20741_/Y VGND VGND VPWR VPWR _20742_/Y sky130_fd_sc_hd__a21oi_4
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25516__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16935__B1 _22564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23461_ _24252_/CLK _20214_/X VGND VGND VPWR VPWR _18139_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_51_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20673_ _20673_/A _14271_/X VGND VGND VPWR VPWR _20675_/B sky130_fd_sc_hd__or2_4
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25200_ _25056_/CLK _14216_/X HRESETn VGND VGND VPWR VPWR _14215_/A sky130_fd_sc_hd__dfstp_4
XFILLER_195_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22412_ _24619_/Q _22275_/X VGND VGND VPWR VPWR _22412_/X sky130_fd_sc_hd__or2_4
XFILLER_149_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23392_ _23391_/CLK _23392_/D VGND VGND VPWR VPWR _20386_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_137_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22971__A _22451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25131_ _25117_/CLK _14439_/X HRESETn VGND VGND VPWR VPWR _25131_/Q sky130_fd_sc_hd__dfstp_4
X_22343_ _22343_/A _22343_/B VGND VGND VPWR VPWR _22345_/B sky130_fd_sc_hd__or2_4
XFILLER_128_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17360__B1 _17284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25062_ _23494_/CLK _25062_/D HRESETn VGND VGND VPWR VPWR _21252_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21587__A _21587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22274_ _21581_/X VGND VGND VPWR VPWR _22274_/X sky130_fd_sc_hd__buf_2
XFILLER_88_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24013_ _24049_/CLK _20737_/X HRESETn VGND VGND VPWR VPWR _13118_/A sky130_fd_sc_hd__dfrtp_4
X_21225_ _24035_/Q VGND VGND VPWR VPWR _21225_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24469__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21156_ _23965_/Q VGND VGND VPWR VPWR _21156_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20107_ _21618_/B _20105_/X _20106_/X _20105_/X VGND VGND VPWR VPWR _23501_/D sky130_fd_sc_hd__a2bb2o_4
X_21087_ _21087_/A VGND VGND VPWR VPWR _22420_/B sky130_fd_sc_hd__buf_2
XANTENNA__12488__B1 _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20038_ _20038_/A VGND VGND VPWR VPWR _20038_/Y sky130_fd_sc_hd__inv_2
X_24915_ _24508_/CLK _15579_/X HRESETn VGND VGND VPWR VPWR _15578_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_236_0_HCLK clkbuf_8_237_0_HCLK/A VGND VGND VPWR VPWR _25043_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24051__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12860_ _12769_/Y _12860_/B VGND VGND VPWR VPWR _12860_/X sky130_fd_sc_hd__or2_4
X_24846_ _25390_/CLK _24846_/D HRESETn VGND VGND VPWR VPWR _24846_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11811_/A VGND VGND VPWR VPWR _22735_/A sky130_fd_sc_hd__inv_2
XFILLER_215_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12912_/A _22714_/A _12912_/A _22714_/A VGND VGND VPWR VPWR _12792_/D sky130_fd_sc_hd__a2bb2o_4
X_24777_ _25380_/CLK _15933_/X HRESETn VGND VGND VPWR VPWR _12205_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_199_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ _21989_/A VGND VGND VPWR VPWR _21990_/D sky130_fd_sc_hd__inv_2
XFILLER_233_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14530_/A _14530_/B VGND VGND VPWR VPWR _25101_/D sky130_fd_sc_hd__or2_4
XFILLER_215_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22711__A2 _22416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ HWDATA[12] VGND VGND VPWR VPWR _16236_/A sky130_fd_sc_hd__buf_2
X_23728_ _23437_/CLK _19464_/X VGND VGND VPWR VPWR _19462_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12660__B1 _12627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16926__B1 _22153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _25121_/Q VGND VGND VPWR VPWR _14461_/Y sky130_fd_sc_hd__inv_2
XFILLER_230_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A _11673_/B _11671_/X _11672_/X VGND VGND VPWR VPWR _15640_/C sky130_fd_sc_hd__or4_4
X_23659_ _24209_/CLK _19669_/X VGND VGND VPWR VPWR _13435_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _23132_/A VGND VGND VPWR VPWR _16200_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23267__A3 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13254_/A _13410_/X _13412_/C VGND VGND VPWR VPWR _13412_/X sky130_fd_sc_hd__and3_4
X_17180_ _24630_/Q _17179_/A _16313_/Y _17179_/Y VGND VGND VPWR VPWR _17180_/X sky130_fd_sc_hd__o22a_4
XFILLER_169_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ _14392_/A VGND VGND VPWR VPWR _14392_/X sky130_fd_sc_hd__buf_2
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16131_ _22662_/A VGND VGND VPWR VPWR _16131_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13343_ _13234_/X _13343_/B VGND VGND VPWR VPWR _13343_/X sky130_fd_sc_hd__or2_4
X_25329_ _23456_/CLK _13355_/X HRESETn VGND VGND VPWR VPWR _25329_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12184__A _21078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16062_ _14407_/A VGND VGND VPWR VPWR _16062_/X sky130_fd_sc_hd__buf_2
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13274_ _13199_/A VGND VGND VPWR VPWR _13312_/A sky130_fd_sc_hd__buf_2
XFILLER_155_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24892__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15013_ _25038_/Q _24476_/Q _14972_/Y _15012_/Y VGND VGND VPWR VPWR _15016_/C sky130_fd_sc_hd__o22a_4
X_12225_ _25447_/Q VGND VGND VPWR VPWR _12273_/B sky130_fd_sc_hd__inv_2
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12912__A _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24821__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19821_ _21752_/B _19814_/X _19820_/X _19814_/X VGND VGND VPWR VPWR _23606_/D sky130_fd_sc_hd__a2bb2o_4
X_12156_ _12155_/X VGND VGND VPWR VPWR _12156_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24139__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_46_0_HCLK clkbuf_6_46_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_93_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19752_ _19751_/Y _19747_/X _19728_/X _19747_/X VGND VGND VPWR VPWR _19752_/X sky130_fd_sc_hd__a2bb2o_4
X_12087_ _16181_/A _12087_/B VGND VGND VPWR VPWR _12087_/X sky130_fd_sc_hd__or2_4
X_16964_ _16964_/A VGND VGND VPWR VPWR _17032_/A sky130_fd_sc_hd__inv_2
XFILLER_238_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18703_ _18703_/A _18703_/B VGND VGND VPWR VPWR _18704_/C sky130_fd_sc_hd__nand2_4
X_15915_ _15681_/X _15913_/Y _15673_/X _15913_/Y VGND VGND VPWR VPWR _24783_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19683_ _19682_/Y _19678_/X _19587_/X _19678_/X VGND VGND VPWR VPWR _19683_/X sky130_fd_sc_hd__a2bb2o_4
X_16895_ _16895_/A VGND VGND VPWR VPWR _16895_/X sky130_fd_sc_hd__buf_2
X_18634_ _24524_/Q _24135_/Q _16596_/Y _18789_/A VGND VGND VPWR VPWR _18634_/X sky130_fd_sc_hd__o22a_4
X_15846_ _21583_/A VGND VGND VPWR VPWR _21579_/B sky130_fd_sc_hd__buf_2
XFILLER_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18565_ _18577_/A _18577_/B VGND VGND VPWR VPWR _18566_/B sky130_fd_sc_hd__or2_4
X_12989_ _13000_/A _12285_/Y _12315_/Y _13000_/D VGND VGND VPWR VPWR _12989_/X sky130_fd_sc_hd__or4_4
X_15777_ _15724_/A VGND VGND VPWR VPWR _15777_/X sky130_fd_sc_hd__buf_2
XFILLER_240_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18906__B2 _11794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_HCLK clkbuf_3_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17516_ _17516_/A VGND VGND VPWR VPWR _17516_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14728_ _14727_/X VGND VGND VPWR VPWR _14728_/Y sky130_fd_sc_hd__inv_2
X_18496_ _18416_/Y _18496_/B VGND VGND VPWR VPWR _18497_/C sky130_fd_sc_hd__or2_4
XFILLER_220_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14659_ _13606_/B _13586_/A VGND VGND VPWR VPWR _20199_/B sky130_fd_sc_hd__or2_4
X_17447_ _21220_/A _21177_/A _17446_/X VGND VGND VPWR VPWR _17448_/A sky130_fd_sc_hd__or3_4
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18691__D _18658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17378_ _17351_/A _17374_/X _17377_/Y VGND VGND VPWR VPWR _24343_/D sky130_fd_sc_hd__and3_4
XFILLER_119_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19117_ _19117_/A _19163_/B _19320_/C VGND VGND VPWR VPWR _19117_/X sky130_fd_sc_hd__or3_4
X_16329_ _24624_/Q VGND VGND VPWR VPWR _16329_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24909__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19048_ _19047_/X VGND VGND VPWR VPWR _19054_/A sky130_fd_sc_hd__inv_2
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24562__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21010_ _24334_/Q _21010_/B VGND VGND VPWR VPWR _21010_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15656__B1 _20822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22669__C _22668_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22961_ _16113_/Y _22559_/X _15855_/B _11710_/Y _21051_/A VGND VGND VPWR VPWR _22961_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24700_ _24753_/CLK _24700_/D HRESETn VGND VGND VPWR VPWR _22909_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_216_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21912_ _22083_/A _20123_/Y VGND VGND VPWR VPWR _21914_/B sky130_fd_sc_hd__or2_4
XFILLER_83_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22892_ _24464_/Q _22431_/X _22891_/X VGND VGND VPWR VPWR _22892_/X sky130_fd_sc_hd__o21a_4
XFILLER_244_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24631_ _24623_/CLK _24631_/D HRESETn VGND VGND VPWR VPWR _24631_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_215_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21843_ _16527_/A _21843_/B _21741_/B VGND VGND VPWR VPWR _21843_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_66_0_HCLK clkbuf_8_67_0_HCLK/A VGND VGND VPWR VPWR _24266_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22154__B1 _25525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17492__A2_N _24114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24562_ _24540_/CLK _16499_/X HRESETn VGND VGND VPWR VPWR _24562_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25350__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21774_ _21769_/X _21772_/X _21773_/X VGND VGND VPWR VPWR _21774_/X sky130_fd_sc_hd__o21a_4
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12642__B1 _12641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23513_ _24199_/CLK _23513_/D VGND VGND VPWR VPWR _23513_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20725_ _15612_/Y _20708_/X _20716_/X _20724_/Y VGND VGND VPWR VPWR _20725_/X sky130_fd_sc_hd__o22a_4
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24493_ _24049_/CLK _16683_/X HRESETn VGND VGND VPWR VPWR _16682_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11901__A _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23444_ _23859_/CLK _23444_/D VGND VGND VPWR VPWR _20257_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20656_ _17393_/A _17393_/B VGND VGND VPWR VPWR _20657_/B sky130_fd_sc_hd__nand2_4
XFILLER_7_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17795__A _16940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23375_ _24907_/CLK _20822_/A VGND VGND VPWR VPWR _23375_/Q sky130_fd_sc_hd__dfxtp_4
X_20587_ _20586_/X VGND VGND VPWR VPWR _23946_/D sky130_fd_sc_hd__inv_2
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25114_ _25109_/CLK _25114_/D HRESETn VGND VGND VPWR VPWR _25114_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22326_ _22325_/X VGND VGND VPWR VPWR _22326_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15895__B1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21417__C1 _21416_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25045_ _25056_/CLK _25045_/D HRESETn VGND VGND VPWR VPWR _14808_/C sky130_fd_sc_hd__dfrtp_4
X_22257_ _22257_/A _22253_/X _22257_/C VGND VGND VPWR VPWR _22257_/X sky130_fd_sc_hd__or3_4
XANTENNA__12732__A _25399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12010_ _24097_/Q _12002_/A _12007_/Y VGND VGND VPWR VPWR _12010_/X sky130_fd_sc_hd__o21a_4
X_21208_ _21208_/A _21208_/B VGND VGND VPWR VPWR _21210_/B sky130_fd_sc_hd__or2_4
XFILLER_2_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18833__B1 _16530_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22188_ _21345_/Y _22174_/X _22176_/X _22180_/Y _22187_/X VGND VGND VPWR VPWR _22195_/C
+ sky130_fd_sc_hd__a2111o_4
XFILLER_133_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24232__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21139_ _14419_/Y _14209_/A _21137_/Y _21348_/A VGND VGND VPWR VPWR _21139_/X sky130_fd_sc_hd__o22a_4
XFILLER_132_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13961_ scl_oen_o_S5 _13955_/X _13956_/Y _13960_/Y VGND VGND VPWR VPWR _13961_/X
+ sky130_fd_sc_hd__o22a_4
XANTENNA__23037__A _21080_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12912_ _12912_/A _12890_/X VGND VGND VPWR VPWR _12912_/X sky130_fd_sc_hd__or2_4
X_15700_ _15699_/Y VGND VGND VPWR VPWR _15700_/X sky130_fd_sc_hd__buf_2
XFILLER_246_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16680_ _16668_/A VGND VGND VPWR VPWR _16680_/X sky130_fd_sc_hd__buf_2
XFILLER_234_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13892_ _13892_/A VGND VGND VPWR VPWR _13935_/A sky130_fd_sc_hd__buf_2
XANTENNA__12881__B1 _12862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16072__B1 _15901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12843_ _12735_/Y _12842_/X VGND VGND VPWR VPWR _12851_/A sky130_fd_sc_hd__or2_4
X_15631_ _21593_/A _15628_/X _15472_/X _15628_/X VGND VGND VPWR VPWR _24895_/D sky130_fd_sc_hd__a2bb2o_4
X_24829_ _25428_/CLK _15822_/X HRESETn VGND VGND VPWR VPWR _24829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14622__A1 _14610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14622__B2 _14611_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15562_ _15559_/Y _15553_/X _15560_/X _15561_/X VGND VGND VPWR VPWR _15562_/X sky130_fd_sc_hd__a2bb2o_4
X_18350_ _18350_/A VGND VGND VPWR VPWR _18350_/Y sky130_fd_sc_hd__inv_2
X_12774_ _12772_/A _22482_/A _12834_/A _12773_/Y VGND VGND VPWR VPWR _12778_/C sky130_fd_sc_hd__o22a_4
XANTENNA__25091__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _21847_/A _14500_/X _25105_/Q _14502_/X VGND VGND VPWR VPWR _14513_/X sky130_fd_sc_hd__o22a_4
X_17301_ _17284_/A _17301_/B _17300_/X VGND VGND VPWR VPWR _17301_/X sky130_fd_sc_hd__or3_4
XFILLER_242_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _25536_/Q VGND VGND VPWR VPWR _11725_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25020__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _11670_/A VGND VGND VPWR VPWR _15493_/Y sky130_fd_sc_hd__inv_2
X_18281_ _18279_/A VGND VGND VPWR VPWR _18282_/A sky130_fd_sc_hd__inv_2
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _20600_/A _14443_/X _14400_/X _14443_/X VGND VGND VPWR VPWR _25129_/D sky130_fd_sc_hd__a2bb2o_4
X_17232_ _24371_/Q VGND VGND VPWR VPWR _17232_/Y sky130_fd_sc_hd__inv_2
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _13453_/A VGND VGND VPWR VPWR _15636_/B sky130_fd_sc_hd__inv_2
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17163_ _16331_/Y _24352_/Q _16331_/Y _24352_/Q VGND VGND VPWR VPWR _17169_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14375_ _25152_/Q VGND VGND VPWR VPWR _14375_/Y sky130_fd_sc_hd__inv_2
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17324__B1 _17276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16114_ _16113_/Y _16111_/X _15946_/X _16111_/X VGND VGND VPWR VPWR _24701_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13326_ _13390_/A _13326_/B _13326_/C VGND VGND VPWR VPWR _13330_/B sky130_fd_sc_hd__and3_4
X_17094_ _17105_/A _17092_/X _17093_/X VGND VGND VPWR VPWR _24394_/D sky130_fd_sc_hd__and3_4
XFILLER_155_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15886__B1 _24797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16045_ _16038_/A VGND VGND VPWR VPWR _16045_/X sky130_fd_sc_hd__buf_2
XANTENNA__21020__A _21019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13257_ _13392_/A _18938_/A VGND VGND VPWR VPWR _13257_/X sky130_fd_sc_hd__or2_4
XFILLER_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12353__A2_N _24824_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12208_ _12208_/A VGND VGND VPWR VPWR _12208_/X sky130_fd_sc_hd__buf_2
X_13188_ _13247_/A VGND VGND VPWR VPWR _13193_/A sky130_fd_sc_hd__buf_2
XFILLER_97_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19804_ _19072_/C _19898_/D _19803_/X VGND VGND VPWR VPWR _19805_/A sky130_fd_sc_hd__or3_4
XFILLER_123_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12139_ _12139_/A _12135_/X VGND VGND VPWR VPWR _12141_/A sky130_fd_sc_hd__and2_4
XANTENNA__15953__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17996_ _18227_/A _17989_/X _17996_/C VGND VGND VPWR VPWR _17996_/X sky130_fd_sc_hd__or3_4
X_19735_ _13443_/B VGND VGND VPWR VPWR _19735_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16947_ _16149_/Y _22190_/A _16157_/Y _24261_/Q VGND VGND VPWR VPWR _16947_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22384__B1 _14666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19666_ _19666_/A VGND VGND VPWR VPWR _19666_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16878_ _19820_/A VGND VGND VPWR VPWR _16878_/X sky130_fd_sc_hd__buf_2
XFILLER_226_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16063__B1 _16062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22786__A _22468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18617_ _16619_/Y _18616_/X _16619_/Y _18616_/X VGND VGND VPWR VPWR _18618_/D sky130_fd_sc_hd__a2bb2o_4
X_15829_ _15813_/A VGND VGND VPWR VPWR _15829_/X sky130_fd_sc_hd__buf_2
XFILLER_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25108__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19597_ _19597_/A _19939_/B _18284_/X VGND VGND VPWR VPWR _19598_/A sky130_fd_sc_hd__or3_4
XFILLER_241_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18548_ _18523_/X _18538_/B _18547_/X VGND VGND VPWR VPWR _24173_/D sky130_fd_sc_hd__and3_4
XANTENNA__22687__A1 _16272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20698__B1 _20696_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18479_ _18556_/A _18479_/B _18478_/X VGND VGND VPWR VPWR _18479_/X sky130_fd_sc_hd__or3_4
X_20510_ _20510_/A _20510_/B VGND VGND VPWR VPWR _20510_/X sky130_fd_sc_hd__and2_4
XANTENNA__11721__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21490_ _21483_/X _21488_/X _21489_/X VGND VGND VPWR VPWR _21490_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22439__B2 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20441_ _14485_/X VGND VGND VPWR VPWR _20441_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17315__B1 _17268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24743__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23160_ _23160_/A _23147_/X _23160_/C _23159_/X VGND VGND VPWR VPWR _23160_/X sky130_fd_sc_hd__or4_4
XFILLER_119_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20372_ _18240_/A VGND VGND VPWR VPWR _20372_/X sky130_fd_sc_hd__buf_2
XFILLER_174_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15877__B1 _11718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22111_ _22111_/A VGND VGND VPWR VPWR _22111_/X sky130_fd_sc_hd__buf_2
XANTENNA__19068__B1 _19067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23091_ _23091_/A _23091_/B _23090_/X VGND VGND VPWR VPWR _23091_/X sky130_fd_sc_hd__and3_4
XANTENNA__16024__A _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22042_ _22043_/A _19592_/Y VGND VGND VPWR VPWR _22042_/X sky130_fd_sc_hd__and2_4
XANTENNA__22611__A1 _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15629__B1 _15469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20622__B1 _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21584__B _21741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23993_ _24340_/CLK _23993_/D HRESETn VGND VGND VPWR VPWR _23993_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_217_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14479__A _18951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22944_ _22944_/A _22821_/B _22817_/C VGND VGND VPWR VPWR _22944_/X sky130_fd_sc_hd__and3_4
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12863__B1 _12862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25531__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22875_ _17179_/Y _22430_/X _25386_/Q _22299_/X VGND VGND VPWR VPWR _22875_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22127__B1 _22095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24614_ _24346_/CLK _16356_/X HRESETn VGND VGND VPWR VPWR _24614_/Q sky130_fd_sc_hd__dfrtp_4
X_21826_ _13772_/D _21826_/B VGND VGND VPWR VPWR _21827_/C sky130_fd_sc_hd__or2_4
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24545_ _24080_/CLK _16545_/X HRESETn VGND VGND VPWR VPWR _24545_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21757_ _21757_/A _21755_/X _21756_/X VGND VGND VPWR VPWR _21757_/X sky130_fd_sc_hd__and3_4
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20708_ _20708_/A VGND VGND VPWR VPWR _20708_/X sky130_fd_sc_hd__buf_2
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _12211_/Y _12493_/B VGND VGND VPWR VPWR _12490_/Y sky130_fd_sc_hd__nand2_4
X_24476_ _25015_/CLK _24476_/D HRESETn VGND VGND VPWR VPWR _24476_/Q sky130_fd_sc_hd__dfrtp_4
X_21688_ _21954_/A _21679_/X _21687_/X VGND VGND VPWR VPWR _21688_/X sky130_fd_sc_hd__or3_4
XFILLER_211_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23427_ _23427_/CLK _20303_/X VGND VGND VPWR VPWR _20302_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23320__A _23320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20639_ _23980_/Q _17389_/B VGND VGND VPWR VPWR _20639_/Y sky130_fd_sc_hd__nand2_4
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24484__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14160_ _14160_/A _23956_/Q VGND VGND VPWR VPWR _14161_/A sky130_fd_sc_hd__or2_4
X_23358_ VGND VGND VPWR VPWR _23358_/HI sda_o_S4 sky130_fd_sc_hd__conb_1
XANTENNA__22850__B2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24413__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13111_ _13111_/A _13111_/B VGND VGND VPWR VPWR _13112_/A sky130_fd_sc_hd__and2_4
X_22309_ _24587_/Q _22701_/B VGND VGND VPWR VPWR _22309_/X sky130_fd_sc_hd__or2_4
X_14091_ _14091_/A _14091_/B _14106_/A VGND VGND VPWR VPWR _14092_/B sky130_fd_sc_hd__or3_4
XFILLER_4_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23289_ _17232_/Y _22485_/X _12818_/A _22444_/X VGND VGND VPWR VPWR _23289_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_111_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_222_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13042_ _12324_/Y _13046_/A _12291_/X _13051_/B VGND VGND VPWR VPWR _13048_/B sky130_fd_sc_hd__or4_4
X_25028_ _25028_/CLK _15213_/Y HRESETn VGND VGND VPWR VPWR _25028_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17850_ _17750_/D _17555_/X VGND VGND VPWR VPWR _17850_/X sky130_fd_sc_hd__or2_4
XFILLER_79_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16293__B1 _15567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16801_ _14962_/Y _16799_/X _16464_/X _16799_/X VGND VGND VPWR VPWR _24442_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17781_ _16913_/Y _17779_/A VGND VGND VPWR VPWR _17782_/C sky130_fd_sc_hd__or2_4
X_14993_ _14903_/X _24446_/Q _14903_/X _24446_/Q VGND VGND VPWR VPWR _14997_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19520_ _21190_/B _19515_/X _19475_/X _19502_/Y VGND VGND VPWR VPWR _23707_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16732_ _24474_/Q VGND VGND VPWR VPWR _16732_/Y sky130_fd_sc_hd__inv_2
X_13944_ _13944_/A _13923_/D _15421_/B VGND VGND VPWR VPWR _13949_/A sky130_fd_sc_hd__or3_4
XANTENNA__25272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19451_ _18209_/B VGND VGND VPWR VPWR _19451_/Y sky130_fd_sc_hd__inv_2
X_13875_ _23993_/Q VGND VGND VPWR VPWR _13956_/A sky130_fd_sc_hd__buf_2
X_16663_ _24501_/Q VGND VGND VPWR VPWR _16663_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22118__B1 _22117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18402_ _18528_/A VGND VGND VPWR VPWR _18468_/A sky130_fd_sc_hd__inv_2
XFILLER_234_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12826_ _12825_/X VGND VGND VPWR VPWR _12967_/A sky130_fd_sc_hd__buf_2
X_15614_ _15612_/Y _15608_/X _11757_/X _15613_/X VGND VGND VPWR VPWR _15614_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19382_ _18168_/B VGND VGND VPWR VPWR _19382_/Y sky130_fd_sc_hd__inv_2
X_16594_ _24525_/Q VGND VGND VPWR VPWR _16594_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18333_ _17460_/A VGND VGND VPWR VPWR _19094_/B sky130_fd_sc_hd__buf_2
X_12757_ _24793_/Q VGND VGND VPWR VPWR _12757_/Y sky130_fd_sc_hd__inv_2
X_15545_ HWDATA[31] VGND VGND VPWR VPWR _15545_/X sky130_fd_sc_hd__buf_2
XFILLER_42_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21341__A1 _24516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11681_/X VGND VGND VPWR VPWR _11708_/X sky130_fd_sc_hd__buf_2
XFILLER_202_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15476_ _14876_/Y _15471_/X _15475_/X _15458_/A VGND VGND VPWR VPWR _15476_/X sky130_fd_sc_hd__a2bb2o_4
X_18264_ _18263_/X _20369_/A VGND VGND VPWR VPWR _18264_/X sky130_fd_sc_hd__or2_4
XFILLER_188_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12688_ _12687_/X VGND VGND VPWR VPWR _12688_/Y sky130_fd_sc_hd__inv_2
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ _14421_/Y _14426_/X _14400_/X _14426_/X VGND VGND VPWR VPWR _25137_/D sky130_fd_sc_hd__a2bb2o_4
X_17215_ _24369_/Q VGND VGND VPWR VPWR _17215_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15948__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18195_ _18099_/A _18195_/B _18194_/X VGND VGND VPWR VPWR _18196_/C sky130_fd_sc_hd__or3_4
XFILLER_144_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ _14344_/A _14357_/X _25481_/Q _14349_/X VGND VGND VPWR VPWR _25156_/D sky130_fd_sc_hd__o22a_4
X_17146_ _17126_/X VGND VGND VPWR VPWR _17147_/B sky130_fd_sc_hd__inv_2
XFILLER_7_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24154__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12292__A2_N _24836_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13309_ _13345_/A _13305_/X _13308_/X VGND VGND VPWR VPWR _13309_/X sky130_fd_sc_hd__or3_4
XFILLER_116_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17077_ _17026_/A _17076_/X _17053_/X VGND VGND VPWR VPWR _17077_/Y sky130_fd_sc_hd__a21oi_4
X_14289_ _14289_/A _14288_/Y VGND VGND VPWR VPWR _14290_/C sky130_fd_sc_hd__or2_4
XFILLER_171_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16028_ _16027_/Y _16025_/X _15951_/X _16025_/X VGND VGND VPWR VPWR _16028_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_16_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17979_ _18054_/A VGND VGND VPWR VPWR _17979_/X sky130_fd_sc_hd__buf_2
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19718_ _19723_/A VGND VGND VPWR VPWR _19718_/X sky130_fd_sc_hd__buf_2
XANTENNA__19222__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20990_ _20990_/A VGND VGND VPWR VPWR _20990_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16036__B1 _11730_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19649_ _20052_/A _20220_/D _19047_/C VGND VGND VPWR VPWR _19650_/A sky130_fd_sc_hd__or3_4
XFILLER_25_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21580__A1 _14932_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23306__C1 _23305_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22660_ _22660_/A VGND VGND VPWR VPWR _22660_/Y sky130_fd_sc_hd__inv_2
XFILLER_240_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24995__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21611_ _21756_/A _21611_/B VGND VGND VPWR VPWR _21612_/C sky130_fd_sc_hd__or2_4
XFILLER_178_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22591_ _16507_/A _22432_/X _22536_/X VGND VGND VPWR VPWR _22591_/X sky130_fd_sc_hd__o21a_4
XFILLER_21_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21332__A1 _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24924__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24330_ _24326_/CLK _24330_/D HRESETn VGND VGND VPWR VPWR _24330_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_178_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21542_ _21030_/A VGND VGND VPWR VPWR _21542_/X sky130_fd_sc_hd__buf_2
XFILLER_178_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15011__B2 _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24261_ _24263_/CLK _24261_/D HRESETn VGND VGND VPWR VPWR _24261_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_16_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21473_ _21473_/A _19955_/Y VGND VGND VPWR VPWR _21475_/B sky130_fd_sc_hd__or2_4
XFILLER_194_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21579__B _21579_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23212_ _24441_/Q _23138_/X _23001_/X _23211_/X VGND VGND VPWR VPWR _23213_/C sky130_fd_sc_hd__a211o_4
XFILLER_193_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20424_ _20424_/A VGND VGND VPWR VPWR _21396_/B sky130_fd_sc_hd__inv_2
X_24192_ _25466_/CLK _18389_/X HRESETn VGND VGND VPWR VPWR _24192_/Q sky130_fd_sc_hd__dfrtp_4
X_23143_ _23115_/X _23118_/X _23127_/Y _23142_/X VGND VGND VPWR VPWR HRDATA[25] sky130_fd_sc_hd__a211o_4
XFILLER_146_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20355_ _20349_/Y VGND VGND VPWR VPWR _20355_/X sky130_fd_sc_hd__buf_2
XFILLER_161_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21595__A _21748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23074_ _23074_/A _22729_/B VGND VGND VPWR VPWR _23074_/X sky130_fd_sc_hd__or2_4
X_20286_ _18276_/X _19960_/X _18284_/X VGND VGND VPWR VPWR _20286_/X sky130_fd_sc_hd__or3_4
XFILLER_161_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22025_ _22021_/X _22024_/X _21686_/X VGND VGND VPWR VPWR _22025_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_103_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11990_ _11990_/A VGND VGND VPWR VPWR _11990_/Y sky130_fd_sc_hd__inv_2
X_23976_ _23976_/CLK _23976_/D HRESETn VGND VGND VPWR VPWR _17385_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_217_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22927_ _22927_/A _22800_/B VGND VGND VPWR VPWR _22927_/X sky130_fd_sc_hd__or2_4
XFILLER_232_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14937__A _25013_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16041__A1_N _16040_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13841__A _23995_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13660_ _13632_/X VGND VGND VPWR VPWR _13660_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22858_ _22146_/X VGND VGND VPWR VPWR _22858_/X sky130_fd_sc_hd__buf_2
XFILLER_188_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23230__A1_N _17231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16671__A1_N _16670_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_36_0_HCLK clkbuf_7_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_36_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12611_ _12580_/Y _12681_/A _12610_/X VGND VGND VPWR VPWR _12614_/B sky130_fd_sc_hd__or3_4
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21809_ _21809_/A _19888_/Y VGND VGND VPWR VPWR _21811_/B sky130_fd_sc_hd__or2_4
XFILLER_25_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13591_ _18026_/A _13597_/A VGND VGND VPWR VPWR _13592_/B sky130_fd_sc_hd__and2_4
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22789_ _22469_/X VGND VGND VPWR VPWR _22789_/X sky130_fd_sc_hd__buf_2
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_99_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24665__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15330_ _15329_/X VGND VGND VPWR VPWR _25002_/D sky130_fd_sc_hd__inv_2
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12542_ _25419_/Q VGND VGND VPWR VPWR _12664_/A sky130_fd_sc_hd__inv_2
X_24528_ _24558_/CLK _24528_/D HRESETn VGND VGND VPWR VPWR _24528_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20674__A _20678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23936__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15261_ _15261_/A _15261_/B VGND VGND VPWR VPWR _15269_/B sky130_fd_sc_hd__or2_4
XFILLER_157_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23050__A _21427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12473_ _12191_/X _12459_/X _12398_/X _12469_/Y VGND VGND VPWR VPWR _12474_/A sky130_fd_sc_hd__a211o_4
X_24459_ _25021_/CLK _16762_/X HRESETn VGND VGND VPWR VPWR _24459_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23076__A1 _24539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14672__A _14672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14212_ _14212_/A _14212_/B VGND VGND VPWR VPWR _14213_/A sky130_fd_sc_hd__nor2_4
X_17000_ _17000_/A _17000_/B _17000_/C _17000_/D VGND VGND VPWR VPWR _17000_/X sky130_fd_sc_hd__or4_4
XFILLER_172_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15192_ _15192_/A _15190_/A VGND VGND VPWR VPWR _15192_/X sky130_fd_sc_hd__or2_4
XFILLER_137_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_HCLK clkbuf_3_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_14143_ _14142_/X VGND VGND VPWR VPWR _14143_/Y sky130_fd_sc_hd__inv_2
X_14074_ _14008_/A _14070_/X _14067_/X _14007_/B _14073_/X VGND VGND VPWR VPWR _14074_/X
+ sky130_fd_sc_hd__a32o_4
X_18951_ _18951_/A VGND VGND VPWR VPWR _18951_/X sky130_fd_sc_hd__buf_2
XANTENNA__22587__B1 _22586_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13025_ _12342_/A _13024_/Y VGND VGND VPWR VPWR _13025_/X sky130_fd_sc_hd__or2_4
X_17902_ _17738_/X VGND VGND VPWR VPWR _17906_/A sky130_fd_sc_hd__inv_2
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18882_ _23948_/Q _18882_/B VGND VGND VPWR VPWR _20593_/A sky130_fd_sc_hd__or2_4
XFILLER_239_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12920__A _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19452__B1 _19408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16266__B1 _15475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17833_ _17758_/Y _17833_/B VGND VGND VPWR VPWR _17833_/X sky130_fd_sc_hd__or2_4
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19204__B1 _19203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17764_ _17764_/A _16940_/Y _17746_/X _17763_/X VGND VGND VPWR VPWR _17764_/X sky130_fd_sc_hd__or4_4
X_14976_ _14970_/Y VGND VGND VPWR VPWR _14976_/X sky130_fd_sc_hd__buf_2
X_19503_ _19502_/Y VGND VGND VPWR VPWR _19503_/X sky130_fd_sc_hd__buf_2
X_16715_ _24479_/Q VGND VGND VPWR VPWR _16715_/Y sky130_fd_sc_hd__inv_2
X_13927_ _13927_/A _13927_/B VGND VGND VPWR VPWR _13928_/B sky130_fd_sc_hd__nand2_4
XFILLER_207_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17695_ _17695_/A _17694_/X _17688_/C VGND VGND VPWR VPWR _24294_/D sky130_fd_sc_hd__and3_4
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19434_ _19434_/A VGND VGND VPWR VPWR _19447_/A sky130_fd_sc_hd__inv_2
X_16646_ _16645_/Y _16643_/X _16459_/X _16643_/X VGND VGND VPWR VPWR _16646_/X sky130_fd_sc_hd__a2bb2o_4
X_13858_ _25250_/Q _13850_/X _25249_/Q _13852_/X VGND VGND VPWR VPWR _13858_/X sky130_fd_sc_hd__o22a_4
XFILLER_223_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12809_ _12807_/X _24789_/Q _12828_/A _12808_/Y VGND VGND VPWR VPWR _12815_/B sky130_fd_sc_hd__a2bb2o_4
X_19365_ _19117_/A _19163_/B _19026_/C _19026_/D VGND VGND VPWR VPWR _19365_/X sky130_fd_sc_hd__and4_4
X_16577_ _16576_/Y _16572_/X _16402_/X _16572_/X VGND VGND VPWR VPWR _16577_/X sky130_fd_sc_hd__a2bb2o_4
X_13789_ _13787_/Y _13784_/X _13788_/X _13784_/X VGND VGND VPWR VPWR _13789_/X sky130_fd_sc_hd__a2bb2o_4
X_18316_ _18315_/X VGND VGND VPWR VPWR _18316_/Y sky130_fd_sc_hd__inv_2
X_15528_ _21138_/A VGND VGND VPWR VPWR _16446_/C sky130_fd_sc_hd__inv_2
XFILLER_203_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19296_ _19294_/Y _19290_/X _19295_/X _19290_/A VGND VGND VPWR VPWR _19296_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21865__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18247_ _22541_/A _18245_/X _15965_/A _18245_/X VGND VGND VPWR VPWR _24236_/D sky130_fd_sc_hd__a2bb2o_4
X_15459_ _15456_/Y _15458_/X _14400_/X _15458_/X VGND VGND VPWR VPWR _15459_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18054__A _18054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18178_ _18146_/A _18970_/A VGND VGND VPWR VPWR _18179_/C sky130_fd_sc_hd__or2_4
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17129_ _16975_/Y _17128_/X VGND VGND VPWR VPWR _17129_/X sky130_fd_sc_hd__or2_4
X_20140_ _20140_/A VGND VGND VPWR VPWR _20140_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22304__A _22195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23970__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20071_ _23512_/Q VGND VGND VPWR VPWR _20071_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19443__B1 _19351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12830__A _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22023__B _19924_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25123__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23830_ _23831_/CLK _19175_/X VGND VGND VPWR VPWR _23830_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19613__A _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23761_ _23767_/CLK _23761_/D VGND VGND VPWR VPWR _23761_/Q sky130_fd_sc_hd__dfxtp_4
X_20973_ _12131_/A _12147_/A VGND VGND VPWR VPWR _20973_/X sky130_fd_sc_hd__and2_4
XFILLER_38_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13491__B1 _11765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22712_ _22712_/A _22709_/X _22711_/X VGND VGND VPWR VPWR _22712_/X sky130_fd_sc_hd__and3_4
X_25500_ _24209_/CLK _11955_/X HRESETn VGND VGND VPWR VPWR _11940_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23692_ _23427_/CLK _19565_/X VGND VGND VPWR VPWR _23692_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22974__A _21080_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25431_ _25428_/CLK _12620_/Y HRESETn VGND VGND VPWR VPWR _25431_/Q sky130_fd_sc_hd__dfrtp_4
X_22643_ _22758_/A _22643_/B VGND VGND VPWR VPWR _22643_/Y sky130_fd_sc_hd__nor2_4
XFILLER_213_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25362_ _25387_/CLK _13012_/X HRESETn VGND VGND VPWR VPWR _12285_/A sky130_fd_sc_hd__dfrtp_4
X_22574_ _12834_/C _22572_/X _22573_/X VGND VGND VPWR VPWR _22574_/X sky130_fd_sc_hd__o21a_4
XFILLER_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24313_ _24310_/CLK _17626_/Y HRESETn VGND VGND VPWR VPWR _24313_/Q sky130_fd_sc_hd__dfrtp_4
X_21525_ _21525_/A _21524_/X VGND VGND VPWR VPWR _21525_/X sky130_fd_sc_hd__and2_4
X_25293_ _25091_/CLK _25293_/D HRESETn VGND VGND VPWR VPWR _11806_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24005__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24244_ _23890_/CLK _24244_/D HRESETn VGND VGND VPWR VPWR _24244_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21456_ _21463_/A VGND VGND VPWR VPWR _21654_/A sky130_fd_sc_hd__buf_2
XFILLER_31_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20407_ _20407_/A VGND VGND VPWR VPWR _20407_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24175_ _24667_/CLK _18543_/X HRESETn VGND VGND VPWR VPWR _24175_/Q sky130_fd_sc_hd__dfrtp_4
X_21387_ _14681_/A _21384_/X _21386_/X VGND VGND VPWR VPWR _21387_/X sky130_fd_sc_hd__and3_4
XFILLER_123_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23126_ _23120_/X _23122_/X _23123_/X _23125_/X VGND VGND VPWR VPWR _23127_/B sky130_fd_sc_hd__o22a_4
X_20338_ _20338_/A VGND VGND VPWR VPWR _21798_/B sky130_fd_sc_hd__inv_2
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23057_ _16659_/Y _22921_/B VGND VGND VPWR VPWR _23057_/X sky130_fd_sc_hd__and2_4
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20269_ _23440_/Q VGND VGND VPWR VPWR _22259_/B sky130_fd_sc_hd__inv_2
XFILLER_89_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12740__A _12740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16248__B1 _16145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22008_ _22007_/X VGND VGND VPWR VPWR _22024_/A sky130_fd_sc_hd__buf_2
XFILLER_237_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14830_ _14830_/A VGND VGND VPWR VPWR _14830_/X sky130_fd_sc_hd__buf_2
XFILLER_248_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12809__B1 _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14274__A2 _14269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11973_ _11973_/A VGND VGND VPWR VPWR _11973_/Y sky130_fd_sc_hd__inv_2
X_14761_ _13730_/A _14761_/B VGND VGND VPWR VPWR _14762_/C sky130_fd_sc_hd__and2_4
XFILLER_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23959_ _25238_/CLK _20608_/X HRESETn VGND VGND VPWR VPWR _23959_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24846__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16500_ _24561_/Q VGND VGND VPWR VPWR _16500_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13712_ _11803_/Y _13670_/X VGND VGND VPWR VPWR _13712_/Y sky130_fd_sc_hd__nand2_4
XFILLER_189_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14692_ _14692_/A _14714_/A _14704_/A _14692_/D VGND VGND VPWR VPWR _14692_/X sky130_fd_sc_hd__or4_4
X_17480_ _17480_/A VGND VGND VPWR VPWR _17480_/X sky130_fd_sc_hd__buf_2
XANTENNA__22884__A _23171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16431_ _16429_/Y _16426_/X _16349_/X _16430_/X VGND VGND VPWR VPWR _16431_/X sky130_fd_sc_hd__a2bb2o_4
X_13643_ _24039_/Q _13642_/X VGND VGND VPWR VPWR _13644_/B sky130_fd_sc_hd__or2_4
XFILLER_60_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19150_ _19148_/Y _19143_/X _19125_/X _19149_/X VGND VGND VPWR VPWR _23840_/D sky130_fd_sc_hd__a2bb2o_4
X_13574_ _13568_/X _13570_/X _13574_/C _13573_/X VGND VGND VPWR VPWR _13574_/X sky130_fd_sc_hd__or4_4
X_16362_ _16360_/Y _16278_/X _16361_/X _16278_/X VGND VGND VPWR VPWR _16362_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18101_ _15691_/X _18081_/X _18100_/X _24247_/Q _18022_/X VGND VGND VPWR VPWR _18101_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _25409_/Q _24863_/Q _12704_/A _12524_/Y VGND VGND VPWR VPWR _12532_/B sky130_fd_sc_hd__o22a_4
X_15313_ _15313_/A _15307_/B _15312_/X VGND VGND VPWR VPWR _15314_/A sky130_fd_sc_hd__or3_4
X_16293_ _16291_/Y _16292_/X _15567_/X _16292_/X VGND VGND VPWR VPWR _24638_/D sky130_fd_sc_hd__a2bb2o_4
X_19081_ _23863_/Q VGND VGND VPWR VPWR _21894_/B sky130_fd_sc_hd__inv_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_123_0_HCLK clkbuf_7_61_0_HCLK/X VGND VGND VPWR VPWR _24910_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__12915__A _12801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18032_ _18032_/A _18032_/B VGND VGND VPWR VPWR _18034_/B sky130_fd_sc_hd__or2_4
Xclkbuf_8_186_0_HCLK clkbuf_7_93_0_HCLK/X VGND VGND VPWR VPWR _23951_/CLK sky130_fd_sc_hd__clkbuf_1
X_12456_ _12184_/Y _12370_/X VGND VGND VPWR VPWR _12456_/X sky130_fd_sc_hd__or2_4
X_15244_ _15244_/A _15244_/B VGND VGND VPWR VPWR _15261_/B sky130_fd_sc_hd__or2_4
XFILLER_138_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15175_ _15168_/A _15173_/A VGND VGND VPWR VPWR _15176_/C sky130_fd_sc_hd__or2_4
X_12387_ _12204_/A _12386_/Y VGND VGND VPWR VPWR _12387_/X sky130_fd_sc_hd__or2_4
XFILLER_207_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14126_ _14099_/X _14124_/X _25142_/Q _14125_/X VGND VGND VPWR VPWR _14126_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_181_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19983_ _19983_/A VGND VGND VPWR VPWR _19983_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14057_ _14028_/B _14054_/X _14046_/X _13989_/X _14055_/X VGND VGND VPWR VPWR _14057_/X
+ sky130_fd_sc_hd__a32o_4
X_18934_ _18947_/A VGND VGND VPWR VPWR _18934_/X sky130_fd_sc_hd__buf_2
XFILLER_140_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12650__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13008_ _13059_/A _13000_/D VGND VGND VPWR VPWR _13008_/X sky130_fd_sc_hd__or2_4
XFILLER_95_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18865_ _16469_/A _18697_/A _16485_/A _18658_/Y VGND VGND VPWR VPWR _18865_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21783__A1 _21766_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22778__B _22654_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17816_ _24279_/Q _17816_/B VGND VGND VPWR VPWR _17818_/B sky130_fd_sc_hd__or2_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18796_ _18795_/X VGND VGND VPWR VPWR _18796_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17747_ _17747_/A VGND VGND VPWR VPWR _17747_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14959_ _25030_/Q VGND VGND VPWR VPWR _14995_/A sky130_fd_sc_hd__inv_2
XFILLER_47_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21535__A1 _16637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17739__B1 _17704_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24587__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21535__B2 _21336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17678_ _17682_/A _17671_/X _17678_/C VGND VGND VPWR VPWR _17678_/X sky130_fd_sc_hd__and3_4
XFILLER_62_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24516__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19417_ _19416_/Y _19413_/X _19392_/X _19413_/X VGND VGND VPWR VPWR _23745_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16629_ _16629_/A VGND VGND VPWR VPWR _16629_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17888__A _21059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23288__B2 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16792__A _16792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19348_ _19343_/A VGND VGND VPWR VPWR _19348_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_82_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_82_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11787__B1 _11786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19279_ _18981_/A VGND VGND VPWR VPWR _19279_/X sky130_fd_sc_hd__buf_2
XFILLER_175_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21310_ _24613_/Q _21309_/X VGND VGND VPWR VPWR _21310_/X sky130_fd_sc_hd__or2_4
X_22290_ _22290_/A VGND VGND VPWR VPWR _22290_/X sky130_fd_sc_hd__buf_2
XFILLER_190_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16516__A1_N _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21241_ _22069_/A _21238_/X _21241_/C VGND VGND VPWR VPWR _21241_/X sky130_fd_sc_hd__and3_4
XANTENNA__21857__B _21843_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25375__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16478__B1 _16301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21172_ _16789_/Y _21583_/A _11701_/X _21171_/X VGND VGND VPWR VPWR _21172_/X sky130_fd_sc_hd__a211o_4
XFILLER_132_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15855__B _15855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20123_ _20123_/A VGND VGND VPWR VPWR _20123_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16032__A _15988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21873__A _11664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20054_ _20054_/A _20054_/B VGND VGND VPWR VPWR _20055_/A sky130_fd_sc_hd__nand2_4
X_24931_ _25070_/CLK _15527_/X HRESETn VGND VGND VPWR VPWR _21133_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_85_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19343__A _19343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24862_ _25403_/CLK _24862_/D HRESETn VGND VGND VPWR VPWR _24862_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20489__A _20496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15453__A1 _14269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23813_ _23853_/CLK _23813_/D VGND VGND VPWR VPWR _23813_/Q sky130_fd_sc_hd__dfxtp_4
X_24793_ _24795_/CLK _24793_/D HRESETn VGND VGND VPWR VPWR _24793_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _23785_/CLK _23744_/D VGND VGND VPWR VPWR _18037_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ _24065_/Q VGND VGND VPWR VPWR _20956_/Y sky130_fd_sc_hd__inv_2
XPHY_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24257__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_5_31_0_HCLK_A clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _23675_/CLK _19623_/X VGND VGND VPWR VPWR _19622_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _20889_/A VGND VGND VPWR VPWR _20887_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23279__B2 _21871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24912__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17721__A2_N _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22626_ _24659_/Q _22532_/B VGND VGND VPWR VPWR _22629_/B sky130_fd_sc_hd__or2_4
X_25414_ _24508_/CLK _12686_/X HRESETn VGND VGND VPWR VPWR _12684_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_241_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25345_ _25341_/CLK _25345_/D HRESETn VGND VGND VPWR VPWR _12980_/A sky130_fd_sc_hd__dfrtp_4
X_22557_ _22632_/A _22556_/X VGND VGND VPWR VPWR _22557_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12735__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12310_ _12308_/A _12309_/A _12308_/Y _12309_/Y VGND VGND VPWR VPWR _12310_/X sky130_fd_sc_hd__o22a_4
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21508_ _21503_/X _21507_/X _11830_/Y _21503_/X VGND VGND VPWR VPWR _21508_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13290_ _13391_/A _19218_/A VGND VGND VPWR VPWR _13292_/B sky130_fd_sc_hd__or2_4
X_25276_ _25098_/CLK _13773_/X HRESETn VGND VGND VPWR VPWR _25276_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22488_ _24621_/Q _22487_/X VGND VGND VPWR VPWR _22488_/X sky130_fd_sc_hd__or2_4
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12241_ _12240_/Y _12247_/A _25443_/Q _12178_/Y VGND VGND VPWR VPWR _12241_/X sky130_fd_sc_hd__a2bb2o_4
X_24227_ _24227_/CLK _24227_/D HRESETn VGND VGND VPWR VPWR _24227_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21439_ _21075_/Y VGND VGND VPWR VPWR _21439_/X sky130_fd_sc_hd__buf_2
XFILLER_135_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12172_ _12172_/A VGND VGND VPWR VPWR _12172_/Y sky130_fd_sc_hd__inv_2
X_24158_ _24159_/CLK _24158_/D HRESETn VGND VGND VPWR VPWR _24158_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25045__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23109_ _24637_/Q _22904_/X VGND VGND VPWR VPWR _23109_/X sky130_fd_sc_hd__or2_4
X_16980_ _24382_/Q VGND VGND VPWR VPWR _17035_/A sky130_fd_sc_hd__inv_2
X_24089_ _24089_/CLK _20961_/X HRESETn VGND VGND VPWR VPWR RsTx_S1 sky130_fd_sc_hd__dfstp_4
X_15931_ _15930_/Y VGND VGND VPWR VPWR _15931_/X sky130_fd_sc_hd__buf_2
XFILLER_77_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16877__A _14777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18650_ _16562_/Y _18739_/A _16562_/Y _24149_/Q VGND VGND VPWR VPWR _18654_/B sky130_fd_sc_hd__a2bb2o_4
X_15862_ _15861_/X VGND VGND VPWR VPWR _15862_/X sky130_fd_sc_hd__buf_2
X_17601_ _17620_/A _17599_/X _17601_/C VGND VGND VPWR VPWR _24320_/D sky130_fd_sc_hd__and3_4
X_14813_ _14812_/X VGND VGND VPWR VPWR _14814_/B sky130_fd_sc_hd__inv_2
X_18581_ _18577_/B _18581_/B _18593_/C VGND VGND VPWR VPWR _18581_/X sky130_fd_sc_hd__and3_4
X_15793_ _15792_/X VGND VGND VPWR VPWR _15793_/X sky130_fd_sc_hd__buf_2
XANTENNA__21517__A1 _21502_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12258__B2 _24751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24680__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17532_ _11741_/Y _24303_/Q _11741_/Y _24303_/Q VGND VGND VPWR VPWR _17532_/X sky130_fd_sc_hd__a2bb2o_4
X_14744_ _22212_/A VGND VGND VPWR VPWR _14744_/X sky130_fd_sc_hd__buf_2
XFILLER_233_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11956_ _11929_/X _11938_/A VGND VGND VPWR VPWR _11956_/X sky130_fd_sc_hd__or2_4
XANTENNA__17197__B2 _17242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17463_ _24208_/Q VGND VGND VPWR VPWR _20220_/A sky130_fd_sc_hd__buf_2
XFILLER_199_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11887_ _11849_/A _11886_/X _11884_/Y VGND VGND VPWR VPWR _11887_/X sky130_fd_sc_hd__o21a_4
X_14675_ _13744_/X _14675_/B VGND VGND VPWR VPWR _14692_/A sky130_fd_sc_hd__nor2_4
XFILLER_220_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16944__B2 _24288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19202_ _18193_/B VGND VGND VPWR VPWR _19202_/Y sky130_fd_sc_hd__inv_2
X_16414_ _16413_/Y _16411_/X _16233_/X _16411_/X VGND VGND VPWR VPWR _24593_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13626_ _13525_/Y _13620_/X _14610_/A VGND VGND VPWR VPWR _25302_/D sky130_fd_sc_hd__a21oi_4
XFILLER_232_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17394_ _17394_/A _17394_/B VGND VGND VPWR VPWR _17394_/X sky130_fd_sc_hd__or2_4
X_19133_ _19133_/A VGND VGND VPWR VPWR _19133_/X sky130_fd_sc_hd__buf_2
X_16345_ _16343_/Y _16344_/X _16059_/X _16344_/X VGND VGND VPWR VPWR _24618_/D sky130_fd_sc_hd__a2bb2o_4
X_13557_ _13555_/A VGND VGND VPWR VPWR _14570_/A sky130_fd_sc_hd__inv_2
XANTENNA__19894__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12508_ _12508_/A VGND VGND VPWR VPWR _12509_/A sky130_fd_sc_hd__inv_2
X_19064_ _19061_/Y _19062_/X _19063_/X _19062_/X VGND VGND VPWR VPWR _23869_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13488_ _13499_/A VGND VGND VPWR VPWR _13488_/X sky130_fd_sc_hd__buf_2
X_16276_ _22505_/B _15986_/Y VGND VGND VPWR VPWR _16277_/A sky130_fd_sc_hd__and2_4
XFILLER_157_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18015_ _18056_/A _18015_/B _18014_/X VGND VGND VPWR VPWR _18015_/X sky130_fd_sc_hd__and3_4
XFILLER_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12439_ _12439_/A VGND VGND VPWR VPWR _25449_/D sky130_fd_sc_hd__inv_2
X_15227_ _15229_/B VGND VGND VPWR VPWR _15228_/B sky130_fd_sc_hd__inv_2
XANTENNA__15956__A _15924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15158_ _15116_/X _15157_/X VGND VGND VPWR VPWR _15242_/B sky130_fd_sc_hd__or2_4
XFILLER_154_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14109_ _14094_/Y _14108_/X VGND VGND VPWR VPWR _14109_/Y sky130_fd_sc_hd__nor2_4
XFILLER_141_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15089_ _15089_/A _15089_/B _15086_/X _15089_/D VGND VGND VPWR VPWR _15116_/B sky130_fd_sc_hd__or4_4
X_19966_ _23553_/Q VGND VGND VPWR VPWR _22247_/B sky130_fd_sc_hd__inv_2
XFILLER_87_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12380__A _12204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22789__A _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18917_ _18917_/A VGND VGND VPWR VPWR _18917_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21693__A _17704_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19897_ _19897_/A VGND VGND VPWR VPWR _22386_/B sky130_fd_sc_hd__inv_2
XFILLER_234_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16787__A _18951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24768__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18848_ _16492_/Y _24143_/Q _24568_/Q _18613_/X VGND VGND VPWR VPWR _18848_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18779_ _18752_/A _18779_/B _18779_/C VGND VGND VPWR VPWR _18779_/X sky130_fd_sc_hd__and3_4
XFILLER_242_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20810_ _20810_/A _20810_/B VGND VGND VPWR VPWR _20810_/X sky130_fd_sc_hd__and2_4
X_21790_ _21783_/Y _21789_/Y _13772_/C VGND VGND VPWR VPWR _21790_/X sky130_fd_sc_hd__o21a_4
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24350__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20741_ _13121_/B VGND VGND VPWR VPWR _20741_/Y sky130_fd_sc_hd__inv_2
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22720__A3 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16935__B2 _16895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23460_ _24252_/CLK _20216_/X VGND VGND VPWR VPWR _18171_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__17411__A _21368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20672_ _20672_/A _20671_/X VGND VGND VPWR VPWR _23988_/D sky130_fd_sc_hd__nor2_4
XFILLER_149_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22411_ _22274_/X _22410_/X _22138_/C _24827_/Q _21082_/X VGND VGND VPWR VPWR _22411_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23391_ _23391_/CLK _23391_/D VGND VGND VPWR VPWR _13206_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_149_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16027__A _24734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25130_ _25117_/CLK _25130_/D HRESETn VGND VGND VPWR VPWR _25130_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22342_ _22338_/X _22341_/X _17725_/A VGND VGND VPWR VPWR _22342_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_176_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21868__A _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17360__A1 _17352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25061_ _23494_/CLK _25061_/D HRESETn VGND VGND VPWR VPWR _25061_/Q sky130_fd_sc_hd__dfrtp_4
X_22273_ _21289_/X VGND VGND VPWR VPWR _22725_/A sky130_fd_sc_hd__buf_2
XANTENNA__19637__B1 _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24012_ _24049_/CLK _24012_/D HRESETn VGND VGND VPWR VPWR _20727_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_26_0_HCLK clkbuf_8_26_0_HCLK/A VGND VGND VPWR VPWR _23555_/CLK sky130_fd_sc_hd__clkbuf_1
X_21224_ _21224_/A _21154_/X _21224_/C _21223_/X VGND VGND VPWR VPWR _21224_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_89_0_HCLK clkbuf_7_44_0_HCLK/X VGND VGND VPWR VPWR _25397_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_105_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12799__A1_N _12838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21155_ _14264_/Y _21155_/B VGND VGND VPWR VPWR _21155_/X sky130_fd_sc_hd__or2_4
XFILLER_120_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20106_ _16875_/A VGND VGND VPWR VPWR _20106_/X sky130_fd_sc_hd__buf_2
X_21086_ _15851_/X VGND VGND VPWR VPWR _21087_/A sky130_fd_sc_hd__buf_2
XANTENNA__12488__A1 _12252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21747__A1 _21597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20037_ _20036_/Y _20034_/X _19810_/X _20034_/X VGND VGND VPWR VPWR _23529_/D sky130_fd_sc_hd__a2bb2o_4
X_24914_ _24508_/CLK _24914_/D HRESETn VGND VGND VPWR VPWR _24914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_219_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23307__B _22658_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24438__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24845_ _25390_/CLK _15799_/X HRESETn VGND VGND VPWR VPWR _24845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/A VGND VGND VPWR VPWR _11810_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12837_/B VGND VGND VPWR VPWR _12912_/A sky130_fd_sc_hd__buf_2
XPHY_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _21510_/X _21917_/X _21957_/X _21972_/Y _21987_/Y VGND VGND VPWR VPWR _21989_/A
+ sky130_fd_sc_hd__a32o_4
X_24776_ _24765_/CLK _24776_/D HRESETn VGND VGND VPWR VPWR _23216_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24091__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _25532_/Q VGND VGND VPWR VPWR _11741_/Y sky130_fd_sc_hd__inv_2
X_20939_ _20941_/A VGND VGND VPWR VPWR _20939_/Y sky130_fd_sc_hd__inv_2
X_23727_ _23437_/CLK _23727_/D VGND VGND VPWR VPWR _19465_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_215_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24020__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _24942_/Q _24941_/Q _24940_/Q _24939_/Q VGND VGND VPWR VPWR _11672_/X sky130_fd_sc_hd__or4_4
X_14460_ _14459_/Y _14455_/X _14389_/X _14455_/A VGND VGND VPWR VPWR _25122_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23658_ _25326_/CLK _19674_/X VGND VGND VPWR VPWR _13141_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ _13312_/A _13411_/B VGND VGND VPWR VPWR _13412_/C sky130_fd_sc_hd__or2_4
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _20606_/A VGND VGND VPWR VPWR _14391_/Y sky130_fd_sc_hd__inv_2
X_22609_ _22609_/A VGND VGND VPWR VPWR _22609_/Y sky130_fd_sc_hd__inv_2
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23589_ _24297_/CLK _19870_/X VGND VGND VPWR VPWR _19868_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__25297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13342_ _13374_/A _23790_/Q VGND VGND VPWR VPWR _13344_/B sky130_fd_sc_hd__or2_4
X_16130_ _16128_/Y _16124_/X _11735_/X _16129_/X VGND VGND VPWR VPWR _16130_/X sky130_fd_sc_hd__a2bb2o_4
X_25328_ _23458_/CLK _13387_/X HRESETn VGND VGND VPWR VPWR _25328_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13273_ _13438_/A _13273_/B VGND VGND VPWR VPWR _13273_/X sky130_fd_sc_hd__or2_4
X_16061_ _24721_/Q VGND VGND VPWR VPWR _16061_/Y sky130_fd_sc_hd__inv_2
X_25259_ _25260_/CLK _25259_/D HRESETn VGND VGND VPWR VPWR _13536_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19628__B1 _19414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12224_ _12418_/B _24760_/Q _12275_/B _24760_/Q VGND VGND VPWR VPWR _12224_/X sky130_fd_sc_hd__a2bb2o_4
X_15012_ _24476_/Q VGND VGND VPWR VPWR _15012_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19820_ _19820_/A VGND VGND VPWR VPWR _19820_/X sky130_fd_sc_hd__buf_2
XFILLER_151_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12155_ _12109_/A _12153_/Y _12154_/X _12149_/X VGND VGND VPWR VPWR _12155_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17991__A _17999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19751_ _23630_/Q VGND VGND VPWR VPWR _19751_/Y sky130_fd_sc_hd__inv_2
X_12086_ _12086_/A VGND VGND VPWR VPWR _12086_/X sky130_fd_sc_hd__buf_2
X_16963_ _24726_/Q _17038_/D _16006_/Y _17023_/A VGND VGND VPWR VPWR _16963_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24861__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18702_ _18703_/A _18703_/B VGND VGND VPWR VPWR _18704_/B sky130_fd_sc_hd__or2_4
XFILLER_238_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15914_ _15673_/X _15913_/Y _15680_/A _15913_/Y VGND VGND VPWR VPWR _24784_/D sky130_fd_sc_hd__a2bb2o_4
X_19682_ _13340_/B VGND VGND VPWR VPWR _19682_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16894_ _24268_/Q VGND VGND VPWR VPWR _16895_/A sky130_fd_sc_hd__inv_2
XANTENNA__16400__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24179__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16614__B1 _16353_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18633_ _18633_/A VGND VGND VPWR VPWR _18789_/A sky130_fd_sc_hd__buf_2
XFILLER_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15845_ _15845_/A VGND VGND VPWR VPWR _21583_/A sky130_fd_sc_hd__inv_2
XFILLER_209_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24108__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18564_ _18471_/D _18579_/B VGND VGND VPWR VPWR _18577_/B sky130_fd_sc_hd__or2_4
XANTENNA__19711__A _19360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15776_ _15544_/Y _15665_/X _15770_/X _13129_/A _15775_/X VGND VGND VPWR VPWR _24852_/D
+ sky130_fd_sc_hd__a32o_4
X_12988_ _13005_/A _12987_/X VGND VGND VPWR VPWR _13000_/D sky130_fd_sc_hd__or2_4
XFILLER_220_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12100__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17515_ _17508_/X _17515_/B _17512_/X _17515_/D VGND VGND VPWR VPWR _17526_/C sky130_fd_sc_hd__or4_4
XFILLER_33_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14727_ _14720_/A _14701_/A _14726_/X VGND VGND VPWR VPWR _14727_/X sky130_fd_sc_hd__a21o_4
XFILLER_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11939_ _11929_/X _11935_/X _18901_/A _11938_/X VGND VGND VPWR VPWR _25502_/D sky130_fd_sc_hd__o22a_4
X_18495_ _24187_/Q _18495_/B VGND VGND VPWR VPWR _18497_/B sky130_fd_sc_hd__or2_4
XFILLER_33_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17446_ _14364_/A _21176_/A VGND VGND VPWR VPWR _17446_/X sky130_fd_sc_hd__or2_4
XFILLER_205_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14658_ _19116_/A VGND VGND VPWR VPWR _19411_/A sky130_fd_sc_hd__buf_2
XFILLER_177_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13609_ _18060_/A _13608_/X _18060_/A _13608_/X VGND VGND VPWR VPWR _13609_/X sky130_fd_sc_hd__a2bb2o_4
X_17377_ _17242_/B _17374_/B VGND VGND VPWR VPWR _17377_/Y sky130_fd_sc_hd__nand2_4
XFILLER_220_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14589_ _14554_/X _14587_/Y _14588_/X _14579_/X _13535_/A VGND VGND VPWR VPWR _14589_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_174_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12375__A _12167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25131__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19116_ _19116_/A _19116_/B _14648_/A VGND VGND VPWR VPWR _19320_/C sky130_fd_sc_hd__or3_4
X_16328_ _16327_/Y _16325_/X _16233_/X _16325_/X VGND VGND VPWR VPWR _16328_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21688__A _21954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25194__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19047_ _19209_/A _19094_/B _19047_/C VGND VGND VPWR VPWR _19047_/X sky130_fd_sc_hd__or3_4
X_16259_ _24650_/Q VGND VGND VPWR VPWR _16259_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_242_0_HCLK clkbuf_8_243_0_HCLK/A VGND VGND VPWR VPWR _24148_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_161_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24949__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16853__B1 _16716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19949_ _19948_/Y _19946_/X _19610_/X _19946_/X VGND VGND VPWR VPWR _19949_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22960_ _12810_/Y _21437_/X _22849_/X _12572_/Y _21085_/X VGND VGND VPWR VPWR _22960_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__24531__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21911_ _21911_/A _21909_/X _21910_/X VGND VGND VPWR VPWR _21911_/X sky130_fd_sc_hd__and3_4
XFILLER_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22891_ _22891_/A VGND VGND VPWR VPWR _22891_/X sky130_fd_sc_hd__buf_2
XFILLER_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21842_ _21842_/A _22932_/A VGND VGND VPWR VPWR _21842_/X sky130_fd_sc_hd__or2_4
X_24630_ _24623_/CLK _16314_/X HRESETn VGND VGND VPWR VPWR _24630_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22154__A1 _15704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22154__B2 _23138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12269__B _12211_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23351__B1 _25546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24561_ _24558_/CLK _16502_/X HRESETn VGND VGND VPWR VPWR _24561_/Q sky130_fd_sc_hd__dfrtp_4
X_21773_ _21247_/X VGND VGND VPWR VPWR _21773_/X sky130_fd_sc_hd__buf_2
XFILLER_224_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20724_ _20722_/A _20718_/A _20723_/X VGND VGND VPWR VPWR _20724_/Y sky130_fd_sc_hd__a21oi_4
X_23512_ _23528_/CLK _20073_/X VGND VGND VPWR VPWR _23512_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24492_ _24487_/CLK _24492_/D HRESETn VGND VGND VPWR VPWR _16684_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23443_ _23499_/CLK _20260_/X VGND VGND VPWR VPWR _23443_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20655_ _20655_/A VGND VGND VPWR VPWR _23983_/D sky130_fd_sc_hd__inv_2
XANTENNA__15592__B1 _11721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25390__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_52_0_HCLK clkbuf_5_26_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23374_ _24907_/CLK _20684_/A VGND VGND VPWR VPWR _13128_/A sky130_fd_sc_hd__dfxtp_4
X_20586_ _14412_/Y _20566_/X _20556_/X _20585_/X VGND VGND VPWR VPWR _20586_/X sky130_fd_sc_hd__a211o_4
XFILLER_149_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22325_ _21569_/A _22323_/X _21575_/A _22324_/X VGND VGND VPWR VPWR _22325_/X sky130_fd_sc_hd__o22a_4
X_25113_ _25113_/CLK _14488_/X HRESETn VGND VGND VPWR VPWR _25113_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12158__B1 SCLK_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25044_ _25056_/CLK _25044_/D HRESETn VGND VGND VPWR VPWR _25044_/Q sky130_fd_sc_hd__dfrtp_4
X_22256_ _22007_/X _22256_/B _22255_/X VGND VGND VPWR VPWR _22257_/C sky130_fd_sc_hd__and3_4
XFILLER_180_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21207_ _21207_/A _21207_/B _21206_/X VGND VGND VPWR VPWR _21207_/X sky130_fd_sc_hd__and3_4
XFILLER_133_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22187_ _22181_/X _22183_/Y _22185_/Y _22186_/X _21556_/Y VGND VGND VPWR VPWR _22187_/X
+ sky130_fd_sc_hd__o41a_4
XANTENNA__24619__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21138_ _21138_/A _17436_/C _14395_/A _13800_/X VGND VGND VPWR VPWR _21348_/A sky130_fd_sc_hd__or4_4
XFILLER_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13960_ _13959_/X VGND VGND VPWR VPWR _13960_/Y sky130_fd_sc_hd__inv_2
X_21069_ _21736_/A _21068_/Y _24713_/Q _21736_/A VGND VGND VPWR VPWR _21069_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24272__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14659__B _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12911_ _12911_/A VGND VGND VPWR VPWR _25384_/D sky130_fd_sc_hd__inv_2
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13891_ _13934_/C VGND VGND VPWR VPWR _13894_/B sky130_fd_sc_hd__inv_2
XFILLER_246_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12881__A1 _12759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24201__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15630_ _24895_/Q VGND VGND VPWR VPWR _21593_/A sky130_fd_sc_hd__inv_2
X_12842_ _12744_/Y _12842_/B VGND VGND VPWR VPWR _12842_/X sky130_fd_sc_hd__or2_4
X_24828_ _25344_/CLK _24828_/D HRESETn VGND VGND VPWR VPWR _24828_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15561_ _15553_/A VGND VGND VPWR VPWR _15561_/X sky130_fd_sc_hd__buf_2
X_12773_ _22482_/A VGND VGND VPWR VPWR _12773_/Y sky130_fd_sc_hd__inv_2
X_24759_ _24800_/CLK _15963_/X HRESETn VGND VGND VPWR VPWR _22597_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_199_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13830__B1 _13829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17253_/X _17264_/X _17219_/Y VGND VGND VPWR VPWR _17300_/X sky130_fd_sc_hd__o21a_4
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14510_/X _14511_/X _14467_/A _14506_/X VGND VGND VPWR VPWR _25107_/D sky130_fd_sc_hd__o22a_4
XFILLER_199_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11724_ _11720_/Y _11714_/X _11721_/X _11723_/X VGND VGND VPWR VPWR _25537_/D sky130_fd_sc_hd__a2bb2o_4
X_18280_ _18280_/A _17706_/X _18280_/C _18279_/X VGND VGND VPWR VPWR _18280_/X sky130_fd_sc_hd__and4_4
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _14178_/B _15489_/X HADDR[20] _15489_/X VGND VGND VPWR VPWR _15492_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17215_/Y VGND VGND VPWR VPWR _17231_/X sky130_fd_sc_hd__buf_2
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _15636_/A VGND VGND VPWR VPWR _15984_/A sky130_fd_sc_hd__buf_2
X_14443_ _14455_/A VGND VGND VPWR VPWR _14443_/X sky130_fd_sc_hd__buf_2
XFILLER_80_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17162_ _17161_/X VGND VGND VPWR VPWR _24373_/D sky130_fd_sc_hd__inv_2
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14374_ _20467_/A _14371_/X _13824_/X _14373_/X VGND VGND VPWR VPWR _25153_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17324__A1 _17314_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25060__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16113_ _24701_/Q VGND VGND VPWR VPWR _16113_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21301__A _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13325_ _13389_/A _23854_/Q VGND VGND VPWR VPWR _13326_/C sky130_fd_sc_hd__or2_4
XANTENNA__15335__B1 _15334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17093_ _17032_/A _17091_/A VGND VGND VPWR VPWR _17093_/X sky130_fd_sc_hd__or2_4
XFILLER_171_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12923__A _22667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16044_ _24727_/Q VGND VGND VPWR VPWR _16044_/Y sky130_fd_sc_hd__inv_2
X_13256_ _13363_/A _13256_/B VGND VGND VPWR VPWR _13256_/X sky130_fd_sc_hd__or2_4
XFILLER_143_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ _12207_/A VGND VGND VPWR VPWR _12208_/A sky130_fd_sc_hd__inv_2
XFILLER_170_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13187_ _13187_/A VGND VGND VPWR VPWR _13293_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_72_0_HCLK clkbuf_7_36_0_HCLK/X VGND VGND VPWR VPWR _24737_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16835__B1 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12138_ _12092_/Y _12137_/X _12092_/Y _12137_/X VGND VGND VPWR VPWR _12145_/B sky130_fd_sc_hd__a2bb2o_4
X_19803_ _13745_/A _13724_/X _13732_/X VGND VGND VPWR VPWR _19803_/X sky130_fd_sc_hd__or3_4
X_17995_ _17990_/X _17992_/X _17994_/X VGND VGND VPWR VPWR _17996_/C sky130_fd_sc_hd__and3_4
XANTENNA__22132__A _24484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12069_ _25482_/Q VGND VGND VPWR VPWR _12069_/Y sky130_fd_sc_hd__inv_2
X_16946_ _23225_/A _16945_/X _16154_/Y _24262_/Q VGND VGND VPWR VPWR _16948_/C sky130_fd_sc_hd__a2bb2o_4
X_19734_ _19733_/Y _19731_/X _19711_/X _19731_/X VGND VGND VPWR VPWR _23636_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19665_ _19663_/Y _19664_/X _19540_/X _19664_/X VGND VGND VPWR VPWR _23661_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16877_ _14777_/X VGND VGND VPWR VPWR _16877_/X sky130_fd_sc_hd__buf_2
XANTENNA__20395__B1 _13829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18616_ _18681_/A VGND VGND VPWR VPWR _18616_/X sky130_fd_sc_hd__buf_2
X_15828_ _12333_/Y _15827_/X _15623_/X _15827_/X VGND VGND VPWR VPWR _24825_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19596_ _23682_/Q VGND VGND VPWR VPWR _19596_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23995__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18547_ _24173_/Q _18547_/B VGND VGND VPWR VPWR _18547_/X sky130_fd_sc_hd__or2_4
X_15759_ _15759_/A VGND VGND VPWR VPWR _15759_/X sky130_fd_sc_hd__buf_2
XANTENNA__22687__A2 _22676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13821__B1 _11753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23924__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14197__A1_N _20517_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18478_ _18478_/A _18478_/B _18477_/X VGND VGND VPWR VPWR _18478_/X sky130_fd_sc_hd__or3_4
XANTENNA__25148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17429_ _17429_/A VGND VGND VPWR VPWR _17429_/X sky130_fd_sc_hd__buf_2
XFILLER_220_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22439__A2 _22417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20440_ _20440_/A VGND VGND VPWR VPWR _20603_/A sky130_fd_sc_hd__buf_2
XANTENNA__17315__A1 _17251_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20371_ _20306_/X _20368_/X _11760_/X _23401_/Q _20370_/X VGND VGND VPWR VPWR _20371_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16305__A _24633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22110_ _20709_/Y _21121_/A VGND VGND VPWR VPWR _22110_/X sky130_fd_sc_hd__or2_4
XFILLER_174_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23090_ _24438_/Q _21542_/X _22098_/X _23089_/X VGND VGND VPWR VPWR _23090_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24783__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22041_ _22041_/A _22040_/X VGND VGND VPWR VPWR _22041_/X sky130_fd_sc_hd__and2_4
XANTENNA__19616__A _19598_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22611__A2 _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24712__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20622__A1 _15468_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23138__A _23138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23992_ _25243_/CLK _23991_/Q HRESETn VGND VGND VPWR VPWR _23992_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22977__A _24633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22943_ _24361_/Q _21058_/X VGND VGND VPWR VPWR _22943_/X sky130_fd_sc_hd__or2_4
XFILLER_217_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22696__B _22696_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22874_ _12187_/Y _22499_/X _24276_/Q _21056_/X VGND VGND VPWR VPWR _22874_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22127__A1 _13772_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24613_ _24662_/CLK _16359_/X HRESETn VGND VGND VPWR VPWR _24613_/Q sky130_fd_sc_hd__dfrtp_4
X_21825_ _21642_/A _21824_/X _24229_/Q _21958_/B VGND VGND VPWR VPWR _21826_/B sky130_fd_sc_hd__o22a_4
XFILLER_36_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13812__B1 _11735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17003__B1 _24744_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21756_ _21756_/A _20189_/Y VGND VGND VPWR VPWR _21756_/X sky130_fd_sc_hd__or2_4
X_24544_ _24574_/CLK _24544_/D HRESETn VGND VGND VPWR VPWR _24544_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25500__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20707_ _20706_/X VGND VGND VPWR VPWR _24007_/D sky130_fd_sc_hd__inv_2
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15565__B1 _15564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21687_ _21682_/X _21685_/X _21686_/X VGND VGND VPWR VPWR _21687_/X sky130_fd_sc_hd__o21a_4
X_24475_ _24477_/CLK _16731_/X HRESETn VGND VGND VPWR VPWR _24475_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_184_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20638_ _20615_/A VGND VGND VPWR VPWR _20638_/X sky130_fd_sc_hd__buf_2
X_23426_ _23675_/CLK _23426_/D VGND VGND VPWR VPWR _20304_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_196_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22217__A _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23357_ VGND VGND VPWR VPWR _23357_/HI scl_o_S5 sky130_fd_sc_hd__conb_1
XANTENNA__13839__A _13839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20569_ _14421_/Y _20566_/X _20557_/X _20568_/X VGND VGND VPWR VPWR _20570_/A sky130_fd_sc_hd__a211o_4
XANTENNA__22850__A2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13110_ _13110_/A _13110_/B VGND VGND VPWR VPWR _13111_/B sky130_fd_sc_hd__nor2_4
X_22308_ _21845_/A _22308_/B _22308_/C VGND VGND VPWR VPWR _22394_/A sky130_fd_sc_hd__and3_4
XFILLER_164_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14090_ _14090_/A _14089_/X _14105_/A VGND VGND VPWR VPWR _14091_/B sky130_fd_sc_hd__or3_4
X_23288_ _12254_/Y _21532_/X _24288_/Q _22493_/X VGND VGND VPWR VPWR _23288_/X sky130_fd_sc_hd__a2bb2o_4
X_13041_ _12976_/C _13041_/B VGND VGND VPWR VPWR _13051_/B sky130_fd_sc_hd__or2_4
X_22239_ _21920_/A VGND VGND VPWR VPWR _22255_/A sky130_fd_sc_hd__buf_2
X_25027_ _25035_/CLK _25027_/D HRESETn VGND VGND VPWR VPWR _25027_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24033__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24453__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16817__B1 HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_59_0_HCLK clkbuf_7_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16800_ _14925_/Y _16794_/X _16459_/X _16799_/X VGND VGND VPWR VPWR _16800_/X sky130_fd_sc_hd__a2bb2o_4
X_17780_ _16913_/A _17780_/B VGND VGND VPWR VPWR _17782_/B sky130_fd_sc_hd__or2_4
X_14992_ _15192_/A _16737_/A _15192_/A _16737_/A VGND VGND VPWR VPWR _14992_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21169__A2 _15662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16731_ _15000_/Y _16726_/X _16459_/X _16730_/X VGND VGND VPWR VPWR _16731_/X sky130_fd_sc_hd__a2bb2o_4
X_13943_ _13943_/A _13934_/C _13935_/A _13943_/D VGND VGND VPWR VPWR _13943_/X sky130_fd_sc_hd__or4_4
XFILLER_101_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19450_ _19449_/Y _19447_/X _19360_/X _19447_/X VGND VGND VPWR VPWR _23732_/D sky130_fd_sc_hd__a2bb2o_4
X_16662_ _16659_/Y _16655_/X _16301_/X _16661_/X VGND VGND VPWR VPWR _24502_/D sky130_fd_sc_hd__a2bb2o_4
X_13874_ _13873_/X VGND VGND VPWR VPWR _13962_/A sky130_fd_sc_hd__buf_2
XFILLER_35_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22118__A1 _21111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18401_ _22548_/A _18400_/Y _16197_/Y _18459_/A VGND VGND VPWR VPWR _18401_/X sky130_fd_sc_hd__a2bb2o_4
X_15613_ _15608_/A VGND VGND VPWR VPWR _15613_/X sky130_fd_sc_hd__buf_2
X_12825_ _12779_/X _12824_/X VGND VGND VPWR VPWR _12825_/X sky130_fd_sc_hd__or2_4
X_19381_ _19379_/Y _19380_/X _19357_/X _19380_/X VGND VGND VPWR VPWR _19381_/X sky130_fd_sc_hd__a2bb2o_4
X_16593_ _16591_/Y _16592_/X _16240_/X _16592_/X VGND VGND VPWR VPWR _24526_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18332_ _19209_/A _18328_/X _19783_/A VGND VGND VPWR VPWR _18332_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_231_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15544_ _15773_/A VGND VGND VPWR VPWR _15544_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21877__B1 _21439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12756_ _12755_/Y VGND VGND VPWR VPWR _12756_/X sky130_fd_sc_hd__buf_2
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21341__A2 _21336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11706_/X VGND VGND VPWR VPWR _11707_/X sky130_fd_sc_hd__buf_2
X_18263_ _13779_/X VGND VGND VPWR VPWR _18263_/X sky130_fd_sc_hd__buf_2
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _16361_/A VGND VGND VPWR VPWR _15475_/X sky130_fd_sc_hd__buf_2
X_12687_ _12553_/Y _12681_/X _12684_/B _12641_/X VGND VGND VPWR VPWR _12687_/X sky130_fd_sc_hd__a211o_4
XFILLER_129_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _16303_/Y _23012_/A _24622_/Q _17347_/C VGND VGND VPWR VPWR _17214_/X sky130_fd_sc_hd__a2bb2o_4
X_14426_ _14431_/A VGND VGND VPWR VPWR _14426_/X sky130_fd_sc_hd__buf_2
XFILLER_30_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18194_ _18098_/A _18194_/B _18193_/X VGND VGND VPWR VPWR _18194_/X sky130_fd_sc_hd__and3_4
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21031__A _22730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17145_ _17128_/X _17143_/Y _17148_/C VGND VGND VPWR VPWR _17145_/X sky130_fd_sc_hd__and3_4
X_14357_ _25156_/Q _14338_/B _25155_/Q _14345_/A VGND VGND VPWR VPWR _14357_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12653__A _12592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13308_ _13268_/X _13308_/B _13307_/X VGND VGND VPWR VPWR _13308_/X sky130_fd_sc_hd__and3_4
XFILLER_143_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17076_ _16973_/Y _17075_/X VGND VGND VPWR VPWR _17076_/X sky130_fd_sc_hd__or2_4
X_14288_ _14288_/A VGND VGND VPWR VPWR _14288_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16027_ _24734_/Q VGND VGND VPWR VPWR _16027_/Y sky130_fd_sc_hd__inv_2
X_13239_ _13350_/A _23617_/Q VGND VGND VPWR VPWR _13239_/X sky130_fd_sc_hd__or2_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24194__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17978_ _14639_/A VGND VGND VPWR VPWR _18054_/A sky130_fd_sc_hd__buf_2
XFILLER_226_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16929_ _16929_/A _16929_/B _16927_/X _16929_/D VGND VGND VPWR VPWR _16929_/X sky130_fd_sc_hd__or4_4
X_19717_ _19716_/X VGND VGND VPWR VPWR _19723_/A sky130_fd_sc_hd__inv_2
XFILLER_38_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19648_ _23666_/Q VGND VGND VPWR VPWR _19648_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25329__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21580__A2 _15704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23306__B1 _23294_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19579_ _19578_/Y _19576_/X _19392_/X _19576_/X VGND VGND VPWR VPWR _19579_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15795__B1 _15560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12828__A _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21610_ _21609_/X _21610_/B VGND VGND VPWR VPWR _21610_/X sky130_fd_sc_hd__or2_4
X_22590_ _22590_/A _16368_/A VGND VGND VPWR VPWR _22590_/X sky130_fd_sc_hd__or2_4
XFILLER_179_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21332__A2 _21325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21541_ _21311_/X VGND VGND VPWR VPWR _21541_/X sky130_fd_sc_hd__buf_2
XFILLER_194_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24260_ _24263_/CLK _24260_/D HRESETn VGND VGND VPWR VPWR _16917_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_178_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21472_ _21472_/A _21472_/B _21472_/C VGND VGND VPWR VPWR _21472_/X sky130_fd_sc_hd__and3_4
XFILLER_166_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23211_ _24473_/Q _23002_/X _23178_/X VGND VGND VPWR VPWR _23211_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24964__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20423_ _21617_/B _20422_/X _19824_/A _20422_/X VGND VGND VPWR VPWR _23379_/D sky130_fd_sc_hd__a2bb2o_4
X_24191_ _25466_/CLK _24191_/D HRESETn VGND VGND VPWR VPWR _24191_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16035__A _16035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23142_ _23182_/A _23131_/Y _23142_/C _23142_/D VGND VGND VPWR VPWR _23142_/X sky130_fd_sc_hd__or4_4
X_20354_ _23407_/Q VGND VGND VPWR VPWR _22033_/B sky130_fd_sc_hd__inv_2
XFILLER_134_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23073_ _23053_/X _23056_/X _23060_/Y _23072_/X VGND VGND VPWR VPWR HRDATA[23] sky130_fd_sc_hd__a211o_4
X_20285_ _23433_/Q VGND VGND VPWR VPWR _22358_/B sky130_fd_sc_hd__inv_2
XFILLER_136_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18250__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22024_ _22024_/A _22024_/B _22024_/C VGND VGND VPWR VPWR _22024_/X sky130_fd_sc_hd__and3_4
XFILLER_88_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11907__A _11897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23975_ _23986_/CLK _20618_/Y HRESETn VGND VGND VPWR VPWR _17385_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22926_ _23062_/A _22926_/B VGND VGND VPWR VPWR _22926_/Y sky130_fd_sc_hd__nor2_4
XFILLER_216_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22857_ _22857_/A _23278_/B VGND VGND VPWR VPWR _22857_/X sky130_fd_sc_hd__or2_4
XFILLER_216_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12610_ _12594_/Y _12503_/Y _12624_/A _12630_/B VGND VGND VPWR VPWR _12610_/X sky130_fd_sc_hd__or4_4
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21808_ _21656_/A _21806_/X _21808_/C VGND VGND VPWR VPWR _21808_/X sky130_fd_sc_hd__and3_4
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13590_ _13590_/A VGND VGND VPWR VPWR _13597_/A sky130_fd_sc_hd__buf_2
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22788_ _16677_/Y _22921_/B VGND VGND VPWR VPWR _22788_/X sky130_fd_sc_hd__and2_4
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12541_ _25403_/Q _24857_/Q _12717_/A _12540_/Y VGND VGND VPWR VPWR _12545_/C sky130_fd_sc_hd__o22a_4
X_24527_ _24558_/CLK _16590_/X HRESETn VGND VGND VPWR VPWR _16589_/A sky130_fd_sc_hd__dfrtp_4
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15538__B1 HADDR[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21739_ _16781_/Y _21579_/B VGND VGND VPWR VPWR _21739_/X sky130_fd_sc_hd__and2_4
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15260_ _15259_/X VGND VGND VPWR VPWR _25016_/D sky130_fd_sc_hd__inv_2
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12472_ _12480_/A _12470_/X _12472_/C VGND VGND VPWR VPWR _12472_/X sky130_fd_sc_hd__and3_4
X_24458_ _24460_/CLK _24458_/D HRESETn VGND VGND VPWR VPWR _16763_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_184_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12367__A2_N _24826_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14211_ _14184_/A VGND VGND VPWR VPWR _14212_/B sky130_fd_sc_hd__buf_2
X_23409_ _23406_/CLK _23409_/D VGND VGND VPWR VPWR _23409_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22284__B1 _22946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_22_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15191_ _25033_/Q _15190_/Y VGND VGND VPWR VPWR _15191_/X sky130_fd_sc_hd__or2_4
XFILLER_165_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24389_ _24315_/CLK _24389_/D HRESETn VGND VGND VPWR VPWR _17027_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24634__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14142_ _14089_/C _14103_/X _14089_/C _14103_/X VGND VGND VPWR VPWR _14142_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_153_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15784__A _15783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14073_ _14073_/A VGND VGND VPWR VPWR _14073_/X sky130_fd_sc_hd__buf_2
X_18950_ _23908_/Q VGND VGND VPWR VPWR _18950_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13024_ _13016_/X VGND VGND VPWR VPWR _13024_/Y sky130_fd_sc_hd__inv_2
X_17901_ _17901_/A VGND VGND VPWR VPWR _17901_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18881_ _23947_/Q _18881_/B VGND VGND VPWR VPWR _18882_/B sky130_fd_sc_hd__or2_4
XANTENNA__23209__C _23208_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17832_ _17831_/X VGND VGND VPWR VPWR _24274_/D sky130_fd_sc_hd__inv_2
XFILLER_239_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17763_ _17811_/D _17763_/B VGND VGND VPWR VPWR _17763_/X sky130_fd_sc_hd__or2_4
XFILLER_248_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14975_ _25014_/Q VGND VGND VPWR VPWR _15265_/A sky130_fd_sc_hd__inv_2
Xclkbuf_8_146_0_HCLK clkbuf_7_73_0_HCLK/X VGND VGND VPWR VPWR _23916_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25493__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16714_ _16713_/Y _16709_/X _16358_/X _16709_/X VGND VGND VPWR VPWR _24480_/D sky130_fd_sc_hd__a2bb2o_4
X_19502_ _19501_/X VGND VGND VPWR VPWR _19502_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13926_ _13944_/A VGND VGND VPWR VPWR _13927_/A sky130_fd_sc_hd__buf_2
X_17694_ _17575_/Y _17697_/A VGND VGND VPWR VPWR _17694_/X sky130_fd_sc_hd__or2_4
XANTENNA__25422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21562__A2 _14182_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18963__B1 _18942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19433_ _19387_/A _13613_/A _19163_/C VGND VGND VPWR VPWR _19434_/A sky130_fd_sc_hd__or3_4
XFILLER_207_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16645_ _16645_/A VGND VGND VPWR VPWR _16645_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21026__A _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13857_ _13841_/X _13855_/X _25192_/Q _13856_/X VGND VGND VPWR VPWR _13857_/X sky130_fd_sc_hd__o22a_4
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12808_ _23219_/A VGND VGND VPWR VPWR _12808_/Y sky130_fd_sc_hd__inv_2
X_19364_ _17949_/B VGND VGND VPWR VPWR _19364_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17537__A1_N _11720_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16576_ _16576_/A VGND VGND VPWR VPWR _16576_/Y sky130_fd_sc_hd__inv_2
X_13788_ _14392_/A VGND VGND VPWR VPWR _13788_/X sky130_fd_sc_hd__buf_2
XFILLER_43_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17518__B2 _17517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18315_ _17732_/Y _18314_/A _24219_/Q _18314_/Y VGND VGND VPWR VPWR _18315_/X sky130_fd_sc_hd__o22a_4
X_15527_ _15526_/Y _15524_/X HADDR[6] _15524_/X VGND VGND VPWR VPWR _15527_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15529__B1 HADDR[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12739_ _12731_/X _12733_/X _12736_/X _12738_/X VGND VGND VPWR VPWR _12779_/A sky130_fd_sc_hd__or4_4
X_19295_ _17440_/A VGND VGND VPWR VPWR _19295_/X sky130_fd_sc_hd__buf_2
XFILLER_175_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18246_ _22584_/A _18236_/X _15748_/X _18245_/X VGND VGND VPWR VPWR _18246_/X sky130_fd_sc_hd__a2bb2o_4
X_15458_ _15458_/A VGND VGND VPWR VPWR _15458_/X sky130_fd_sc_hd__buf_2
X_14409_ _14405_/Y _14398_/X _14407_/X _14408_/X VGND VGND VPWR VPWR _14409_/X sky130_fd_sc_hd__a2bb2o_4
X_18177_ _18113_/A _19449_/A VGND VGND VPWR VPWR _18177_/X sky130_fd_sc_hd__or2_4
XFILLER_175_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15389_ _15106_/Y _15395_/B VGND VGND VPWR VPWR _15390_/B sky130_fd_sc_hd__or2_4
XANTENNA__24375__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17128_ _16957_/Y _17127_/X VGND VGND VPWR VPWR _17128_/X sky130_fd_sc_hd__or2_4
XFILLER_156_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24304__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15694__A _15694_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17059_ _16978_/A _17058_/Y VGND VGND VPWR VPWR _17061_/B sky130_fd_sc_hd__or2_4
XANTENNA__22304__B _22272_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20070_ _22203_/B _20067_/X _19810_/X _20067_/X VGND VGND VPWR VPWR _23513_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12830__B _12781_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20105__A _20088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_42_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_85_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20972_ _12126_/X _20971_/B VGND VGND VPWR VPWR _20972_/X sky130_fd_sc_hd__and2_4
X_23760_ _24088_/CLK _23760_/D VGND VGND VPWR VPWR _23760_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18954__B1 _17440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22711_ _24730_/Q _22416_/B _21118_/X _22710_/X VGND VGND VPWR VPWR _22711_/X sky130_fd_sc_hd__a211o_4
XPHY_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15768__B1 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23691_ _23691_/CLK _23691_/D VGND VGND VPWR VPWR _19566_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25430_ _25428_/CLK _25430_/D HRESETn VGND VGND VPWR VPWR _12623_/A sky130_fd_sc_hd__dfrtp_4
X_22642_ _21592_/A _22640_/X _22111_/X _22641_/X VGND VGND VPWR VPWR _22643_/B sky130_fd_sc_hd__o22a_4
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14440__B1 _14389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12277__B _12240_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22573_ _16895_/X _22435_/A _12267_/Y _21531_/X VGND VGND VPWR VPWR _22573_/X sky130_fd_sc_hd__o22a_4
X_25361_ _25346_/CLK _13015_/Y HRESETn VGND VGND VPWR VPWR _25361_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24312_ _24305_/CLK _24312_/D HRESETn VGND VGND VPWR VPWR _17502_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_194_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21524_ _21520_/X _21521_/X _21522_/X _25522_/Q _22522_/B VGND VGND VPWR VPWR _21524_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25292_ _25292_/CLK _25292_/D HRESETn VGND VGND VPWR VPWR _11804_/A sky130_fd_sc_hd__dfrtp_4
X_21455_ _21208_/A VGND VGND VPWR VPWR _21463_/A sky130_fd_sc_hd__buf_2
X_24243_ _24889_/CLK _18198_/X HRESETn VGND VGND VPWR VPWR _24243_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21069__B2 _21736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15940__B1 _15939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12293__A _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19131__B1 _19106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20406_ _20405_/Y _20401_/X _15643_/X _20389_/A VGND VGND VPWR VPWR _23385_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12754__B1 _12838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24174_ _24667_/CLK _18545_/X HRESETn VGND VGND VPWR VPWR _24174_/Q sky130_fd_sc_hd__dfrtp_4
X_21386_ _21385_/X _21386_/B VGND VGND VPWR VPWR _21386_/X sky130_fd_sc_hd__or2_4
XANTENNA__24045__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20337_ _20336_/Y _20334_/X _19610_/A _20334_/X VGND VGND VPWR VPWR _20337_/X sky130_fd_sc_hd__a2bb2o_4
X_23125_ _15569_/Y _23292_/B VGND VGND VPWR VPWR _23125_/X sky130_fd_sc_hd__and2_4
XANTENNA__23215__C1 _23214_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23056_ _23054_/X _23055_/X _22919_/X VGND VGND VPWR VPWR _23056_/X sky130_fd_sc_hd__or3_4
X_20268_ _22337_/B _20267_/X _19964_/X _20267_/X VGND VGND VPWR VPWR _23441_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22007_ _17707_/X VGND VGND VPWR VPWR _22007_/X sky130_fd_sc_hd__buf_2
X_20199_ _19116_/A _20199_/B _19387_/A _13596_/A VGND VGND VPWR VPWR _20200_/A sky130_fd_sc_hd__or4_4
XFILLER_163_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23326__A _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_219_0_HCLK clkbuf_8_219_0_HCLK/A VGND VGND VPWR VPWR _24419_/CLK sky130_fd_sc_hd__clkbuf_1
X_14760_ _13725_/A VGND VGND VPWR VPWR _14765_/A sky130_fd_sc_hd__buf_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11972_ _11967_/A _11973_/A _11964_/Y _11971_/Y VGND VGND VPWR VPWR _25497_/D sky130_fd_sc_hd__o22a_4
X_23958_ _23958_/CLK _23958_/D HRESETn VGND VGND VPWR VPWR _23958_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_17_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18945__B1 _16783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13711_ _13673_/B _13710_/Y _13708_/X _13701_/X _11823_/A VGND VGND VPWR VPWR _25286_/D
+ sky130_fd_sc_hd__a32o_4
X_22909_ _22909_/A _22909_/B VGND VGND VPWR VPWR _22909_/X sky130_fd_sc_hd__or2_4
X_14691_ _13744_/X _14675_/B VGND VGND VPWR VPWR _14692_/D sky130_fd_sc_hd__and2_4
X_23889_ _23889_/CLK _19009_/X VGND VGND VPWR VPWR _19008_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12468__A _12191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16430_ _16375_/A VGND VGND VPWR VPWR _16430_/X sky130_fd_sc_hd__buf_2
X_13642_ _24038_/Q _13641_/Y VGND VGND VPWR VPWR _13642_/X sky130_fd_sc_hd__or2_4
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24886__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16361_ _16361_/A VGND VGND VPWR VPWR _16361_/X sky130_fd_sc_hd__buf_2
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _25255_/Q _14549_/B _13820_/A _14557_/A VGND VGND VPWR VPWR _13573_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18155__A _18056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18100_ _18132_/A _18089_/X _18100_/C VGND VGND VPWR VPWR _18100_/X sky130_fd_sc_hd__and3_4
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19370__B1 _19279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24815__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15312_ _15304_/X _15320_/D _15150_/Y VGND VGND VPWR VPWR _15312_/X sky130_fd_sc_hd__o21a_4
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ _24863_/Q VGND VGND VPWR VPWR _12524_/Y sky130_fd_sc_hd__inv_2
X_19080_ _22067_/B _19074_/X _16869_/X _19079_/X VGND VGND VPWR VPWR _23864_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _16284_/X VGND VGND VPWR VPWR _16292_/X sky130_fd_sc_hd__buf_2
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18031_ _17999_/A VGND VGND VPWR VPWR _18032_/A sky130_fd_sc_hd__buf_2
X_15243_ _15243_/A _15243_/B VGND VGND VPWR VPWR _15244_/B sky130_fd_sc_hd__or2_4
XFILLER_145_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12455_ _12263_/A VGND VGND VPWR VPWR _12480_/A sky130_fd_sc_hd__buf_2
XFILLER_157_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15174_ _25037_/Q _15173_/Y VGND VGND VPWR VPWR _15174_/X sky130_fd_sc_hd__or2_4
X_12386_ _12385_/X VGND VGND VPWR VPWR _12386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22405__A _22405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14125_ _14115_/A VGND VGND VPWR VPWR _14125_/X sky130_fd_sc_hd__buf_2
X_19982_ _21677_/B _19980_/X _19981_/X _19980_/X VGND VGND VPWR VPWR _19982_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_181_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14056_ _13989_/X _14054_/X _14046_/X _13990_/C _14055_/X VGND VGND VPWR VPWR _14056_/X
+ sky130_fd_sc_hd__a32o_4
X_18933_ _18932_/X VGND VGND VPWR VPWR _18947_/A sky130_fd_sc_hd__inv_2
XFILLER_140_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ _13007_/A VGND VGND VPWR VPWR _13007_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12244__A2_N _24752_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_29_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18864_ _16469_/Y _24152_/Q _16485_/Y _24146_/Q VGND VGND VPWR VPWR _18864_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17815_ _17817_/B VGND VGND VPWR VPWR _17816_/B sky130_fd_sc_hd__inv_2
XFILLER_0_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18795_ _18789_/C _18794_/X _18724_/X _18791_/B VGND VGND VPWR VPWR _18795_/X sky130_fd_sc_hd__a211o_4
XFILLER_95_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22140__A _22140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19189__B1 _19122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13762__A _21283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17746_ _17746_/A _16906_/Y VGND VGND VPWR VPWR _17746_/X sky130_fd_sc_hd__or2_4
X_14958_ _14949_/X _14952_/X _14958_/C _14957_/X VGND VGND VPWR VPWR _14958_/X sky130_fd_sc_hd__or4_4
XFILLER_36_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13909_ _13878_/B VGND VGND VPWR VPWR _13931_/B sky130_fd_sc_hd__buf_2
X_17677_ _17519_/Y _17670_/X VGND VGND VPWR VPWR _17678_/C sky130_fd_sc_hd__nand2_4
X_14889_ _14888_/Y VGND VGND VPWR VPWR _15192_/A sky130_fd_sc_hd__buf_2
XANTENNA__12378__A _12370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16628_ _16628_/A _16631_/A _16632_/B VGND VGND VPWR VPWR _16629_/A sky130_fd_sc_hd__or3_4
X_19416_ _19416_/A VGND VGND VPWR VPWR _19416_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17888__B _17625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20595__A _14083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16792__B _16792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15765__A3 _15764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16559_ _24539_/Q VGND VGND VPWR VPWR _16559_/Y sky130_fd_sc_hd__inv_2
X_19347_ _23768_/Q VGND VGND VPWR VPWR _19347_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22496__B1 _25529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14973__B2 _16796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19361__B1 _19360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24556__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19278_ _23793_/Q VGND VGND VPWR VPWR _19278_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18229_ _15691_/A _18213_/X _18228_/X _24243_/Q _18022_/A VGND VGND VPWR VPWR _18229_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_248_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21240_ _21884_/A _21240_/B VGND VGND VPWR VPWR _21241_/C sky130_fd_sc_hd__or2_4
XANTENNA__21857__C _21741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21171_ _15331_/A _15845_/A _21327_/B VGND VGND VPWR VPWR _21171_/X sky130_fd_sc_hd__and3_4
XFILLER_190_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17409__A _20628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20122_ _20120_/Y _20116_/X _20095_/X _20121_/X VGND VGND VPWR VPWR _23496_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17427__B1 _16783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20053_ _20054_/A VGND VGND VPWR VPWR _20053_/X sky130_fd_sc_hd__buf_2
X_24930_ _23388_/CLK _15529_/X HRESETn VGND VGND VPWR VPWR _14180_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_112_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25344__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24861_ _25409_/CLK _15758_/X HRESETn VGND VGND VPWR VPWR _24861_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23812_ _23873_/CLK _23812_/D VGND VGND VPWR VPWR _19226_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_227_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24792_ _24795_/CLK _24792_/D HRESETn VGND VGND VPWR VPWR _22420_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_38_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23743_ _23785_/CLK _23743_/D VGND VGND VPWR VPWR _23743_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_192_0_HCLK clkbuf_7_96_0_HCLK/X VGND VGND VPWR VPWR _24675_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ _20828_/X _20954_/X _16645_/A _20874_/X VGND VGND VPWR VPWR _20955_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_49_0_HCLK clkbuf_8_49_0_HCLK/A VGND VGND VPWR VPWR _24947_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_199_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23674_ _25326_/CLK _23674_/D VGND VGND VPWR VPWR _13147_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20870_/X _20885_/X _16684_/A _20875_/X VGND VGND VPWR VPWR _24048_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_214_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14413__B1 _14392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25413_ _24032_/CLK _12688_/Y HRESETn VGND VGND VPWR VPWR _12553_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22625_ _22624_/X VGND VGND VPWR VPWR _22650_/B sky130_fd_sc_hd__inv_2
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19352__B1 _19351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24297__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11920__A _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25344_ _25344_/CLK _13081_/X HRESETn VGND VGND VPWR VPWR _25344_/Q sky130_fd_sc_hd__dfrtp_4
X_22556_ _22552_/X _22553_/X _22135_/C _12511_/A _22555_/X VGND VGND VPWR VPWR _22556_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24226__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21507_ _21504_/X _21377_/X _21507_/C VGND VGND VPWR VPWR _21507_/X sky130_fd_sc_hd__and3_4
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25275_ _23388_/CLK _25275_/D HRESETn VGND VGND VPWR VPWR _25275_/Q sky130_fd_sc_hd__dfrtp_4
X_22487_ _21309_/A VGND VGND VPWR VPWR _22487_/X sky130_fd_sc_hd__buf_2
XFILLER_158_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19104__B1 _19057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12240_ _12240_/A VGND VGND VPWR VPWR _12240_/Y sky130_fd_sc_hd__inv_2
X_24226_ _24233_/CLK _18261_/X HRESETn VGND VGND VPWR VPWR _24226_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21438_ _16637_/A _21435_/X _21436_/X _25521_/Q _21437_/X VGND VGND VPWR VPWR _21438_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22225__A _22225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14963__A2_N _24418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12171_ _25439_/Q _12169_/Y _12279_/A _23184_/A VGND VGND VPWR VPWR _12171_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16008__A1_N _16006_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21369_ _21367_/Y _21159_/X _17431_/Y _21722_/B VGND VGND VPWR VPWR _21369_/X sky130_fd_sc_hd__o22a_4
X_24157_ _24080_/CLK _18704_/X HRESETn VGND VGND VPWR VPWR _24157_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17319__A _17179_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23108_ _22543_/A VGND VGND VPWR VPWR _23108_/X sky130_fd_sc_hd__buf_2
X_24088_ _24088_/CLK _20962_/X HRESETn VGND VGND VPWR VPWR RsTx_S0 sky130_fd_sc_hd__dfstp_4
XFILLER_107_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15930_ _15924_/X VGND VGND VPWR VPWR _15930_/Y sky130_fd_sc_hd__inv_2
X_23039_ _23103_/A _23038_/X VGND VGND VPWR VPWR _23039_/X sky130_fd_sc_hd__and2_4
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19534__A _11774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22411__B1 _24827_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25085__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15861_ _15889_/A VGND VGND VPWR VPWR _15861_/X sky130_fd_sc_hd__buf_2
XANTENNA__25014__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17600_ _17516_/Y _17600_/B VGND VGND VPWR VPWR _17601_/C sky130_fd_sc_hd__or2_4
X_14812_ _25052_/Q _14811_/X _14812_/C VGND VGND VPWR VPWR _14812_/X sky130_fd_sc_hd__or3_4
XFILLER_18_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13582__A _19522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18580_ _18580_/A VGND VGND VPWR VPWR _18593_/C sky130_fd_sc_hd__buf_2
X_15792_ _15820_/A VGND VGND VPWR VPWR _15792_/X sky130_fd_sc_hd__buf_2
XFILLER_190_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17531_ _25521_/Q _17580_/C _25525_/Q _17530_/Y VGND VGND VPWR VPWR _17531_/X sky130_fd_sc_hd__a2bb2o_4
X_14743_ _14705_/A VGND VGND VPWR VPWR _22212_/A sky130_fd_sc_hd__buf_2
X_11955_ _11940_/A _11954_/X _11944_/A VGND VGND VPWR VPWR _11955_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19591__B1 _19540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17462_ _13162_/X _17450_/X _18342_/A VGND VGND VPWR VPWR _17462_/X sky130_fd_sc_hd__o21a_4
XFILLER_199_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14674_ _14666_/X _14671_/X _14741_/A VGND VGND VPWR VPWR _14675_/B sky130_fd_sc_hd__o21a_4
XFILLER_60_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11886_ _11849_/B _11883_/Y VGND VGND VPWR VPWR _11886_/X sky130_fd_sc_hd__and2_4
XANTENNA__14404__B1 _14403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15747__A3 _15746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16413_ _24593_/Q VGND VGND VPWR VPWR _16413_/Y sky130_fd_sc_hd__inv_2
X_19201_ _19198_/Y _19199_/X _19200_/X _19199_/X VGND VGND VPWR VPWR _19201_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13625_ _13625_/A VGND VGND VPWR VPWR _14610_/A sky130_fd_sc_hd__buf_2
XFILLER_177_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17393_ _17393_/A _17393_/B VGND VGND VPWR VPWR _17394_/B sky130_fd_sc_hd__or2_4
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19132_ _23845_/Q VGND VGND VPWR VPWR _19132_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22119__B _22119_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16344_ _16344_/A VGND VGND VPWR VPWR _16344_/X sky130_fd_sc_hd__buf_2
X_13556_ _13556_/A VGND VGND VPWR VPWR _13556_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21150__B1 _25170_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_200_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12507_ _12507_/A _12501_/X _12507_/C _12506_/X VGND VGND VPWR VPWR _12507_/X sky130_fd_sc_hd__or4_4
X_19063_ _19063_/A VGND VGND VPWR VPWR _19063_/X sky130_fd_sc_hd__buf_2
X_16275_ _23313_/A VGND VGND VPWR VPWR _16275_/Y sky130_fd_sc_hd__inv_2
X_13487_ _12000_/Y _13485_/X _11757_/X _13485_/X VGND VGND VPWR VPWR _13487_/X sky130_fd_sc_hd__a2bb2o_4
X_18014_ _18014_/A _23841_/Q VGND VGND VPWR VPWR _18014_/X sky130_fd_sc_hd__or2_4
XFILLER_218_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15226_ _15039_/X _15205_/C VGND VGND VPWR VPWR _15229_/B sky130_fd_sc_hd__or2_4
XFILLER_157_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12438_ _12428_/C _12428_/D _12390_/X _12436_/B VGND VGND VPWR VPWR _12439_/A sky130_fd_sc_hd__a211o_4
XANTENNA__22135__A _21303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15157_ _15127_/X _15136_/X _15157_/C _15156_/X VGND VGND VPWR VPWR _15157_/X sky130_fd_sc_hd__or4_4
XANTENNA__23949__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12369_ _12369_/A _12369_/B _12359_/X _12368_/X VGND VGND VPWR VPWR _12370_/B sky130_fd_sc_hd__or4_4
XFILLER_153_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14108_ _14108_/A _14108_/B _14095_/A VGND VGND VPWR VPWR _14108_/X sky130_fd_sc_hd__and3_4
X_15088_ _15087_/Y _24580_/Q _15087_/Y _24580_/Q VGND VGND VPWR VPWR _15089_/D sky130_fd_sc_hd__a2bb2o_4
X_19965_ _22359_/B _19963_/X _19964_/X _19963_/X VGND VGND VPWR VPWR _19965_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12380__B _12264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14039_ _14030_/Y _14032_/Y _14039_/C _14038_/X VGND VGND VPWR VPWR _14039_/X sky130_fd_sc_hd__or4_4
X_18916_ _18915_/Y _18913_/X _17418_/X _18913_/X VGND VGND VPWR VPWR _18916_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21693__B _21649_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19896_ _21184_/B _19891_/X _19874_/X _19878_/Y VGND VGND VPWR VPWR _23579_/D sky130_fd_sc_hd__a2bb2o_4
X_18847_ _24552_/Q _18804_/A _16510_/A _18789_/C VGND VGND VPWR VPWR _18847_/X sky130_fd_sc_hd__a2bb2o_4
X_18778_ _18778_/A _18778_/B VGND VGND VPWR VPWR _18779_/C sky130_fd_sc_hd__or2_4
XFILLER_242_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_202_0_HCLK clkbuf_8_202_0_HCLK/A VGND VGND VPWR VPWR _24980_/CLK sky130_fd_sc_hd__clkbuf_1
X_17729_ _17725_/X _17728_/X _17725_/X _17728_/X VGND VGND VPWR VPWR _17736_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19582__B1 _19395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24737__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_8_0_HCLK clkbuf_7_4_0_HCLK/X VGND VGND VPWR VPWR _23806_/CLK sky130_fd_sc_hd__clkbuf_1
X_20740_ _20731_/X _20739_/X _24904_/Q _20736_/X VGND VGND VPWR VPWR _20740_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16396__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20671_ _14207_/Y _17401_/A _17384_/A _17398_/A VGND VGND VPWR VPWR _20671_/X sky130_fd_sc_hd__o22a_4
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12836__A _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24390__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22410_ _22410_/A _22275_/X VGND VGND VPWR VPWR _22410_/X sky130_fd_sc_hd__or2_4
XFILLER_149_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16148__B1 _16055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23390_ _23912_/CLK _23390_/D VGND VGND VPWR VPWR _13256_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22341_ _21933_/A _22341_/B _22341_/C VGND VGND VPWR VPWR _22341_/X sky130_fd_sc_hd__and3_4
XFILLER_149_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22272_ _22271_/X VGND VGND VPWR VPWR _22272_/Y sky130_fd_sc_hd__inv_2
X_25060_ _23665_/CLK _14770_/X HRESETn VGND VGND VPWR VPWR _25060_/Q sky130_fd_sc_hd__dfrtp_4
X_21223_ _21955_/A _21213_/X _21222_/Y VGND VGND VPWR VPWR _21223_/X sky130_fd_sc_hd__or3_4
X_24011_ _24049_/CLK _20726_/Y HRESETn VGND VGND VPWR VPWR _20722_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20491__C _20477_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12185__B2 _21088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25525__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21154_ _17436_/B _21146_/X _12058_/C _21153_/X VGND VGND VPWR VPWR _21154_/X sky130_fd_sc_hd__o22a_4
XFILLER_105_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20105_ _20088_/A VGND VGND VPWR VPWR _20105_/X sky130_fd_sc_hd__buf_2
XANTENNA__23197__B2 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21085_ _22451_/A VGND VGND VPWR VPWR _21085_/X sky130_fd_sc_hd__buf_2
XANTENNA__14882__B1 _15249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20036_ _23529_/Q VGND VGND VPWR VPWR _20036_/Y sky130_fd_sc_hd__inv_2
X_24913_ _24508_/CLK _15585_/X HRESETn VGND VGND VPWR VPWR _15583_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11696__B1 _11695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_12_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_218_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16623__A1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11915__A _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24844_ _25390_/CLK _24844_/D HRESETn VGND VGND VPWR VPWR _12309_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_160_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24775_ _24765_/CLK _15936_/X HRESETn VGND VGND VPWR VPWR _23184_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_61_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21987_ _22041_/A _21986_/X _21510_/X VGND VGND VPWR VPWR _21987_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_160_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23198__A1_N _17175_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24478__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11737_/Y _11733_/X _11739_/X _11733_/X VGND VGND VPWR VPWR _11740_/X sky130_fd_sc_hd__a2bb2o_4
X_23726_ _23437_/CLK _23726_/D VGND VGND VPWR VPWR _23726_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20919_/X _20937_/X _24504_/Q _20923_/X VGND VGND VPWR VPWR _20938_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23323__B _16792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20183__B2 _20180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24407__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _24938_/Q _24937_/Q VGND VGND VPWR VPWR _11671_/X sky130_fd_sc_hd__or2_4
X_23657_ _23665_/CLK _23657_/D VGND VGND VPWR VPWR _13223_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_187_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _20868_/X VGND VGND VPWR VPWR _20869_/Y sky130_fd_sc_hd__inv_2
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19325__B1 _19279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13220_/X _13410_/B VGND VGND VPWR VPWR _13410_/X sky130_fd_sc_hd__or2_4
XFILLER_168_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14664__C _13584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22608_ _21055_/X _22603_/X _21832_/X _22607_/Y VGND VGND VPWR VPWR _22609_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16139__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14390_ _14388_/Y _14383_/X _14389_/X _14372_/X VGND VGND VPWR VPWR _25147_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23588_ _24297_/CLK _19872_/X VGND VGND VPWR VPWR _19871_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12465__B _12191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24060__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13341_ _13219_/X _13339_/X _13341_/C VGND VGND VPWR VPWR _13341_/X sky130_fd_sc_hd__and3_4
X_25327_ _23458_/CLK _25327_/D HRESETn VGND VGND VPWR VPWR _25327_/Q sky130_fd_sc_hd__dfrtp_4
X_22539_ _22539_/A _22539_/B _22539_/C VGND VGND VPWR VPWR _22539_/X sky130_fd_sc_hd__and3_4
XFILLER_139_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16060_ _16057_/Y _16058_/X _16059_/X _16058_/X VGND VGND VPWR VPWR _24722_/D sky130_fd_sc_hd__a2bb2o_4
X_13272_ _13345_/A _13267_/X _13271_/X VGND VGND VPWR VPWR _13272_/X sky130_fd_sc_hd__or3_4
X_25258_ _25325_/CLK _13833_/X HRESETn VGND VGND VPWR VPWR _13559_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15011_ _14886_/A _15010_/Y _15272_/A _16786_/A VGND VGND VPWR VPWR _15011_/X sky130_fd_sc_hd__a2bb2o_4
X_12223_ _12275_/B VGND VGND VPWR VPWR _12418_/B sky130_fd_sc_hd__buf_2
X_24209_ _24209_/CLK _24209_/D HRESETn VGND VGND VPWR VPWR _17460_/A sky130_fd_sc_hd__dfrtp_4
X_25189_ _25249_/CLK _14255_/X HRESETn VGND VGND VPWR VPWR _25189_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12154_ _12154_/A _18372_/B VGND VGND VPWR VPWR _12154_/X sky130_fd_sc_hd__and2_4
XFILLER_150_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19750_ _19749_/Y _19747_/X _19702_/X _19747_/X VGND VGND VPWR VPWR _23631_/D sky130_fd_sc_hd__a2bb2o_4
X_12085_ _21570_/A VGND VGND VPWR VPWR _12086_/A sky130_fd_sc_hd__buf_2
X_16962_ _24383_/Q VGND VGND VPWR VPWR _17038_/D sky130_fd_sc_hd__inv_2
XFILLER_49_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18701_ _18700_/X VGND VGND VPWR VPWR _18703_/B sky130_fd_sc_hd__inv_2
XFILLER_1_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15913_ _15912_/X VGND VGND VPWR VPWR _15913_/Y sky130_fd_sc_hd__inv_2
X_16893_ _16122_/Y _24274_/Q _16122_/Y _24274_/Q VGND VGND VPWR VPWR _16901_/A sky130_fd_sc_hd__a2bb2o_4
X_19681_ _19680_/Y _19678_/X _19534_/X _19678_/X VGND VGND VPWR VPWR _19681_/X sky130_fd_sc_hd__a2bb2o_4
X_15844_ _11676_/B _14442_/A VGND VGND VPWR VPWR _15845_/A sky130_fd_sc_hd__or2_4
X_18632_ _24135_/Q VGND VGND VPWR VPWR _18633_/A sky130_fd_sc_hd__inv_2
XFILLER_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15775_ _15773_/A _15670_/X VGND VGND VPWR VPWR _15775_/X sky130_fd_sc_hd__or2_4
X_18563_ _18563_/A _18563_/B VGND VGND VPWR VPWR _18579_/B sky130_fd_sc_hd__or2_4
XANTENNA__22699__B1 _22468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12987_ _13017_/A _12349_/Y _12987_/C _12986_/X VGND VGND VPWR VPWR _12987_/X sky130_fd_sc_hd__or4_4
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24830__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14726_ _14721_/X _14725_/Y _14718_/Y VGND VGND VPWR VPWR _14726_/X sky130_fd_sc_hd__a21o_4
X_17514_ _25527_/Q _17513_/A _11759_/Y _17513_/Y VGND VGND VPWR VPWR _17515_/D sky130_fd_sc_hd__o22a_4
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11938_ _11938_/A _11938_/B _11945_/A _11940_/A VGND VGND VPWR VPWR _11938_/X sky130_fd_sc_hd__and4_4
X_18494_ _18496_/B VGND VGND VPWR VPWR _18495_/B sky130_fd_sc_hd__inv_2
XANTENNA__16378__B1 _16001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22330__A1_N _20628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24148__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17445_ _15636_/A _15636_/B _11660_/A _12039_/D VGND VGND VPWR VPWR _21176_/A sky130_fd_sc_hd__or4_4
XFILLER_220_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21034__A _22525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14657_ _14648_/A _14656_/X _19002_/B _13588_/X VGND VGND VPWR VPWR _14657_/X sky130_fd_sc_hd__o22a_4
XFILLER_178_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_32_0_HCLK clkbuf_7_16_0_HCLK/X VGND VGND VPWR VPWR _23610_/CLK sky130_fd_sc_hd__clkbuf_1
X_11869_ _11869_/A _11864_/B VGND VGND VPWR VPWR _11869_/Y sky130_fd_sc_hd__nor2_4
XFILLER_232_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19316__B1 _19203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_95_0_HCLK clkbuf_8_95_0_HCLK/A VGND VGND VPWR VPWR _25428_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13608_ _13606_/A _13606_/B _14650_/A VGND VGND VPWR VPWR _13608_/X sky130_fd_sc_hd__a21o_4
X_17376_ _17241_/Y _17374_/X _17375_/Y VGND VGND VPWR VPWR _17376_/X sky130_fd_sc_hd__o21a_4
X_14588_ _14566_/D VGND VGND VPWR VPWR _14588_/X sky130_fd_sc_hd__buf_2
XFILLER_220_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16327_ _24625_/Q VGND VGND VPWR VPWR _16327_/Y sky130_fd_sc_hd__inv_2
X_19115_ _23850_/Q VGND VGND VPWR VPWR _19115_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13539_ _25084_/Q VGND VGND VPWR VPWR _14549_/A sky130_fd_sc_hd__inv_2
XFILLER_9_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19046_ _19046_/A VGND VGND VPWR VPWR _19046_/Y sky130_fd_sc_hd__inv_2
X_16258_ _16256_/Y _16252_/X _15466_/X _16257_/X VGND VGND VPWR VPWR _24651_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17167__A2_N _17366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15209_ _14898_/X _15209_/B VGND VGND VPWR VPWR _15211_/B sky130_fd_sc_hd__or2_4
XFILLER_127_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22623__B1 _22622_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16189_ _23248_/A VGND VGND VPWR VPWR _16189_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16302__B1 _16301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19948_ _19948_/A VGND VGND VPWR VPWR _19948_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24989__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19879_ _19878_/Y VGND VGND VPWR VPWR _19879_/X sky130_fd_sc_hd__buf_2
XANTENNA__24918__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21910_ _21913_/A _20041_/Y VGND VGND VPWR VPWR _21910_/X sky130_fd_sc_hd__or2_4
XANTENNA__11735__A _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22890_ _24598_/Q _22890_/B VGND VGND VPWR VPWR _22890_/X sky130_fd_sc_hd__or2_4
XANTENNA__13419__B2 _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21841_ _21315_/X _21831_/X _21840_/X VGND VGND VPWR VPWR _21841_/X sky130_fd_sc_hd__a21bo_4
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24571__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24560_ _24148_/CLK _16504_/X HRESETn VGND VGND VPWR VPWR _24560_/Q sky130_fd_sc_hd__dfrtp_4
X_21772_ _22380_/A _21772_/B _21772_/C VGND VGND VPWR VPWR _21772_/X sky130_fd_sc_hd__and3_4
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24500__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23511_ _23575_/CLK _20075_/X VGND VGND VPWR VPWR _23511_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20723_ _20723_/A _20718_/Y VGND VGND VPWR VPWR _20723_/X sky130_fd_sc_hd__and2_4
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24491_ _24487_/CLK _16688_/X HRESETn VGND VGND VPWR VPWR _24491_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_196_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16038__A _16038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19307__B1 _19282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23442_ _23972_/CLK _20263_/X VGND VGND VPWR VPWR _23442_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21879__A _21019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20654_ _14224_/Y _20638_/X _20629_/A _20653_/X VGND VGND VPWR VPWR _20655_/A sky130_fd_sc_hd__a211o_4
XFILLER_210_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_3_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_6_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20585_ _18881_/B _20584_/Y _20572_/X VGND VGND VPWR VPWR _20585_/X sky130_fd_sc_hd__and3_4
X_23373_ _23972_/CLK scl_oen_o_S5 VGND VGND VPWR VPWR _20997_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__17795__C _17555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25112_ _23958_/CLK _14493_/X HRESETn VGND VGND VPWR VPWR _25112_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22324_ _12119_/A _12086_/A _18371_/Y _12057_/A VGND VGND VPWR VPWR _22324_/X sky130_fd_sc_hd__o22a_4
XFILLER_137_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25043_ _25043_/CLK _14870_/Y HRESETn VGND VGND VPWR VPWR _14859_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_164_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13397__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22255_ _22255_/A _19922_/Y VGND VGND VPWR VPWR _22255_/X sky130_fd_sc_hd__or2_4
XFILLER_191_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21206_ _21209_/A _21206_/B VGND VGND VPWR VPWR _21206_/X sky130_fd_sc_hd__or2_4
X_22186_ _20510_/A _21849_/X _23968_/Q _21364_/B VGND VGND VPWR VPWR _22186_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22090__B2 _22089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22503__A _15008_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18604__A1_N _16605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21137_ _23927_/Q VGND VGND VPWR VPWR _21137_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21068_ _21068_/A VGND VGND VPWR VPWR _21068_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16944__A2_N _24288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24659__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ _12741_/X _12892_/B _12862_/X _12907_/Y VGND VGND VPWR VPWR _12911_/A sky130_fd_sc_hd__a211o_4
X_20019_ _22016_/B _20013_/X _19970_/X _20018_/X VGND VGND VPWR VPWR _23536_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19794__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13890_ _13898_/B VGND VGND VPWR VPWR _13934_/C sky130_fd_sc_hd__buf_2
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12841_ _12796_/Y _12804_/Y _12841_/C _12841_/D VGND VGND VPWR VPWR _12842_/B sky130_fd_sc_hd__or4_4
X_24827_ _25428_/CLK _15825_/X HRESETn VGND VGND VPWR VPWR _24827_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19546__B1 _19408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13860__A _23995_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15560_ HWDATA[28] VGND VGND VPWR VPWR _15560_/X sky130_fd_sc_hd__buf_2
X_12772_ _12772_/A VGND VGND VPWR VPWR _12834_/A sky130_fd_sc_hd__inv_2
X_24758_ _25369_/CLK _15966_/X HRESETn VGND VGND VPWR VPWR _22558_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_203_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24241__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _25107_/Q _14500_/X _21847_/A _14502_/X VGND VGND VPWR VPWR _14511_/X sky130_fd_sc_hd__o22a_4
XFILLER_199_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11766_/A VGND VGND VPWR VPWR _11723_/X sky130_fd_sc_hd__buf_2
X_23709_ _23691_/CLK _23709_/D VGND VGND VPWR VPWR _23709_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _16364_/A _15489_/X HADDR[21] _15489_/X VGND VGND VPWR VPWR _15491_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24689_ _24744_/CLK _24689_/D HRESETn VGND VGND VPWR VPWR _16144_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_19_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17341_/A VGND VGND VPWR VPWR _17230_/X sky130_fd_sc_hd__buf_2
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14442_/A _14442_/B VGND VGND VPWR VPWR _14455_/A sky130_fd_sc_hd__nor2_4
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _14364_/A VGND VGND VPWR VPWR _16366_/A sky130_fd_sc_hd__buf_2
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16780__B1 _16778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17161_ _17040_/Y _17062_/X _17064_/X _17159_/B VGND VGND VPWR VPWR _17161_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15787__A _15786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14373_ _14372_/X VGND VGND VPWR VPWR _14373_/X sky130_fd_sc_hd__buf_2
XANTENNA__12626__D _12626_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19259__A _19253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16112_ _16110_/Y _16111_/X _16020_/X _16111_/X VGND VGND VPWR VPWR _16112_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _13388_/A _23870_/Q VGND VGND VPWR VPWR _13326_/B sky130_fd_sc_hd__or2_4
X_17092_ _16964_/A _17091_/Y VGND VGND VPWR VPWR _17092_/X sky130_fd_sc_hd__or2_4
XFILLER_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16043_ _16042_/Y _16038_/X _11743_/X _16038_/X VGND VGND VPWR VPWR _24728_/D sky130_fd_sc_hd__a2bb2o_4
X_13255_ _13293_/A _13255_/B _13255_/C VGND VGND VPWR VPWR _13263_/B sky130_fd_sc_hd__or3_4
XFILLER_142_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12206_ _12204_/A _12205_/A _12204_/Y _12205_/Y VGND VGND VPWR VPWR _12214_/B sky130_fd_sc_hd__o22a_4
X_13186_ _13186_/A VGND VGND VPWR VPWR _13186_/X sky130_fd_sc_hd__buf_2
XFILLER_151_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19802_ _23610_/Q VGND VGND VPWR VPWR _22364_/B sky130_fd_sc_hd__inv_2
XFILLER_151_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12137_ _12135_/A _12116_/X _12136_/Y VGND VGND VPWR VPWR _12137_/X sky130_fd_sc_hd__o21a_4
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17994_ _18151_/A _23905_/Q VGND VGND VPWR VPWR _17994_/X sky130_fd_sc_hd__or2_4
X_19733_ _13411_/B VGND VGND VPWR VPWR _19733_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23030__B1 _11694_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12068_ _12067_/Y _12065_/X _11775_/X _12065_/X VGND VGND VPWR VPWR _25483_/D sky130_fd_sc_hd__a2bb2o_4
X_16945_ _16945_/A VGND VGND VPWR VPWR _16945_/X sky130_fd_sc_hd__buf_2
XFILLER_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19785__B1 _18250_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15538__A2_N _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19664_ _19650_/Y VGND VGND VPWR VPWR _19664_/X sky130_fd_sc_hd__buf_2
XFILLER_64_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16876_ _19824_/A VGND VGND VPWR VPWR _16876_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16599__B1 _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24329__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18615_ _16566_/A _18613_/X _24542_/Q _18698_/A VGND VGND VPWR VPWR _18618_/C sky130_fd_sc_hd__a2bb2o_4
X_15827_ _15820_/A VGND VGND VPWR VPWR _15827_/X sky130_fd_sc_hd__buf_2
X_19595_ _19594_/Y _19590_/X _19408_/X _19576_/A VGND VGND VPWR VPWR _19595_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_231_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19537__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17242__A _17241_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15758_ _12502_/Y _15755_/X _15619_/X _15755_/X VGND VGND VPWR VPWR _15758_/X sky130_fd_sc_hd__a2bb2o_4
X_18546_ _18533_/X VGND VGND VPWR VPWR _18547_/B sky130_fd_sc_hd__inv_2
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14709_ _25064_/Q VGND VGND VPWR VPWR _14710_/A sky130_fd_sc_hd__buf_2
X_15689_ _18022_/A VGND VGND VPWR VPWR _15690_/A sky130_fd_sc_hd__inv_2
X_18477_ _18563_/A _18562_/A _18561_/C _18477_/D VGND VGND VPWR VPWR _18477_/X sky130_fd_sc_hd__or4_4
XFILLER_61_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17428_ _24328_/Q VGND VGND VPWR VPWR _21558_/A sky130_fd_sc_hd__inv_2
XANTENNA__16771__B1 _16601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15697__A _14366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23964__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17359_ _17351_/A _17359_/B _17359_/C VGND VGND VPWR VPWR _17359_/X sky130_fd_sc_hd__and3_4
XANTENNA__25188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20370_ _20369_/X VGND VGND VPWR VPWR _20370_/X sky130_fd_sc_hd__buf_2
XFILLER_9_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16523__B1 _16522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19029_ _19024_/Y _19028_/X _19006_/X _19028_/X VGND VGND VPWR VPWR _23882_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22040_ _22393_/A _21999_/Y _22006_/X _21510_/X _22039_/X VGND VGND VPWR VPWR _22040_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_115_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12736__A1_N _25374_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11899__B1 RsRx_S1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23991_ _25243_/CLK sda_i_S5 HRESETn VGND VGND VPWR VPWR _23991_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24752__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22942_ _23251_/A _22939_/X _22941_/X VGND VGND VPWR VPWR _22942_/X sky130_fd_sc_hd__and3_4
XFILLER_217_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24124__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22873_ _22781_/A _22860_/X _22873_/C _22873_/D VGND VGND VPWR VPWR _22873_/X sky130_fd_sc_hd__or4_4
XFILLER_28_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22127__A2 _22090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24612_ _24623_/CLK _16362_/X HRESETn VGND VGND VPWR VPWR _24612_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15801__A2 _15789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21824_ _21643_/X _21823_/X _24224_/Q _21278_/X VGND VGND VPWR VPWR _21824_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24543_ _24574_/CLK _16551_/X HRESETn VGND VGND VPWR VPWR _16550_/A sky130_fd_sc_hd__dfrtp_4
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21755_ _21609_/X _21755_/B VGND VGND VPWR VPWR _21755_/X sky130_fd_sc_hd__or2_4
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20706_ _15625_/Y _20687_/X _20696_/X _20705_/Y VGND VGND VPWR VPWR _20706_/X sky130_fd_sc_hd__o22a_4
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24474_ _24477_/CLK _16733_/X HRESETn VGND VGND VPWR VPWR _24474_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21686_ _18296_/A VGND VGND VPWR VPWR _21686_/X sky130_fd_sc_hd__buf_2
XFILLER_212_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16762__B1 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23425_ _23425_/CLK _20311_/X VGND VGND VPWR VPWR _22400_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20637_ _20637_/A VGND VGND VPWR VPWR _20637_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19079__A _19074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25540__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23356_ VGND VGND VPWR VPWR _23356_/HI scl_o_S4 sky130_fd_sc_hd__conb_1
XANTENNA__16514__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20568_ _18876_/X _20567_/Y _20553_/C VGND VGND VPWR VPWR _20568_/X sky130_fd_sc_hd__and3_4
XANTENNA__22850__A3 _22849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22307_ _24522_/Q _22807_/A _23001_/A _22306_/X VGND VGND VPWR VPWR _22308_/C sky130_fd_sc_hd__a211o_4
X_23287_ _22286_/X _23277_/X _23287_/C _23286_/X VGND VGND VPWR VPWR _23287_/X sky130_fd_sc_hd__or4_4
X_20499_ _25207_/Q _20497_/X _20477_/C _20498_/X VGND VGND VPWR VPWR _20500_/B sky130_fd_sc_hd__a22oi_4
XFILLER_4_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13040_ _12976_/D _13032_/B VGND VGND VPWR VPWR _13041_/B sky130_fd_sc_hd__or2_4
X_25026_ _25035_/CLK _25026_/D HRESETn VGND VGND VPWR VPWR _25026_/Q sky130_fd_sc_hd__dfrtp_4
X_22238_ _22251_/A _22238_/B VGND VGND VPWR VPWR _22238_/X sky130_fd_sc_hd__or2_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22169_ _22169_/A VGND VGND VPWR VPWR _22174_/B sky130_fd_sc_hd__inv_2
XFILLER_182_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14828__B1 _20664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14991_ _14983_/X _14984_/X _14987_/X _14991_/D VGND VGND VPWR VPWR _15017_/A sky130_fd_sc_hd__or4_4
XFILLER_115_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24493__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13500__B1 _11786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13942_ _13924_/A _15421_/B _13942_/C VGND VGND VPWR VPWR _13957_/A sky130_fd_sc_hd__or3_4
X_16730_ _16730_/A VGND VGND VPWR VPWR _16730_/X sky130_fd_sc_hd__buf_2
XANTENNA__14887__A1_N _25014_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24422__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16661_ _16668_/A VGND VGND VPWR VPWR _16661_/X sky130_fd_sc_hd__buf_2
XFILLER_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13873_ _23967_/Q VGND VGND VPWR VPWR _13873_/X sky130_fd_sc_hd__buf_2
XANTENNA__22118__A2 _22114_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15612_ _24901_/Q VGND VGND VPWR VPWR _15612_/Y sky130_fd_sc_hd__inv_2
X_18400_ _18400_/A VGND VGND VPWR VPWR _18400_/Y sky130_fd_sc_hd__inv_2
X_12824_ _12792_/X _12824_/B _12815_/X _12824_/D VGND VGND VPWR VPWR _12824_/X sky130_fd_sc_hd__or4_4
X_16592_ _16598_/A VGND VGND VPWR VPWR _16592_/X sky130_fd_sc_hd__buf_2
X_19380_ _19372_/A VGND VGND VPWR VPWR _19380_/X sky130_fd_sc_hd__buf_2
XFILLER_62_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15543_ _14366_/A _21290_/A VGND VGND VPWR VPWR _15773_/A sky130_fd_sc_hd__or2_4
X_18331_ _19273_/A _20387_/B _19094_/C VGND VGND VPWR VPWR _19783_/A sky130_fd_sc_hd__or3_4
X_12755_ _12755_/A VGND VGND VPWR VPWR _12755_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _22684_/B VGND VGND VPWR VPWR _11706_/X sky130_fd_sc_hd__buf_2
X_18262_ _24225_/Q VGND VGND VPWR VPWR _23346_/A sky130_fd_sc_hd__inv_2
XFILLER_91_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _14871_/Y _15471_/X _14479_/X _15471_/X VGND VGND VPWR VPWR _15474_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12686_/A _12686_/B _12686_/C VGND VGND VPWR VPWR _12686_/X sky130_fd_sc_hd__and3_4
XANTENNA__16753__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _15457_/A _14425_/B VGND VGND VPWR VPWR _14431_/A sky130_fd_sc_hd__nor2_4
X_17213_ _17213_/A _17210_/X _17211_/X _17213_/D VGND VGND VPWR VPWR _17227_/B sky130_fd_sc_hd__or4_4
XFILLER_202_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18193_ _18193_/A _18193_/B VGND VGND VPWR VPWR _18193_/X sky130_fd_sc_hd__or2_4
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_106_0_HCLK clkbuf_7_53_0_HCLK/X VGND VGND VPWR VPWR _24667_/CLK sky130_fd_sc_hd__clkbuf_1
X_17144_ _17087_/A VGND VGND VPWR VPWR _17148_/C sky130_fd_sc_hd__buf_2
XFILLER_7_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15310__A _15282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _14344_/A _14355_/X _25482_/Q _14349_/X VGND VGND VPWR VPWR _25157_/D sky130_fd_sc_hd__o22a_4
XFILLER_190_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12653__B _12606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_169_0_HCLK clkbuf_7_84_0_HCLK/X VGND VGND VPWR VPWR _23774_/CLK sky130_fd_sc_hd__clkbuf_1
X_13307_ _13227_/X _13307_/B VGND VGND VPWR VPWR _13307_/X sky130_fd_sc_hd__or2_4
X_17075_ _17045_/A _17074_/X VGND VGND VPWR VPWR _17075_/X sky130_fd_sc_hd__or2_4
XFILLER_116_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14287_ _14280_/A _14285_/X _14286_/Y VGND VGND VPWR VPWR _14287_/X sky130_fd_sc_hd__o21a_4
XFILLER_170_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16026_ _16024_/Y _16019_/X _15948_/X _16025_/X VGND VGND VPWR VPWR _16026_/X sky130_fd_sc_hd__a2bb2o_4
X_13238_ _13421_/A VGND VGND VPWR VPWR _13350_/A sky130_fd_sc_hd__buf_2
XFILLER_124_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22143__A _23138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13765__A _13765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13169_ _13169_/A _13169_/B _13169_/C VGND VGND VPWR VPWR _13169_/X sky130_fd_sc_hd__and3_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16141__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17977_ _18113_/A _23785_/Q VGND VGND VPWR VPWR _17981_/B sky130_fd_sc_hd__or2_4
XANTENNA__15492__B1 HADDR[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19716_ _19273_/A _20387_/B _19716_/C _18932_/B VGND VGND VPWR VPWR _19716_/X sky130_fd_sc_hd__or4_4
X_16928_ _16128_/Y _24272_/Q _16128_/Y _24272_/Q VGND VGND VPWR VPWR _16929_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24163__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19647_ _19645_/Y _19641_/X _19646_/X _19641_/A VGND VGND VPWR VPWR _23667_/D sky130_fd_sc_hd__a2bb2o_4
X_16859_ _16858_/X VGND VGND VPWR VPWR _16859_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19578_ _19578_/A VGND VGND VPWR VPWR _19578_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16992__B1 _24721_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18529_ _18468_/A _18526_/X VGND VGND VPWR VPWR _18530_/C sky130_fd_sc_hd__or2_4
XANTENNA__25369__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21540_ _24614_/Q _22130_/B VGND VGND VPWR VPWR _21540_/X sky130_fd_sc_hd__or2_4
XANTENNA__16744__B1 _16391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16961__A1_N _16031_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21471_ _21665_/A _21471_/B VGND VGND VPWR VPWR _21472_/C sky130_fd_sc_hd__or2_4
XFILLER_147_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_65_0_HCLK clkbuf_7_65_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_65_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12844__A _12617_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23210_ _15085_/A _23301_/B VGND VGND VPWR VPWR _23210_/X sky130_fd_sc_hd__or2_4
X_20422_ _20409_/Y VGND VGND VPWR VPWR _20422_/X sky130_fd_sc_hd__buf_2
XFILLER_146_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24190_ _24645_/CLK _24190_/D HRESETn VGND VGND VPWR VPWR _21013_/B sky130_fd_sc_hd__dfrtp_4
X_23141_ _23005_/A _23141_/B _23141_/C VGND VGND VPWR VPWR _23142_/D sky130_fd_sc_hd__and3_4
XFILLER_146_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20353_ _22243_/B _20350_/X _19603_/A _20350_/X VGND VGND VPWR VPWR _23408_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18249__B1 _16601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20284_ _20283_/Y _20279_/X _20008_/X _20266_/Y VGND VGND VPWR VPWR _23434_/D sky130_fd_sc_hd__a2bb2o_4
X_23072_ _23072_/A _23072_/B _23072_/C _23072_/D VGND VGND VPWR VPWR _23072_/X sky130_fd_sc_hd__or4_4
XFILLER_115_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24933__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22023_ _22016_/A _19924_/Y VGND VGND VPWR VPWR _22024_/C sky130_fd_sc_hd__or2_4
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22988__A _16665_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_5_25_0_HCLK_A clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23974_ _23972_/CLK _23972_/Q HRESETn VGND VGND VPWR VPWR _21006_/C sky130_fd_sc_hd__dfstp_4
XFILLER_68_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22925_ _24022_/Q _21292_/X _13636_/D _21315_/X VGND VGND VPWR VPWR _22926_/B sky130_fd_sc_hd__a22oi_4
XFILLER_72_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17224__B2 _21856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11923__A _19620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22856_ _22819_/X _22856_/B _22845_/X _22856_/D VGND VGND VPWR VPWR HRDATA[17] sky130_fd_sc_hd__or4_4
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23034__D _23033_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21807_ _21677_/A _21807_/B VGND VGND VPWR VPWR _21808_/C sky130_fd_sc_hd__or2_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22787_ _22730_/A VGND VGND VPWR VPWR _22921_/B sky130_fd_sc_hd__buf_2
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12540_ _24857_/Q VGND VGND VPWR VPWR _12540_/Y sky130_fd_sc_hd__inv_2
X_24526_ _24555_/CLK _24526_/D HRESETn VGND VGND VPWR VPWR _16591_/A sky130_fd_sc_hd__dfrtp_4
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21738_ _21737_/X VGND VGND VPWR VPWR _21738_/X sky130_fd_sc_hd__buf_2
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15538__B2 _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25039__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22228__A _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21132__A _17438_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12471_ _12208_/X _12468_/X VGND VGND VPWR VPWR _12472_/C sky130_fd_sc_hd__or2_4
X_24457_ _24443_/CLK _24457_/D HRESETn VGND VGND VPWR VPWR _16765_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21669_ _17730_/X VGND VGND VPWR VPWR _21954_/A sky130_fd_sc_hd__buf_2
X_14210_ _14209_/X VGND VGND VPWR VPWR _14212_/A sky130_fd_sc_hd__buf_2
X_23408_ _23441_/CLK _23408_/D VGND VGND VPWR VPWR _20352_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22284__A1 _21077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15190_ _15190_/A VGND VGND VPWR VPWR _15190_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24388_ _24390_/CLK _17112_/X HRESETn VGND VGND VPWR VPWR _24388_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14141_ _14133_/X _14140_/Y _14090_/A _14133_/X VGND VGND VPWR VPWR _25218_/D sky130_fd_sc_hd__a2bb2o_4
X_23339_ _23339_/A _23339_/B VGND VGND VPWR VPWR _23339_/X sky130_fd_sc_hd__or2_4
XFILLER_180_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14072_ _14007_/B _14070_/X _14067_/X _14007_/A _14065_/X VGND VGND VPWR VPWR _25233_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_152_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13023_ _12970_/X _13018_/X _13023_/C VGND VGND VPWR VPWR _13023_/X sky130_fd_sc_hd__and3_4
X_17900_ _17907_/A _17899_/Y VGND VGND VPWR VPWR _17901_/A sky130_fd_sc_hd__and2_4
X_25009_ _25015_/CLK _15279_/X HRESETn VGND VGND VPWR VPWR _25009_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13585__A _14364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22587__A2 _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24674__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18880_ _23946_/Q _18880_/B VGND VGND VPWR VPWR _18881_/B sky130_fd_sc_hd__or2_4
XANTENNA__18255__A3 _15830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24603__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17831_ _17760_/Y _17813_/B _17783_/X _17829_/B VGND VGND VPWR VPWR _17831_/X sky130_fd_sc_hd__a211o_4
XFILLER_86_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20062__A3 _20061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15474__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17762_ _17755_/Y _17756_/Y _17762_/C _17762_/D VGND VGND VPWR VPWR _17763_/B sky130_fd_sc_hd__or4_4
X_14974_ _25036_/Q _14962_/Y _15244_/A _24418_/Q VGND VGND VPWR VPWR _14974_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19501_ _18280_/A _18289_/X _18276_/X _18285_/B VGND VGND VPWR VPWR _19501_/X sky130_fd_sc_hd__or4_4
XFILLER_75_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16713_ _24480_/Q VGND VGND VPWR VPWR _16713_/Y sky130_fd_sc_hd__inv_2
X_13925_ _13925_/A VGND VGND VPWR VPWR _14236_/D sky130_fd_sc_hd__inv_2
XFILLER_35_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17693_ _17575_/Y _17697_/A VGND VGND VPWR VPWR _17695_/A sky130_fd_sc_hd__nand2_4
XFILLER_208_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19432_ _17958_/B VGND VGND VPWR VPWR _19432_/Y sky130_fd_sc_hd__inv_2
X_13856_ _13845_/Y VGND VGND VPWR VPWR _13856_/X sky130_fd_sc_hd__buf_2
X_16644_ _16639_/Y _16643_/X _16373_/X _16643_/X VGND VGND VPWR VPWR _16644_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12807_ _12830_/C VGND VGND VPWR VPWR _12807_/X sky130_fd_sc_hd__buf_2
X_19363_ _19362_/Y _19356_/X _19295_/X _19343_/A VGND VGND VPWR VPWR _23763_/D sky130_fd_sc_hd__a2bb2o_4
X_13787_ _25274_/Q VGND VGND VPWR VPWR _13787_/Y sky130_fd_sc_hd__inv_2
X_16575_ _16574_/Y _16572_/X _16400_/X _16572_/X VGND VGND VPWR VPWR _24533_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18314_ _18314_/A VGND VGND VPWR VPWR _18314_/Y sky130_fd_sc_hd__inv_2
X_12738_ _12879_/A _24810_/Q _12879_/A _24810_/Q VGND VGND VPWR VPWR _12738_/X sky130_fd_sc_hd__a2bb2o_4
X_15526_ _21133_/B VGND VGND VPWR VPWR _15526_/Y sky130_fd_sc_hd__inv_2
X_19294_ _23787_/Q VGND VGND VPWR VPWR _19294_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15529__B2 _15524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22138__A _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15457_ _15457_/A _14212_/B VGND VGND VPWR VPWR _15458_/A sky130_fd_sc_hd__nor2_4
X_18245_ _18236_/A VGND VGND VPWR VPWR _18245_/X sky130_fd_sc_hd__buf_2
X_12669_ _12664_/A _12672_/B VGND VGND VPWR VPWR _12670_/C sky130_fd_sc_hd__nand2_4
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16136__A _16124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ _14408_/A VGND VGND VPWR VPWR _14408_/X sky130_fd_sc_hd__buf_2
XFILLER_163_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15388_ _15294_/B _15400_/B VGND VGND VPWR VPWR _15395_/B sky130_fd_sc_hd__or2_4
X_18176_ _14636_/A _18174_/X _18175_/X VGND VGND VPWR VPWR _18180_/B sky130_fd_sc_hd__and3_4
X_14339_ _14339_/A _14339_/B _14339_/C VGND VGND VPWR VPWR _25163_/D sky130_fd_sc_hd__and3_4
X_17127_ _16991_/Y _17126_/X VGND VGND VPWR VPWR _17127_/X sky130_fd_sc_hd__or2_4
XFILLER_116_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17058_ _17057_/X VGND VGND VPWR VPWR _17058_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16009_ _16009_/A VGND VGND VPWR VPWR _16009_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_7_0_HCLK clkbuf_4_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__24344__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18651__B1 _16566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20971_ _20971_/A _20971_/B VGND VGND VPWR VPWR _24102_/D sky130_fd_sc_hd__and2_4
XANTENNA__20121__A _20116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22710_ _22710_/A _21864_/B _21864_/C VGND VGND VPWR VPWR _22710_/X sky130_fd_sc_hd__and3_4
XANTENNA__11743__A _16236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18954__B2 _18947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23690_ _23706_/CLK _19577_/X VGND VGND VPWR VPWR _23690_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22641_ _16687_/Y _22641_/B VGND VGND VPWR VPWR _22641_/X sky130_fd_sc_hd__and2_4
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25360_ _25387_/CLK _13021_/X HRESETn VGND VGND VPWR VPWR _25360_/Q sky130_fd_sc_hd__dfrtp_4
X_22572_ _21019_/X VGND VGND VPWR VPWR _22572_/X sky130_fd_sc_hd__buf_2
XANTENNA__16717__B1 _16716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21710__B1 _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24311_ _24305_/CLK _17636_/Y HRESETn VGND VGND VPWR VPWR _17543_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_178_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21523_ _21232_/X VGND VGND VPWR VPWR _22522_/B sky130_fd_sc_hd__buf_2
X_25291_ _24236_/CLK _13698_/X HRESETn VGND VGND VPWR VPWR _11826_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24242_ _24889_/CLK _24242_/D HRESETn VGND VGND VPWR VPWR _24242_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21887__A _22056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21454_ _17709_/A VGND VGND VPWR VPWR _21803_/A sky130_fd_sc_hd__buf_2
XFILLER_147_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12754__A1 _25386_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20405_ _13427_/B VGND VGND VPWR VPWR _20405_/Y sky130_fd_sc_hd__inv_2
X_24173_ _24172_/CLK _24173_/D HRESETn VGND VGND VPWR VPWR _24173_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19357__A _11785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21385_ _21239_/A VGND VGND VPWR VPWR _21385_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_152_0_HCLK clkbuf_7_76_0_HCLK/X VGND VGND VPWR VPWR _25308_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23124_ _22684_/B VGND VGND VPWR VPWR _23292_/B sky130_fd_sc_hd__buf_2
XFILLER_190_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20336_ _23414_/Q VGND VGND VPWR VPWR _20336_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23215__B1 _23203_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11918__A _19617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23055_ _17234_/Y _22916_/X _12796_/A _22917_/X VGND VGND VPWR VPWR _23055_/X sky130_fd_sc_hd__a2bb2o_4
X_20267_ _20266_/Y VGND VGND VPWR VPWR _20267_/X sky130_fd_sc_hd__buf_2
XANTENNA__24085__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22006_ _24231_/Q _22735_/B _21511_/X _22005_/Y VGND VGND VPWR VPWR _22006_/X sky130_fd_sc_hd__a211o_4
XFILLER_1_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20198_ _17952_/B VGND VGND VPWR VPWR _20198_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24014__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21529__B1 _24857_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16853__A1_N _16852_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11971_ _11967_/A _11932_/B _11970_/Y VGND VGND VPWR VPWR _11971_/Y sky130_fd_sc_hd__a21oi_4
X_23957_ _23958_/CLK _23957_/D HRESETn VGND VGND VPWR VPWR _23957_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12749__A _21027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13710_ _11823_/Y _13672_/B VGND VGND VPWR VPWR _13710_/Y sky130_fd_sc_hd__nand2_4
XFILLER_72_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22908_ _22136_/B VGND VGND VPWR VPWR _22908_/X sky130_fd_sc_hd__buf_2
XFILLER_205_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14690_ _21764_/A _14685_/Y _21757_/A _14684_/X VGND VGND VPWR VPWR _14704_/A sky130_fd_sc_hd__o22a_4
XFILLER_205_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23888_ _23887_/CLK _23888_/D VGND VGND VPWR VPWR _18045_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__16956__B1 _15980_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13641_ _13640_/X VGND VGND VPWR VPWR _13641_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22839_ _22928_/A VGND VGND VPWR VPWR _22839_/X sky130_fd_sc_hd__buf_2
XFILLER_32_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16360_ _24612_/Q VGND VGND VPWR VPWR _16360_/Y sky130_fd_sc_hd__inv_2
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _25256_/Q _14549_/A _25255_/Q _14549_/B VGND VGND VPWR VPWR _13574_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15311_ _15323_/A _15311_/B VGND VGND VPWR VPWR _15320_/D sky130_fd_sc_hd__and2_4
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _25409_/Q VGND VGND VPWR VPWR _12704_/A sky130_fd_sc_hd__inv_2
X_24509_ _24032_/CLK _16644_/X HRESETn VGND VGND VPWR VPWR _16639_/A sky130_fd_sc_hd__dfrtp_4
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16291_ _16291_/A VGND VGND VPWR VPWR _16291_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25489_ _25466_/CLK _25489_/D HRESETn VGND VGND VPWR VPWR _12029_/A sky130_fd_sc_hd__dfrtp_4
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15242_ _14903_/X _15242_/B VGND VGND VPWR VPWR _15243_/B sky130_fd_sc_hd__or2_4
X_18030_ _18030_/A _18030_/B _18030_/C VGND VGND VPWR VPWR _18035_/B sky130_fd_sc_hd__and3_4
XANTENNA__14195__B1 _13829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12454_ _12454_/A VGND VGND VPWR VPWR _25445_/D sky130_fd_sc_hd__inv_2
XANTENNA__24855__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15173_ _15173_/A VGND VGND VPWR VPWR _15173_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20807__A2 _20708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12745__B2 _24811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12385_ _12264_/Y _12385_/B VGND VGND VPWR VPWR _12385_/X sky130_fd_sc_hd__or2_4
XANTENNA__17133__B1 _17053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14124_ _14092_/A _14092_/B _14092_/A _14092_/B VGND VGND VPWR VPWR _14124_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22405__B _21064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19981_ _19981_/A VGND VGND VPWR VPWR _19981_/X sky130_fd_sc_hd__buf_2
XFILLER_153_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14055_ _14049_/B VGND VGND VPWR VPWR _14055_/X sky130_fd_sc_hd__buf_2
X_18932_ _19716_/C _18932_/B _20387_/A _20387_/B VGND VGND VPWR VPWR _18932_/X sky130_fd_sc_hd__or4_4
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13006_ _13000_/A _13005_/X _12998_/A _13001_/Y VGND VGND VPWR VPWR _13007_/A sky130_fd_sc_hd__a211o_4
XFILLER_140_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18863_ _16450_/Y _18703_/A _16450_/Y _18703_/A VGND VGND VPWR VPWR _18866_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17814_ _16938_/Y _17814_/B VGND VGND VPWR VPWR _17817_/B sky130_fd_sc_hd__or2_4
XFILLER_223_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18794_ _18789_/A _18797_/A _18797_/B VGND VGND VPWR VPWR _18794_/X sky130_fd_sc_hd__or3_4
XFILLER_239_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21037__A _24785_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17745_ _24283_/Q VGND VGND VPWR VPWR _17746_/A sky130_fd_sc_hd__inv_2
X_14957_ _15229_/A _24429_/Q _15061_/A _24429_/Q VGND VGND VPWR VPWR _14957_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11776__A1_N _11772_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13908_ _13908_/A VGND VGND VPWR VPWR _13931_/A sky130_fd_sc_hd__buf_2
X_17676_ _17682_/A _17676_/B _17676_/C VGND VGND VPWR VPWR _17676_/X sky130_fd_sc_hd__and3_4
XFILLER_223_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14888_ _25033_/Q VGND VGND VPWR VPWR _14888_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19415_ _19410_/Y _19413_/X _19414_/X _19413_/X VGND VGND VPWR VPWR _23746_/D sky130_fd_sc_hd__a2bb2o_4
X_16627_ _13728_/B VGND VGND VPWR VPWR _16631_/A sky130_fd_sc_hd__inv_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17458__A2_N _13157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13839_ _13839_/A VGND VGND VPWR VPWR _13840_/C sky130_fd_sc_hd__inv_2
XFILLER_211_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18346__A _13157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19346_ _19345_/Y _19343_/X _19279_/X _19343_/X VGND VGND VPWR VPWR _19346_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22496__A1 _11681_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16558_ _16557_/Y _16555_/X _16295_/X _16555_/X VGND VGND VPWR VPWR _24540_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15509_ _15508_/Y _15506_/X HADDR[13] _15506_/X VGND VGND VPWR VPWR _15509_/X sky130_fd_sc_hd__a2bb2o_4
X_19277_ _19272_/Y _19276_/X _19144_/X _19276_/X VGND VGND VPWR VPWR _19277_/X sky130_fd_sc_hd__a2bb2o_4
X_16489_ _16487_/Y _16482_/X _16397_/X _16488_/X VGND VGND VPWR VPWR _24566_/D sky130_fd_sc_hd__a2bb2o_4
X_18228_ _18132_/A _18220_/X _18228_/C VGND VGND VPWR VPWR _18228_/X sky130_fd_sc_hd__and3_4
XFILLER_164_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24596__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18159_ _18094_/A _18159_/B _18159_/C VGND VGND VPWR VPWR _18163_/B sky130_fd_sc_hd__and3_4
XFILLER_144_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23288__A2_N _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24525__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21170_ _16852_/Y _21519_/A VGND VGND VPWR VPWR _21170_/X sky130_fd_sc_hd__or2_4
XFILLER_172_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_225_0_HCLK clkbuf_7_112_0_HCLK/X VGND VGND VPWR VPWR _24976_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12841__B _12804_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20116__A _20116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20121_ _20116_/A VGND VGND VPWR VPWR _20121_/X sky130_fd_sc_hd__buf_2
XANTENNA__11738__A HWDATA[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19905__A _19900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20052_ _20052_/A VGND VGND VPWR VPWR _20054_/A sky130_fd_sc_hd__buf_2
XFILLER_219_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24860_ _25403_/CLK _15760_/X HRESETn VGND VGND VPWR VPWR _12551_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22050__B _23342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23811_ _23873_/CLK _19229_/X VGND VGND VPWR VPWR _23811_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24791_ _24795_/CLK _15895_/X HRESETn VGND VGND VPWR VPWR _22295_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22184__B1 _17417_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25384__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23742_ _25073_/CLK _23742_/D VGND VGND VPWR VPWR _18111_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_199_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ _20952_/Y _20949_/X _20953_/X VGND VGND VPWR VPWR _20954_/X sky130_fd_sc_hd__o21a_4
XFILLER_214_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _25326_/CLK _19631_/X VGND VGND VPWR VPWR _13228_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _20883_/Y _20880_/Y _20888_/A VGND VGND VPWR VPWR _20885_/X sky130_fd_sc_hd__o21a_4
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25412_ _24032_/CLK _25412_/D HRESETn VGND VGND VPWR VPWR _25412_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_241_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22624_ _22521_/B _22621_/X _22423_/X _22623_/X VGND VGND VPWR VPWR _22624_/X sky130_fd_sc_hd__o22a_4
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25343_ _25344_/CLK _13083_/X HRESETn VGND VGND VPWR VPWR _12305_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_166_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22555_ _22554_/X VGND VGND VPWR VPWR _22555_/X sky130_fd_sc_hd__buf_2
XFILLER_10_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21506_ _21379_/B _21505_/X VGND VGND VPWR VPWR _21507_/C sky130_fd_sc_hd__or2_4
X_25274_ _25325_/CLK _13789_/X HRESETn VGND VGND VPWR VPWR _25274_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22486_ _21864_/B VGND VGND VPWR VPWR _22486_/X sky130_fd_sc_hd__buf_2
XFILLER_155_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_35_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24225_ _24227_/CLK _24225_/D HRESETn VGND VGND VPWR VPWR _24225_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21437_ _21232_/X VGND VGND VPWR VPWR _21437_/X sky130_fd_sc_hd__buf_2
XFILLER_135_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24266__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12170_ _12170_/A VGND VGND VPWR VPWR _12279_/A sky130_fd_sc_hd__inv_2
X_24156_ _24080_/CLK _18711_/Y HRESETn VGND VGND VPWR VPWR _24156_/Q sky130_fd_sc_hd__dfrtp_4
X_21368_ _21368_/A VGND VGND VPWR VPWR _21722_/B sky130_fd_sc_hd__buf_2
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23107_ _23280_/A _23107_/B VGND VGND VPWR VPWR _23115_/C sky130_fd_sc_hd__and2_4
XFILLER_1_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20319_ _20306_/X _19573_/X _18257_/X _20318_/X _20310_/X VGND VGND VPWR VPWR _23421_/D
+ sky130_fd_sc_hd__a32o_4
X_24087_ _25226_/CLK _20470_/X HRESETn VGND VGND VPWR VPWR _20445_/A sky130_fd_sc_hd__dfrtp_4
X_21299_ _21298_/X VGND VGND VPWR VPWR _21300_/A sky130_fd_sc_hd__buf_2
XFILLER_1_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23038_ _23035_/X _23036_/X _22858_/X _24843_/Q _23037_/X VGND VGND VPWR VPWR _23038_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_110_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22411__B2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22962__A2 _22960_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15860_ _15881_/A VGND VGND VPWR VPWR _15889_/A sky130_fd_sc_hd__inv_2
X_14811_ _14811_/A _14811_/B _25051_/Q VGND VGND VPWR VPWR _14811_/X sky130_fd_sc_hd__or3_4
XFILLER_91_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15791_ _15811_/A VGND VGND VPWR VPWR _15820_/A sky130_fd_sc_hd__inv_2
X_24989_ _24976_/CLK _24989_/D HRESETn VGND VGND VPWR VPWR _24989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22175__B1 _25439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17530_ _17530_/A VGND VGND VPWR VPWR _17530_/Y sky130_fd_sc_hd__inv_2
X_11954_ _11938_/A _11938_/B _11929_/X VGND VGND VPWR VPWR _11954_/X sky130_fd_sc_hd__and3_4
X_14742_ _14711_/X _14741_/X _14711_/X _14741_/X VGND VGND VPWR VPWR _25064_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25054__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14673_ _14673_/A VGND VGND VPWR VPWR _14741_/A sky130_fd_sc_hd__inv_2
X_17461_ _20387_/B VGND VGND VPWR VPWR _18911_/B sky130_fd_sc_hd__buf_2
X_11885_ _11797_/A _11856_/X _11883_/Y _25514_/Q _11884_/Y VGND VGND VPWR VPWR _11885_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_233_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14694__A _22213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19200_ _19063_/A VGND VGND VPWR VPWR _19200_/X sky130_fd_sc_hd__buf_2
XFILLER_32_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13624_ _13623_/X VGND VGND VPWR VPWR _13625_/A sky130_fd_sc_hd__inv_2
X_16412_ _16410_/Y _16406_/X _16229_/X _16411_/X VGND VGND VPWR VPWR _24594_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_117_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_234_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17392_ _17392_/A _17392_/B VGND VGND VPWR VPWR _17393_/B sky130_fd_sc_hd__or2_4
XFILLER_220_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19131_ _19130_/Y _19126_/X _19106_/X _19126_/X VGND VGND VPWR VPWR _23846_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13555_ _13555_/A VGND VGND VPWR VPWR _14563_/C sky130_fd_sc_hd__buf_2
X_16343_ _24618_/Q VGND VGND VPWR VPWR _16343_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12506_ _12505_/Y _24880_/Q _12505_/Y _24880_/Q VGND VGND VPWR VPWR _12506_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16274_ _15665_/X _15986_/Y _16267_/X _24644_/Q _16273_/X VGND VGND VPWR VPWR _16274_/X
+ sky130_fd_sc_hd__a32o_4
X_19062_ _19054_/A VGND VGND VPWR VPWR _19062_/X sky130_fd_sc_hd__buf_2
XFILLER_173_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ _12009_/Y _13485_/X _11753_/X _13485_/X VGND VGND VPWR VPWR _13486_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15225_ _15225_/A VGND VGND VPWR VPWR _25024_/D sky130_fd_sc_hd__inv_2
X_18013_ _18017_/A VGND VGND VPWR VPWR _18014_/A sky130_fd_sc_hd__buf_2
X_12437_ _12434_/A _12433_/B _12437_/C VGND VGND VPWR VPWR _12437_/X sky130_fd_sc_hd__and3_4
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12942__A _12772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15156_ _15149_/X _15156_/B _15156_/C _15155_/X VGND VGND VPWR VPWR _15156_/X sky130_fd_sc_hd__or4_4
X_12368_ _12368_/A _12363_/X _12364_/X _12368_/D VGND VGND VPWR VPWR _12368_/X sky130_fd_sc_hd__or4_4
XFILLER_99_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14107_ _14106_/X VGND VGND VPWR VPWR _14108_/B sky130_fd_sc_hd__inv_2
XFILLER_113_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15087_ _15087_/A VGND VGND VPWR VPWR _15087_/Y sky130_fd_sc_hd__inv_2
X_19964_ _19964_/A VGND VGND VPWR VPWR _19964_/X sky130_fd_sc_hd__buf_2
X_12299_ _12299_/A VGND VGND VPWR VPWR _12983_/D sky130_fd_sc_hd__inv_2
XFILLER_234_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22938__C1 _22937_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14038_ _13995_/A _14038_/B _13989_/X _14038_/D VGND VGND VPWR VPWR _14038_/X sky130_fd_sc_hd__and4_4
X_18915_ _23921_/Q VGND VGND VPWR VPWR _18915_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23989__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19895_ _19895_/A VGND VGND VPWR VPWR _21184_/B sky130_fd_sc_hd__inv_2
Xclkbuf_8_55_0_HCLK clkbuf_8_55_0_HCLK/A VGND VGND VPWR VPWR _24357_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_110_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18846_ _18830_/X _18835_/X _18840_/X _18845_/X VGND VGND VPWR VPWR _18846_/X sky130_fd_sc_hd__or4_4
XFILLER_110_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16093__B1 _15996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21990__A _21841_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18777_ _24139_/Q _18777_/B VGND VGND VPWR VPWR _18779_/B sky130_fd_sc_hd__or2_4
XANTENNA__24955__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15989_ _15988_/X VGND VGND VPWR VPWR _15990_/A sky130_fd_sc_hd__buf_2
XFILLER_209_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17728_ _18279_/A _17726_/B _17727_/Y VGND VGND VPWR VPWR _17728_/X sky130_fd_sc_hd__o21a_4
XFILLER_82_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19031__B1 _18981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17659_ _17659_/A _17659_/B VGND VGND VPWR VPWR _17661_/B sky130_fd_sc_hd__or2_4
X_20670_ _20670_/A VGND VGND VPWR VPWR _20670_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24777__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19329_ _23775_/Q VGND VGND VPWR VPWR _19329_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24706__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22340_ _21926_/A _22340_/B VGND VGND VPWR VPWR _22341_/C sky130_fd_sc_hd__or2_4
XFILLER_148_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22271_ _21284_/X _22233_/X _21956_/X _22270_/X VGND VGND VPWR VPWR _22271_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12852__A _12769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24010_ _24900_/CLK _24010_/D HRESETn VGND VGND VPWR VPWR _13117_/A sky130_fd_sc_hd__dfrtp_4
X_21222_ _21222_/A VGND VGND VPWR VPWR _21222_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21153_ _21149_/X _21152_/X VGND VGND VPWR VPWR _21153_/X sky130_fd_sc_hd__and2_4
XFILLER_171_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20104_ _23501_/Q VGND VGND VPWR VPWR _21618_/B sky130_fd_sc_hd__inv_2
X_21084_ _22840_/A VGND VGND VPWR VPWR _22451_/A sky130_fd_sc_hd__buf_2
XFILLER_247_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20404__B1 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14882__B2 _24425_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20035_ _20031_/Y _20034_/X _19807_/X _20034_/X VGND VGND VPWR VPWR _20035_/X sky130_fd_sc_hd__a2bb2o_4
X_24912_ _24032_/CLK _24912_/D HRESETn VGND VGND VPWR VPWR _24912_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22996__A _22996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24843_ _25390_/CLK _15801_/X HRESETn VGND VGND VPWR VPWR _24843_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15831__B1 _24824_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24774_ _25380_/CLK _24774_/D HRESETn VGND VGND VPWR VPWR _23144_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ _21281_/B _21973_/X _21977_/Y _21511_/X _21985_/X VGND VGND VPWR VPWR _21986_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_233_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _23427_/CLK _19471_/X VGND VGND VPWR VPWR _19469_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_215_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20937_ _20935_/Y _20932_/Y _20941_/B VGND VGND VPWR VPWR _20937_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17602__B _17602_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11670_/A _15496_/A _15518_/A VGND VGND VPWR VPWR _15640_/B sky130_fd_sc_hd__or3_4
X_23656_ _23665_/CLK _23656_/D VGND VGND VPWR VPWR _13266_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _16694_/Y _20846_/X _20855_/X _20867_/X VGND VGND VPWR VPWR _20868_/X sky130_fd_sc_hd__o22a_4
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22607_ _22758_/A _22607_/B VGND VGND VPWR VPWR _22607_/Y sky130_fd_sc_hd__nor2_4
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14664__D _21283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23587_ _23555_/CLK _23587_/D VGND VGND VPWR VPWR _23587_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20799_ _20780_/X _20798_/X _24918_/Q _20784_/X VGND VGND VPWR VPWR _20799_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24447__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13340_ _13443_/A _13340_/B VGND VGND VPWR VPWR _13341_/C sky130_fd_sc_hd__or2_4
X_25326_ _25326_/CLK _25326_/D HRESETn VGND VGND VPWR VPWR _25326_/Q sky130_fd_sc_hd__dfrtp_4
X_22538_ _24424_/Q _21031_/X _22533_/X _22537_/X VGND VGND VPWR VPWR _22539_/C sky130_fd_sc_hd__a211o_4
XFILLER_155_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15898__B1 _24789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13271_ _13268_/X _13271_/B _13270_/X VGND VGND VPWR VPWR _13271_/X sky130_fd_sc_hd__and3_4
X_25257_ _25325_/CLK _13834_/X HRESETn VGND VGND VPWR VPWR _13552_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_127_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22469_ _22290_/X VGND VGND VPWR VPWR _22469_/X sky130_fd_sc_hd__buf_2
X_15010_ _24473_/Q VGND VGND VPWR VPWR _15010_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18849__A1_N _16527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12222_ _25445_/Q VGND VGND VPWR VPWR _12275_/B sky130_fd_sc_hd__inv_2
X_24208_ _24208_/CLK _18338_/X HRESETn VGND VGND VPWR VPWR _24208_/Q sky130_fd_sc_hd__dfrtp_4
X_25188_ _25249_/CLK _14257_/X HRESETn VGND VGND VPWR VPWR _14256_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13577__B _13577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12153_ _14339_/A VGND VGND VPWR VPWR _12153_/Y sky130_fd_sc_hd__inv_2
X_24139_ _24139_/CLK _18779_/X HRESETn VGND VGND VPWR VPWR _24139_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12084_ _12084_/A VGND VGND VPWR VPWR _21570_/A sky130_fd_sc_hd__buf_2
X_16961_ _16031_/Y _17027_/A _16031_/Y _17027_/A VGND VGND VPWR VPWR _16968_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18700_ _18707_/A _18707_/B _18700_/C _18699_/X VGND VGND VPWR VPWR _18700_/X sky130_fd_sc_hd__or4_4
X_15912_ _15678_/X _15694_/X _15906_/X _15911_/X VGND VGND VPWR VPWR _15912_/X sky130_fd_sc_hd__a211o_4
X_19680_ _13304_/B VGND VGND VPWR VPWR _19680_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12811__A2_N _24811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16892_ _16887_/X _16892_/B _16890_/X _16891_/X VGND VGND VPWR VPWR _16892_/X sky130_fd_sc_hd__or4_4
XFILLER_238_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20946__A1 _16650_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18631_ _24544_/Q _24155_/Q _16546_/Y _18707_/A VGND VGND VPWR VPWR _18637_/B sky130_fd_sc_hd__o22a_4
X_15843_ _15700_/X VGND VGND VPWR VPWR _15843_/X sky130_fd_sc_hd__buf_2
XFILLER_237_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22148__B1 _22525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15822__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18562_ _18562_/A _18562_/B VGND VGND VPWR VPWR _18563_/B sky130_fd_sc_hd__or2_4
X_12986_ _12978_/X _12985_/X VGND VGND VPWR VPWR _12986_/X sky130_fd_sc_hd__or2_4
X_15774_ _15544_/Y _15651_/X _15770_/X _20684_/A _15773_/X VGND VGND VPWR VPWR _15774_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22699__B2 _22698_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17513_ _17513_/A VGND VGND VPWR VPWR _17513_/Y sky130_fd_sc_hd__inv_2
X_14725_ _14722_/Y _14702_/X _14724_/Y VGND VGND VPWR VPWR _14725_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21315__A _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11937_ _17442_/B VGND VGND VPWR VPWR _11938_/B sky130_fd_sc_hd__inv_2
X_18493_ _18493_/A _18493_/B VGND VGND VPWR VPWR _18496_/B sky130_fd_sc_hd__or2_4
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21371__B2 _21721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17444_ _13584_/X VGND VGND VPWR VPWR _21177_/A sky130_fd_sc_hd__buf_2
X_11868_ _11797_/Y VGND VGND VPWR VPWR _11869_/A sky130_fd_sc_hd__buf_2
X_14656_ _25073_/Q _19026_/C _14784_/A VGND VGND VPWR VPWR _14656_/X sky130_fd_sc_hd__o21a_4
XFILLER_220_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24870__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ _14647_/B VGND VGND VPWR VPWR _14650_/A sky130_fd_sc_hd__inv_2
XPHY_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17375_ _17241_/Y _17374_/X _17268_/X VGND VGND VPWR VPWR _17375_/Y sky130_fd_sc_hd__a21oi_4
X_11799_ _11799_/A VGND VGND VPWR VPWR _11799_/X sky130_fd_sc_hd__buf_2
X_14587_ _14554_/A _14554_/B VGND VGND VPWR VPWR _14587_/Y sky130_fd_sc_hd__nand2_4
XFILLER_229_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19114_ _19113_/Y _19109_/X _18998_/X _19101_/A VGND VGND VPWR VPWR _23851_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24188__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16326_ _16324_/Y _16319_/X _16229_/X _16325_/X VGND VGND VPWR VPWR _16326_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13538_ _13538_/A VGND VGND VPWR VPWR _13538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22871__A1 _11681_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15138__A2_N _24602_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24117__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19045_ _19044_/Y _19040_/X _18998_/X _19028_/A VGND VGND VPWR VPWR _23875_/D sky130_fd_sc_hd__a2bb2o_4
X_13469_ _13464_/A VGND VGND VPWR VPWR _13469_/X sky130_fd_sc_hd__buf_2
X_16257_ _16183_/Y VGND VGND VPWR VPWR _16257_/X sky130_fd_sc_hd__buf_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15208_ _15207_/X VGND VGND VPWR VPWR _15209_/B sky130_fd_sc_hd__inv_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18827__B1 _16498_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16188_ _16187_/Y _16185_/X _15554_/X _16185_/X VGND VGND VPWR VPWR _16188_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15983__A _23138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15139_ _24980_/Q VGND VGND VPWR VPWR _15139_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19947_ _19945_/Y _19941_/X _19606_/X _19946_/X VGND VGND VPWR VPWR _19947_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15656__A3 _15643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22312__C _22311_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19878_ _19878_/A VGND VGND VPWR VPWR _19878_/Y sky130_fd_sc_hd__inv_2
XFILLER_228_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16066__B1 _15466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17802__A1 _16906_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18829_ _16463_/Y _24154_/Q _16463_/Y _24154_/Q VGND VGND VPWR VPWR _18830_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21840_ _21122_/X _21834_/Y _21556_/A _21839_/X VGND VGND VPWR VPWR _21840_/X sky130_fd_sc_hd__o22a_4
XANTENNA__17703__A _13807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23351__A2 _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22154__A3 _21427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21771_ _21771_/A _20168_/Y VGND VGND VPWR VPWR _21772_/C sky130_fd_sc_hd__or2_4
XANTENNA__12847__A _25399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23510_ _23526_/CLK _23510_/D VGND VGND VPWR VPWR _23510_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20722_ _20722_/A VGND VGND VPWR VPWR _20723_/A sky130_fd_sc_hd__inv_2
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14765__C _13577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24490_ _24487_/CLK _16690_/X HRESETn VGND VGND VPWR VPWR _16689_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_224_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23441_ _23441_/CLK _23441_/D VGND VGND VPWR VPWR _20264_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20653_ _17393_/B _20652_/Y _20661_/C VGND VGND VPWR VPWR _20653_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_100_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_201_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14977__A2_N _14885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24540__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23372_ _23932_/CLK scl_oen_o_S4 VGND VGND VPWR VPWR _23372_/Q sky130_fd_sc_hd__dfxtp_4
X_20584_ _23946_/Q _18880_/B VGND VGND VPWR VPWR _20584_/Y sky130_fd_sc_hd__nand2_4
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22056__A _22056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25111_ _23958_/CLK _14498_/X HRESETn VGND VGND VPWR VPWR _25111_/Q sky130_fd_sc_hd__dfrtp_4
X_22323_ _11976_/Y _21570_/A _11975_/Y _12057_/A VGND VGND VPWR VPWR _22323_/X sky130_fd_sc_hd__o22a_4
XFILLER_164_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16054__A _24723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25042_ _25043_/CLK _14874_/Y HRESETn VGND VGND VPWR VPWR _14859_/B sky130_fd_sc_hd__dfrtp_4
X_22254_ _22261_/A _19943_/Y VGND VGND VPWR VPWR _22256_/B sky130_fd_sc_hd__or2_4
XFILLER_118_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21205_ _21205_/A _20345_/Y VGND VGND VPWR VPWR _21207_/B sky130_fd_sc_hd__or2_4
X_22185_ _22184_/X VGND VGND VPWR VPWR _22185_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22503__B _22505_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21136_ _14388_/Y _14182_/A _14459_/Y _21368_/A VGND VGND VPWR VPWR _21141_/B sky130_fd_sc_hd__o22a_4
XANTENNA__15647__A3 _15643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21067_ _24714_/Q _15649_/Y _21042_/X _21066_/X VGND VGND VPWR VPWR _21068_/A sky130_fd_sc_hd__a211o_4
XFILLER_247_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21050__B1 _21047_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20018_ _20012_/Y VGND VGND VPWR VPWR _20018_/X sky130_fd_sc_hd__buf_2
XFILLER_235_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15804__B1 _15581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12840_ _12835_/X _12839_/X VGND VGND VPWR VPWR _12841_/D sky130_fd_sc_hd__or2_4
X_24826_ _25428_/CLK _24826_/D HRESETn VGND VGND VPWR VPWR _24826_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24699__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12771_ _25397_/Q _12770_/A _12769_/Y _12770_/Y VGND VGND VPWR VPWR _12771_/X sky130_fd_sc_hd__o22a_4
X_21969_ _23690_/Q _19578_/A _19580_/A _21969_/D VGND VGND VPWR VPWR _21969_/X sky130_fd_sc_hd__or4_4
X_24757_ _25369_/CLK _15967_/X HRESETn VGND VGND VPWR VPWR _22476_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16229__A _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11682_/Y VGND VGND VPWR VPWR _11766_/A sky130_fd_sc_hd__buf_2
X_14510_ _23957_/Q VGND VGND VPWR VPWR _14510_/X sky130_fd_sc_hd__buf_2
XANTENNA__24628__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _14177_/B _15486_/X HADDR[22] _15489_/X VGND VGND VPWR VPWR _15490_/X sky130_fd_sc_hd__a2bb2o_4
X_23708_ _23691_/CLK _19518_/X VGND VGND VPWR VPWR _19517_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_42_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24688_ _24744_/CLK _24688_/D HRESETn VGND VGND VPWR VPWR _22405_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15032__B2 _24453_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11651_/Y _17703_/B VGND VGND VPWR VPWR _14364_/A sky130_fd_sc_hd__or2_4
X_14441_ _14096_/A VGND VGND VPWR VPWR _20600_/A sky130_fd_sc_hd__buf_2
X_23639_ _23627_/CLK _23639_/D VGND VGND VPWR VPWR _19725_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_187_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13043__B1 _13019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22302__B1 _22301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24281__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14372_ _14370_/Y VGND VGND VPWR VPWR _14372_/X sky130_fd_sc_hd__buf_2
X_17160_ _17151_/X _17159_/X _17148_/C VGND VGND VPWR VPWR _24374_/D sky130_fd_sc_hd__and3_4
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24210__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13323_ _13189_/A VGND VGND VPWR VPWR _13388_/A sky130_fd_sc_hd__buf_2
X_16111_ _16111_/A VGND VGND VPWR VPWR _16111_/X sky130_fd_sc_hd__buf_2
XANTENNA__20864__B1 _20855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25309_ _25466_/CLK _25309_/D HRESETn VGND VGND VPWR VPWR _13498_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17091_ _17091_/A VGND VGND VPWR VPWR _17091_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21301__C _21306_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13254_ _13254_/A _13254_/B _13253_/X VGND VGND VPWR VPWR _13255_/C sky130_fd_sc_hd__and3_4
X_16042_ _16042_/A VGND VGND VPWR VPWR _16042_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15886__A3 _16236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25487__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12205_ _12205_/A VGND VGND VPWR VPWR _12205_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19275__A _19274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13185_ _13164_/X _13181_/X _13184_/A _25333_/Q _13186_/A VGND VGND VPWR VPWR _25333_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19801_ _19800_/Y _19796_/X _19759_/X _19784_/A VGND VGND VPWR VPWR _23611_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16296__B1 _16295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12136_ _12135_/X VGND VGND VPWR VPWR _12136_/Y sky130_fd_sc_hd__inv_2
X_17993_ _18054_/A VGND VGND VPWR VPWR _18151_/A sky130_fd_sc_hd__buf_2
XFILLER_215_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12750__A2_N _24785_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19732_ _19730_/Y _19731_/X _19708_/X _19731_/X VGND VGND VPWR VPWR _23637_/D sky130_fd_sc_hd__a2bb2o_4
X_12067_ _25483_/Q VGND VGND VPWR VPWR _12067_/Y sky130_fd_sc_hd__inv_2
X_16944_ _16088_/Y _24288_/Q _16088_/Y _24288_/Q VGND VGND VPWR VPWR _16944_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14212__A _14212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23030__B2 _21051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16048__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19663_ _13371_/B VGND VGND VPWR VPWR _19663_/Y sky130_fd_sc_hd__inv_2
X_16875_ _16875_/A VGND VGND VPWR VPWR _19824_/A sky130_fd_sc_hd__buf_2
X_18614_ _24153_/Q VGND VGND VPWR VPWR _18698_/A sky130_fd_sc_hd__inv_2
XFILLER_231_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_129_0_HCLK clkbuf_7_64_0_HCLK/X VGND VGND VPWR VPWR _25326_/CLK sky130_fd_sc_hd__clkbuf_1
X_15826_ _12284_/Y _15823_/X _15619_/X _15823_/X VGND VGND VPWR VPWR _24826_/D sky130_fd_sc_hd__a2bb2o_4
X_19594_ _19594_/A VGND VGND VPWR VPWR _19594_/Y sky130_fd_sc_hd__inv_2
X_18545_ _18523_/X _18538_/X _18545_/C VGND VGND VPWR VPWR _18545_/X sky130_fd_sc_hd__and3_4
X_15757_ _12530_/Y _15755_/X _15616_/X _15755_/X VGND VGND VPWR VPWR _24862_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17242__B _17242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12969_ _21016_/A _12854_/X _12968_/Y VGND VGND VPWR VPWR _12969_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17548__B1 _25521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24369__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14708_ _14707_/X _13748_/Y _14707_/X _13748_/Y VGND VGND VPWR VPWR _14708_/X sky130_fd_sc_hd__a2bb2o_4
X_18476_ _24158_/Q VGND VGND VPWR VPWR _18477_/D sky130_fd_sc_hd__inv_2
X_15688_ _15688_/A _15681_/A VGND VGND VPWR VPWR _18022_/A sky130_fd_sc_hd__or2_4
XANTENNA__16220__B1 _15953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17427_ _21722_/A _17422_/X _16783_/X _17422_/X VGND VGND VPWR VPWR _24329_/D sky130_fd_sc_hd__a2bb2o_4
X_14639_ _14639_/A VGND VGND VPWR VPWR _18017_/A sky130_fd_sc_hd__buf_2
XFILLER_159_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17358_ _17358_/A _17358_/B VGND VGND VPWR VPWR _17359_/C sky130_fd_sc_hd__or2_4
XANTENNA__15697__B _15697_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16309_ _16308_/Y _16306_/X _15946_/X _16306_/X VGND VGND VPWR VPWR _24632_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17289_ _17234_/Y _17288_/X VGND VGND VPWR VPWR _17299_/B sky130_fd_sc_hd__or2_4
XFILLER_162_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19028_ _19028_/A VGND VGND VPWR VPWR _19028_/X sky130_fd_sc_hd__buf_2
XFILLER_162_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11746__A _25531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19225__B1 _19200_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23990_ _24340_/CLK _23989_/Q HRESETn VGND VGND VPWR VPWR _23990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16039__B1 _11735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_25_0_HCLK clkbuf_7_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22941_ _16569_/A _22730_/X _15663_/X _22940_/X VGND VGND VPWR VPWR _22941_/X sky130_fd_sc_hd__a211o_4
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_88_0_HCLK clkbuf_7_89_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_88_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22780__B1 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22872_ _22774_/X _22867_/Y _22868_/X _22871_/X VGND VGND VPWR VPWR _22873_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21823_ _23421_/Q _20307_/X _23397_/Q _21960_/B VGND VGND VPWR VPWR _21823_/X sky130_fd_sc_hd__o22a_4
X_24611_ _24597_/CLK _16371_/X HRESETn VGND VGND VPWR VPWR _16363_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_83_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24792__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15801__A3 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16049__A _24725_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24721__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24542_ _24574_/CLK _16553_/X HRESETn VGND VGND VPWR VPWR _24542_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21754_ _21769_/A _21754_/B _21753_/X VGND VGND VPWR VPWR _21754_/X sky130_fd_sc_hd__and3_4
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16211__B1 _16020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24039__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20705_ _13114_/A _13113_/X _20704_/Y VGND VGND VPWR VPWR _20705_/Y sky130_fd_sc_hd__a21oi_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24473_ _24443_/CLK _24473_/D HRESETn VGND VGND VPWR VPWR _24473_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_196_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21685_ _21803_/A _21685_/B _21684_/X VGND VGND VPWR VPWR _21685_/X sky130_fd_sc_hd__and3_4
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23424_ _23706_/CLK _20312_/X VGND VGND VPWR VPWR _22266_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_184_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20636_ _15460_/Y _20615_/X _20629_/X _20635_/X VGND VGND VPWR VPWR _20637_/A sky130_fd_sc_hd__a211o_4
XFILLER_149_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23355_ VGND VGND VPWR VPWR _23355_/HI IRQ[31] sky130_fd_sc_hd__conb_1
X_20567_ _18876_/A _18875_/X VGND VGND VPWR VPWR _20567_/Y sky130_fd_sc_hd__nand2_4
XFILLER_165_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22306_ _16517_/A _21441_/X _22891_/A VGND VGND VPWR VPWR _22306_/X sky130_fd_sc_hd__o21a_4
XFILLER_125_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13201__A _13254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15868__A3 _15721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23286_ _23108_/X _23283_/Y _23155_/X _23285_/X VGND VGND VPWR VPWR _23286_/X sky130_fd_sc_hd__a2bb2o_4
X_20498_ _23966_/Q _20495_/C VGND VGND VPWR VPWR _20498_/X sky130_fd_sc_hd__and2_4
XFILLER_164_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25025_ _25035_/CLK _25025_/D HRESETn VGND VGND VPWR VPWR _25025_/Q sky130_fd_sc_hd__dfrtp_4
X_22237_ _21674_/X _22235_/X _22236_/X VGND VGND VPWR VPWR _22237_/X sky130_fd_sc_hd__and3_4
XANTENNA__18267__A1 _13783_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19095__A _19094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22168_ _14428_/Y _21365_/A _14445_/Y _21368_/A VGND VGND VPWR VPWR _22169_/A sky130_fd_sc_hd__o22a_4
XANTENNA__20034__A _20034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21119_ _21118_/X VGND VGND VPWR VPWR _21119_/X sky130_fd_sc_hd__buf_2
XFILLER_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19823__A _19805_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14990_ _15168_/B _24474_/Q _14989_/A _24474_/Q VGND VGND VPWR VPWR _14991_/D sky130_fd_sc_hd__a2bb2o_4
X_22099_ _24552_/Q _21064_/B _21339_/X VGND VGND VPWR VPWR _22099_/X sky130_fd_sc_hd__o21a_4
X_13941_ _13927_/A _13932_/B _13932_/C _13941_/D VGND VGND VPWR VPWR _14238_/A sky130_fd_sc_hd__and4_4
XFILLER_208_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24809__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16660_ _16660_/A VGND VGND VPWR VPWR _16668_/A sky130_fd_sc_hd__buf_2
X_13872_ _23995_/Q _13871_/X _14264_/A _13845_/Y VGND VGND VPWR VPWR _13872_/X sky130_fd_sc_hd__o22a_4
X_15611_ _15610_/Y _15608_/X _11753_/X _15608_/X VGND VGND VPWR VPWR _15611_/X sky130_fd_sc_hd__a2bb2o_4
X_12823_ _12823_/A _12823_/B _12820_/X _12823_/D VGND VGND VPWR VPWR _12824_/D sky130_fd_sc_hd__or4_4
X_24809_ _24809_/CLK _15869_/X HRESETn VGND VGND VPWR VPWR _24809_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17062__B _17333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16591_ _16591_/A VGND VGND VPWR VPWR _16591_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12487__A _12211_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18330_ _18910_/A _18910_/B _18336_/A VGND VGND VPWR VPWR _19094_/C sky130_fd_sc_hd__or3_4
XFILLER_131_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24462__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15542_ _15984_/A _14365_/B _15636_/C _15636_/D VGND VGND VPWR VPWR _21290_/A sky130_fd_sc_hd__or4_4
X_12754_ _25386_/Q _22861_/A _12838_/A _12753_/Y VGND VGND VPWR VPWR _12754_/X sky130_fd_sc_hd__o22a_4
XFILLER_187_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _22807_/A VGND VGND VPWR VPWR _22684_/B sky130_fd_sc_hd__buf_2
X_18261_ _13807_/D _18256_/X _16267_/X _24226_/Q _18241_/A VGND VGND VPWR VPWR _18261_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_98_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12558_/Y _12682_/X VGND VGND VPWR VPWR _12686_/C sky130_fd_sc_hd__or2_4
X_15473_ _14863_/Y _15471_/X _15472_/X _15471_/X VGND VGND VPWR VPWR _15473_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _16322_/Y _24356_/Q _16322_/Y _24356_/Q VGND VGND VPWR VPWR _17213_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424_ _22327_/B VGND VGND VPWR VPWR _15457_/A sky130_fd_sc_hd__buf_2
X_18192_ _18128_/A _23828_/Q VGND VGND VPWR VPWR _18194_/B sky130_fd_sc_hd__or2_4
XFILLER_230_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17143_ _16957_/Y _17127_/X VGND VGND VPWR VPWR _17143_/Y sky130_fd_sc_hd__nand2_4
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14355_ _25157_/Q _14338_/B _25156_/Q _14345_/A VGND VGND VPWR VPWR _14355_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13306_ _13374_/A _19285_/A VGND VGND VPWR VPWR _13308_/B sky130_fd_sc_hd__or2_4
XFILLER_171_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14286_ _14280_/A _14285_/X _13627_/X VGND VGND VPWR VPWR _14286_/Y sky130_fd_sc_hd__a21oi_4
X_17074_ _17062_/A _17088_/B _17006_/Y _17032_/X VGND VGND VPWR VPWR _17074_/X sky130_fd_sc_hd__or4_4
XANTENNA__15859__A3 _15710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13237_ _13167_/A _23633_/Q VGND VGND VPWR VPWR _13240_/B sky130_fd_sc_hd__or2_4
X_16025_ _15998_/A VGND VGND VPWR VPWR _16025_/X sky130_fd_sc_hd__buf_2
XFILLER_40_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13168_ _13168_/A _23858_/Q VGND VGND VPWR VPWR _13169_/C sky130_fd_sc_hd__or2_4
XFILLER_123_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12119_ _12119_/A _12119_/B VGND VGND VPWR VPWR _12119_/Y sky130_fd_sc_hd__nor2_4
X_13099_ _12321_/Y _13095_/B VGND VGND VPWR VPWR _13100_/B sky130_fd_sc_hd__nand2_4
X_17976_ _17999_/A VGND VGND VPWR VPWR _18113_/A sky130_fd_sc_hd__buf_2
XFILLER_242_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19715_ _23642_/Q VGND VGND VPWR VPWR _19715_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16927_ _16133_/Y _24270_/Q _16133_/Y _24270_/Q VGND VGND VPWR VPWR _16927_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19646_ _19646_/A VGND VGND VPWR VPWR _19646_/X sky130_fd_sc_hd__buf_2
X_16858_ _24412_/Q VGND VGND VPWR VPWR _16858_/X sky130_fd_sc_hd__buf_2
XFILLER_93_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15809_ _12329_/Y _15806_/X _11721_/X _15806_/X VGND VGND VPWR VPWR _24837_/D sky130_fd_sc_hd__a2bb2o_4
X_19577_ _19568_/Y _19576_/X _19414_/X _19576_/X VGND VGND VPWR VPWR _19577_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16789_ _24446_/Q VGND VGND VPWR VPWR _16789_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18528_ _18528_/A _18528_/B VGND VGND VPWR VPWR _18530_/B sky130_fd_sc_hd__or2_4
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15204__C _15059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24132__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18459_ _18459_/A VGND VGND VPWR VPWR _18499_/A sky130_fd_sc_hd__inv_2
XFILLER_194_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21470_ _21661_/A _20343_/Y VGND VGND VPWR VPWR _21472_/B sky130_fd_sc_hd__or2_4
X_20421_ _23379_/Q VGND VGND VPWR VPWR _21617_/B sky130_fd_sc_hd__inv_2
XFILLER_147_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16943__A2_N _24261_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25338__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23140_ _16806_/A _23138_/X _23001_/X _23139_/X VGND VGND VPWR VPWR _23141_/C sky130_fd_sc_hd__a211o_4
X_20352_ _20352_/A VGND VGND VPWR VPWR _22243_/B sky130_fd_sc_hd__inv_2
X_23071_ _23005_/A _23071_/B _23071_/C VGND VGND VPWR VPWR _23072_/D sky130_fd_sc_hd__and3_4
X_20283_ _23434_/Q VGND VGND VPWR VPWR _20283_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12860__A _12769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22022_ _22014_/A _19945_/Y VGND VGND VPWR VPWR _22024_/B sky130_fd_sc_hd__or2_4
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24973__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23973_ _23972_/CLK _14790_/A HRESETn VGND VGND VPWR VPWR _20261_/B sky130_fd_sc_hd__dfstp_4
XFILLER_68_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24902__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22924_ _23060_/A _22924_/B VGND VGND VPWR VPWR _22924_/Y sky130_fd_sc_hd__nor2_4
XFILLER_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_112_0_HCLK clkbuf_7_56_0_HCLK/X VGND VGND VPWR VPWR _25375_/CLK sky130_fd_sc_hd__clkbuf_1
X_22855_ _22848_/Y _22853_/Y _22854_/X VGND VGND VPWR VPWR _22856_/D sky130_fd_sc_hd__o21a_4
XFILLER_216_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16983__A1 _24718_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_175_0_HCLK clkbuf_7_87_0_HCLK/X VGND VGND VPWR VPWR _23846_/CLK sky130_fd_sc_hd__clkbuf_1
X_21806_ _21670_/X _21806_/B VGND VGND VPWR VPWR _21806_/X sky130_fd_sc_hd__or2_4
X_22786_ _22468_/A VGND VGND VPWR VPWR _22786_/X sky130_fd_sc_hd__buf_2
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15522__A2_N _15519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21737_ _22928_/A VGND VGND VPWR VPWR _21737_/X sky130_fd_sc_hd__buf_2
X_24525_ _24555_/CLK _24525_/D HRESETn VGND VGND VPWR VPWR _24525_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12470_ _12207_/A _12469_/Y VGND VGND VPWR VPWR _12470_/X sky130_fd_sc_hd__or2_4
XANTENNA__22808__A1 _16494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21668_ _21453_/X _21668_/B _21668_/C VGND VGND VPWR VPWR _21668_/X sky130_fd_sc_hd__or3_4
X_24456_ _24443_/CLK _24456_/D HRESETn VGND VGND VPWR VPWR _15018_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20619_ _17385_/A _17385_/B VGND VGND VPWR VPWR _20619_/Y sky130_fd_sc_hd__nand2_4
X_23407_ _23441_/CLK _23407_/D VGND VGND VPWR VPWR _23407_/Q sky130_fd_sc_hd__dfxtp_4
X_24387_ _24390_/CLK _17114_/Y HRESETn VGND VGND VPWR VPWR _17029_/A sky130_fd_sc_hd__dfrtp_4
X_21599_ _13640_/A _21597_/X _13109_/A _21598_/X VGND VGND VPWR VPWR _21599_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25079__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14140_ _14118_/X _14139_/X _25138_/Q _14125_/X VGND VGND VPWR VPWR _14140_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__16499__B1 _16226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12782__A1_N _25385_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23338_ _23319_/X _23322_/X _23326_/Y _23337_/X VGND VGND VPWR VPWR HRDATA[31] sky130_fd_sc_hd__a211o_4
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25008__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14071_ _14007_/A _14070_/X _14067_/X _25234_/Q _14065_/X VGND VGND VPWR VPWR _14071_/X
+ sky130_fd_sc_hd__a32o_4
X_23269_ _12770_/Y _21863_/X _22280_/X _12534_/Y _22294_/X VGND VGND VPWR VPWR _23269_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_106_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13022_ _12308_/Y _13017_/X VGND VGND VPWR VPWR _13023_/C sky130_fd_sc_hd__nand2_4
XFILLER_4_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25008_ _25015_/CLK _25008_/D HRESETn VGND VGND VPWR VPWR _14902_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_106_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13585__B _21283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17830_ _17818_/A _17826_/B _17830_/C VGND VGND VPWR VPWR _24275_/D sky130_fd_sc_hd__and3_4
XFILLER_248_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16671__B1 _16397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23075__A _24571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17761_ _17761_/A _16921_/Y _16911_/Y _17760_/Y VGND VGND VPWR VPWR _17762_/D sky130_fd_sc_hd__or4_4
XFILLER_66_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14973_ _14972_/Y _16796_/A _14972_/Y _16796_/A VGND VGND VPWR VPWR _14973_/X sky130_fd_sc_hd__a2bb2o_4
X_19500_ _23714_/Q VGND VGND VPWR VPWR _22351_/B sky130_fd_sc_hd__inv_2
X_16712_ _16711_/Y _16709_/X _16435_/X _16709_/X VGND VGND VPWR VPWR _24481_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24643__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13924_ _13924_/A _13938_/B _13913_/X _13937_/A VGND VGND VPWR VPWR _13925_/A sky130_fd_sc_hd__or4_4
XFILLER_207_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17692_ _17521_/Y _17696_/B VGND VGND VPWR VPWR _17697_/A sky130_fd_sc_hd__or2_4
Xclkbuf_7_71_0_HCLK clkbuf_7_71_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_71_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16423__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19431_ _19430_/Y _19426_/X _19408_/X _19426_/A VGND VGND VPWR VPWR _23739_/D sky130_fd_sc_hd__a2bb2o_4
X_16643_ _16655_/A VGND VGND VPWR VPWR _16643_/X sky130_fd_sc_hd__buf_2
XFILLER_47_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13855_ _20673_/A _13850_/X _25250_/Q _13852_/X VGND VGND VPWR VPWR _13855_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16974__A1 _24740_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12806_ _12806_/A VGND VGND VPWR VPWR _12830_/C sky130_fd_sc_hd__inv_2
X_19362_ _19362_/A VGND VGND VPWR VPWR _19362_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16574_ _16574_/A VGND VGND VPWR VPWR _16574_/Y sky130_fd_sc_hd__inv_2
X_13786_ _13774_/Y _13784_/X _13785_/X _13784_/X VGND VGND VPWR VPWR _25275_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23971__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22419__A _21748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18313_ _18313_/A VGND VGND VPWR VPWR _18320_/A sky130_fd_sc_hd__inv_2
X_15525_ _15523_/Y _15519_/X HADDR[7] _15524_/X VGND VGND VPWR VPWR _15525_/X sky130_fd_sc_hd__a2bb2o_4
X_12737_ _12878_/A VGND VGND VPWR VPWR _12879_/A sky130_fd_sc_hd__inv_2
X_19293_ _19292_/Y _19290_/X _19203_/X _19290_/X VGND VGND VPWR VPWR _19293_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_231_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23241__C _23240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18244_ _18238_/X _18240_/X _16236_/A _22620_/A _18241_/X VGND VGND VPWR VPWR _18244_/X
+ sky130_fd_sc_hd__a32o_4
X_15456_ _24958_/Q VGND VGND VPWR VPWR _15456_/Y sky130_fd_sc_hd__inv_2
X_12668_ _12671_/A _12668_/B VGND VGND VPWR VPWR _12672_/B sky130_fd_sc_hd__or2_4
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _14407_/A VGND VGND VPWR VPWR _14407_/X sky130_fd_sc_hd__buf_2
X_18175_ _17972_/A _18175_/B VGND VGND VPWR VPWR _18175_/X sky130_fd_sc_hd__or2_4
XANTENNA__19728__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15387_ _15294_/C _15386_/X VGND VGND VPWR VPWR _15400_/B sky130_fd_sc_hd__or2_4
X_12599_ _12596_/Y _12655_/A _12598_/X VGND VGND VPWR VPWR _12599_/X sky130_fd_sc_hd__or3_4
XFILLER_117_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17126_ _17039_/Y _17126_/B VGND VGND VPWR VPWR _17126_/X sky130_fd_sc_hd__or2_4
X_14338_ _14338_/A _14338_/B VGND VGND VPWR VPWR _14339_/C sky130_fd_sc_hd__or2_4
XFILLER_190_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17057_ _17047_/C _17069_/B VGND VGND VPWR VPWR _17057_/X sky130_fd_sc_hd__or2_4
XFILLER_116_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14269_ _15432_/A VGND VGND VPWR VPWR _14269_/X sky130_fd_sc_hd__buf_2
XANTENNA__12680__A _12680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16152__A _22153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16008_ _16006_/Y _16007_/X _15567_/X _16007_/X VGND VGND VPWR VPWR _16008_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15991__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18651__B2 _18613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16662__B1 _16301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17959_ _17944_/A _17959_/B VGND VGND VPWR VPWR _17959_/X sky130_fd_sc_hd__or2_4
XANTENNA__24384__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20970_ _24101_/Q _12150_/Y VGND VGND VPWR VPWR _20970_/Y sky130_fd_sc_hd__nor2_4
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14400__A _14400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25137__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16414__B1 _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24313__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19629_ _13228_/B VGND VGND VPWR VPWR _19629_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22640_ _15603_/Y _22756_/B VGND VGND VPWR VPWR _22640_/X sky130_fd_sc_hd__and2_4
XFILLER_213_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_248_0_HCLK clkbuf_7_124_0_HCLK/X VGND VGND VPWR VPWR _24139_/CLK sky130_fd_sc_hd__clkbuf_1
X_22571_ _22570_/X VGND VGND VPWR VPWR _22571_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16717__B2 _16655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12581__A2_N _24885_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25519__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21522_ _21298_/X VGND VGND VPWR VPWR _21522_/X sky130_fd_sc_hd__buf_2
X_24310_ _24310_/CLK _24310_/D HRESETn VGND VGND VPWR VPWR _17507_/A sky130_fd_sc_hd__dfrtp_4
X_25290_ _24236_/CLK _13702_/X HRESETn VGND VGND VPWR VPWR _25290_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24241_ _24341_/CLK _18237_/X HRESETn VGND VGND VPWR VPWR _11811_/A sky130_fd_sc_hd__dfrtp_4
X_21453_ _18314_/Y VGND VGND VPWR VPWR _21453_/X sky130_fd_sc_hd__buf_2
XANTENNA__19667__B1 _19543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18542__A _18467_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20404_ _20403_/Y _20401_/X _11788_/X _20401_/X VGND VGND VPWR VPWR _23386_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24172_ _24172_/CLK _24172_/D HRESETn VGND VGND VPWR VPWR _18465_/A sky130_fd_sc_hd__dfrtp_4
X_21384_ _14668_/X _21384_/B VGND VGND VPWR VPWR _21384_/X sky130_fd_sc_hd__or2_4
XFILLER_107_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23123_ _22469_/X VGND VGND VPWR VPWR _23123_/X sky130_fd_sc_hd__buf_2
X_20335_ _20333_/Y _20329_/X _19606_/A _20334_/X VGND VGND VPWR VPWR _23415_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12590__A _12617_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16062__A _14407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23054_ _12232_/Y _22984_/X _17744_/A _22914_/X VGND VGND VPWR VPWR _23054_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20266_ _20266_/A VGND VGND VPWR VPWR _20266_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22005_ _22004_/X VGND VGND VPWR VPWR _22005_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24339__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20197_ _21245_/B _20192_/X _20133_/X _20180_/A VGND VGND VPWR VPWR _23467_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16653__B1 _16382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21408__A _22197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13467__B1 _11765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21529__B2 _22522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11970_ _11956_/X VGND VGND VPWR VPWR _11970_/Y sky130_fd_sc_hd__inv_2
X_23956_ _23932_/CLK _23956_/D HRESETn VGND VGND VPWR VPWR _23956_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24054__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_58_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22907_ _22907_/A VGND VGND VPWR VPWR _22907_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23887_ _23887_/CLK _19014_/X VGND VGND VPWR VPWR _18083_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_204_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13640_ _13640_/A _13640_/B VGND VGND VPWR VPWR _13640_/X sky130_fd_sc_hd__and2_4
XFILLER_244_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22838_ _21030_/A VGND VGND VPWR VPWR _22838_/X sky130_fd_sc_hd__buf_2
XANTENNA__23342__B _23342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _25083_/Q VGND VGND VPWR VPWR _14549_/B sky130_fd_sc_hd__inv_2
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12549__A2_N _12547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22769_ _22769_/A _22768_/X VGND VGND VPWR VPWR _22781_/B sky130_fd_sc_hd__and2_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15310_ _15282_/B VGND VGND VPWR VPWR _15313_/A sky130_fd_sc_hd__buf_2
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12522_ _25420_/Q _12521_/A _12597_/A _12521_/Y VGND VGND VPWR VPWR _12532_/A sky130_fd_sc_hd__o22a_4
X_24508_ _24508_/CLK _16646_/X HRESETn VGND VGND VPWR VPWR _16645_/A sky130_fd_sc_hd__dfrtp_4
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14719__B1 _13726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16290_ _16289_/Y _16285_/X _16004_/X _16285_/X VGND VGND VPWR VPWR _24639_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25488_ _25466_/CLK _12031_/X HRESETn VGND VGND VPWR VPWR _25488_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15241_ _15241_/A VGND VGND VPWR VPWR _15269_/A sky130_fd_sc_hd__buf_2
XFILLER_173_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12453_ _12418_/B _12447_/X _12398_/X _12450_/B VGND VGND VPWR VPWR _12454_/A sky130_fd_sc_hd__a211o_4
X_24439_ _25021_/CLK _16807_/X HRESETn VGND VGND VPWR VPWR _16806_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12384_ _12384_/A VGND VGND VPWR VPWR _12384_/Y sky130_fd_sc_hd__inv_2
X_15172_ _15168_/B _15161_/D VGND VGND VPWR VPWR _15173_/A sky130_fd_sc_hd__or2_4
XFILLER_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14123_ _23955_/D _14122_/X _20592_/A _23955_/D VGND VGND VPWR VPWR _25223_/D sky130_fd_sc_hd__a2bb2o_4
X_19980_ _19962_/Y VGND VGND VPWR VPWR _19980_/X sky130_fd_sc_hd__buf_2
XFILLER_99_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12931__C _12781_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18931_ _23914_/Q VGND VGND VPWR VPWR _18931_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24895__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14054_ _14054_/A VGND VGND VPWR VPWR _14054_/X sky130_fd_sc_hd__buf_2
XANTENNA__22702__A _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13005_ _13005_/A _12987_/X _12285_/Y _13005_/D VGND VGND VPWR VPWR _13005_/X sky130_fd_sc_hd__or4_4
XANTENNA__24824__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18862_ _16507_/Y _18791_/A _16527_/A _18787_/A VGND VGND VPWR VPWR _18862_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17813_ _17762_/D _17813_/B VGND VGND VPWR VPWR _17814_/B sky130_fd_sc_hd__or2_4
XANTENNA__16644__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18793_ _18793_/A _18793_/B _18792_/X VGND VGND VPWR VPWR _18793_/X sky130_fd_sc_hd__and3_4
XFILLER_208_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17744_ _17744_/A VGND VGND VPWR VPWR _17764_/A sky130_fd_sc_hd__inv_2
X_14956_ _15061_/A VGND VGND VPWR VPWR _15229_/A sky130_fd_sc_hd__buf_2
XFILLER_236_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21037__B _21064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22193__A1 _25526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13907_ _13907_/A _13907_/B _13907_/C _13883_/Y VGND VGND VPWR VPWR _13907_/X sky130_fd_sc_hd__and4_4
X_17675_ _17499_/Y _17671_/X VGND VGND VPWR VPWR _17676_/C sky130_fd_sc_hd__nand2_4
X_14887_ _25014_/Q _14885_/Y _15182_/A _24441_/Q VGND VGND VPWR VPWR _14891_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16947__B2 _24261_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19414_ _19006_/A VGND VGND VPWR VPWR _19414_/X sky130_fd_sc_hd__buf_2
X_16626_ _13728_/A VGND VGND VPWR VPWR _16628_/A sky130_fd_sc_hd__inv_2
X_13838_ _13837_/Y _13810_/A _13798_/X _13810_/A VGND VGND VPWR VPWR _13838_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23252__B _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22149__A _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19345_ _23769_/Q VGND VGND VPWR VPWR _19345_/Y sky130_fd_sc_hd__inv_2
X_16557_ _16557_/A VGND VGND VPWR VPWR _16557_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_1_0_HCLK clkbuf_6_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_13769_ _13768_/X VGND VGND VPWR VPWR _13769_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16147__A _22405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_15_0_HCLK clkbuf_7_7_0_HCLK/X VGND VGND VPWR VPWR _23559_/CLK sky130_fd_sc_hd__clkbuf_1
X_15508_ _24938_/Q VGND VGND VPWR VPWR _15508_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19276_ _19290_/A VGND VGND VPWR VPWR _19276_/X sky130_fd_sc_hd__buf_2
X_16488_ _16470_/A VGND VGND VPWR VPWR _16488_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_78_0_HCLK clkbuf_8_79_0_HCLK/A VGND VGND VPWR VPWR _24681_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_175_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18227_ _18227_/A _18227_/B _18227_/C VGND VGND VPWR VPWR _18228_/C sky130_fd_sc_hd__or3_4
X_15439_ _15429_/A VGND VGND VPWR VPWR _15439_/X sky130_fd_sc_hd__buf_2
XANTENNA__15922__A2 _15783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18158_ _18126_/A _18158_/B VGND VGND VPWR VPWR _18159_/C sky130_fd_sc_hd__or2_4
XANTENNA__22175__A1_N _17366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17109_ _17105_/A _17103_/B _17108_/Y VGND VGND VPWR VPWR _24389_/D sky130_fd_sc_hd__and3_4
XFILLER_116_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18089_ _18124_/A _18085_/X _18089_/C VGND VGND VPWR VPWR _18089_/X sky130_fd_sc_hd__or3_4
X_20120_ _23496_/Q VGND VGND VPWR VPWR _20120_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24565__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20051_ _20050_/Y _20046_/X _19852_/X _20034_/A VGND VGND VPWR VPWR _20051_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18624__A1 _24539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17550__A2_N _24113_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21228__A _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16928__A1_N _16128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23810_ _23610_/CLK _23810_/D VGND VGND VPWR VPWR _19230_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_245_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24790_ _24795_/CLK _15897_/X HRESETn VGND VGND VPWR VPWR _22130_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ _20953_/A _20953_/B _13653_/X VGND VGND VPWR VPWR _20953_/X sky130_fd_sc_hd__or3_4
X_23741_ _23747_/CLK _23741_/D VGND VGND VPWR VPWR _18143_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_38_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20884_ _24048_/Q _13649_/X VGND VGND VPWR VPWR _20888_/A sky130_fd_sc_hd__or2_4
X_23672_ _23644_/CLK _23672_/D VGND VGND VPWR VPWR _13270_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25411_ _25403_/CLK _12701_/X HRESETn VGND VGND VPWR VPWR _25411_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_242_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22623_ _17246_/Y _22543_/X _22622_/Y VGND VGND VPWR VPWR _22623_/X sky130_fd_sc_hd__o21a_4
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16057__A _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25353__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14195__A1_N _20517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22554_ _22641_/B VGND VGND VPWR VPWR _22554_/X sky130_fd_sc_hd__buf_2
X_25342_ _25344_/CLK _13085_/X HRESETn VGND VGND VPWR VPWR _25342_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21898__A _22386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21505_ _23419_/Q _20307_/X _23395_/Q _22229_/B VGND VGND VPWR VPWR _21505_/X sky130_fd_sc_hd__o22a_4
XFILLER_210_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22485_ _22429_/X VGND VGND VPWR VPWR _22485_/X sky130_fd_sc_hd__buf_2
X_25273_ _25272_/CLK _25273_/D HRESETn VGND VGND VPWR VPWR _25273_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21436_ _21298_/X VGND VGND VPWR VPWR _21436_/X sky130_fd_sc_hd__buf_2
X_24224_ _23398_/CLK _18267_/X HRESETn VGND VGND VPWR VPWR _24224_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24155_ _24080_/CLK _24155_/D HRESETn VGND VGND VPWR VPWR _24155_/Q sky130_fd_sc_hd__dfrtp_4
X_21367_ _25245_/Q VGND VGND VPWR VPWR _21367_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20318_ _23421_/Q VGND VGND VPWR VPWR _20318_/X sky130_fd_sc_hd__buf_2
X_23106_ _22971_/X _23105_/X _22973_/X _24880_/Q _22974_/X VGND VGND VPWR VPWR _23107_/B
+ sky130_fd_sc_hd__a32o_4
X_24086_ _25226_/CLK _24086_/D HRESETn VGND VGND VPWR VPWR _20440_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21298_ _21297_/Y VGND VGND VPWR VPWR _21298_/X sky130_fd_sc_hd__buf_2
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22522__A _16694_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23037_ _21080_/X VGND VGND VPWR VPWR _23037_/X sky130_fd_sc_hd__buf_2
X_20249_ _22075_/B _20243_/X _16863_/A _20248_/X VGND VGND VPWR VPWR _20249_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16520__A _16520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24235__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14810_ _14810_/A _14810_/B _14796_/A VGND VGND VPWR VPWR _14811_/B sky130_fd_sc_hd__or3_4
XFILLER_67_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11664__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15790_ _15777_/X _15789_/X _15710_/X _24850_/Q _15787_/X VGND VGND VPWR VPWR _24850_/D
+ sky130_fd_sc_hd__a32o_4
X_24988_ _24976_/CLK _24988_/D HRESETn VGND VGND VPWR VPWR _24988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12112__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14741_ _14741_/A _14740_/Y VGND VGND VPWR VPWR _14741_/X sky130_fd_sc_hd__or2_4
XFILLER_218_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11953_ _11945_/A _11944_/Y _11942_/X _11952_/X VGND VGND VPWR VPWR _25501_/D sky130_fd_sc_hd__o22a_4
X_23939_ _23938_/CLK _20555_/Y HRESETn VGND VGND VPWR VPWR _23939_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14975__A _25014_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17460_ _17460_/A VGND VGND VPWR VPWR _20387_/B sky130_fd_sc_hd__inv_2
X_14672_ _14672_/A _14671_/X VGND VGND VPWR VPWR _14673_/A sky130_fd_sc_hd__and2_4
XFILLER_60_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11884_ _11856_/B _11873_/X _11883_/Y VGND VGND VPWR VPWR _11884_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_244_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16411_ _16418_/A VGND VGND VPWR VPWR _16411_/X sky130_fd_sc_hd__buf_2
X_13623_ _13622_/X VGND VGND VPWR VPWR _13623_/X sky130_fd_sc_hd__buf_2
X_17391_ _23982_/Q _20645_/A VGND VGND VPWR VPWR _17392_/B sky130_fd_sc_hd__or2_4
XANTENNA__25094__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_231_0_HCLK clkbuf_8_231_0_HCLK/A VGND VGND VPWR VPWR _24133_/CLK sky130_fd_sc_hd__clkbuf_1
X_19130_ _23846_/Q VGND VGND VPWR VPWR _19130_/Y sky130_fd_sc_hd__inv_2
X_16342_ _16341_/Y _16337_/X _16055_/X _16337_/X VGND VGND VPWR VPWR _16342_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13554_ _13552_/A _25085_/Q _13552_/Y _14550_/A VGND VGND VPWR VPWR _13565_/A sky130_fd_sc_hd__o22a_4
XFILLER_201_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25023__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14168__A1 _14166_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12505_ _25426_/Q VGND VGND VPWR VPWR _12505_/Y sky130_fd_sc_hd__inv_2
X_19061_ _19061_/A VGND VGND VPWR VPWR _19061_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16273_ _16272_/X _16270_/B VGND VGND VPWR VPWR _16273_/X sky130_fd_sc_hd__or2_4
XFILLER_146_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13485_ _13499_/A VGND VGND VPWR VPWR _13485_/X sky130_fd_sc_hd__buf_2
XFILLER_200_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18012_ _18053_/A _18012_/B VGND VGND VPWR VPWR _18015_/B sky130_fd_sc_hd__or2_4
XFILLER_185_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22416__B _22416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15224_ _15214_/C _15214_/D _15194_/X _15221_/Y VGND VGND VPWR VPWR _15225_/A sky130_fd_sc_hd__a211o_4
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21438__B1 _25521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12436_ _12234_/A _12436_/B VGND VGND VPWR VPWR _12437_/C sky130_fd_sc_hd__or2_4
XFILLER_138_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22135__C _22135_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15155_ _15294_/D _15072_/A _15296_/A _16432_/A VGND VGND VPWR VPWR _15155_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12367_ _12979_/D _24826_/Q _13097_/A _24823_/Q VGND VGND VPWR VPWR _12368_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_153_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14106_ _14106_/A _14106_/B _14092_/A VGND VGND VPWR VPWR _14106_/X sky130_fd_sc_hd__or3_4
XFILLER_113_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12298_ _25356_/Q _12296_/Y _12285_/A _12297_/Y VGND VGND VPWR VPWR _12298_/X sky130_fd_sc_hd__a2bb2o_4
X_15086_ _24997_/Q _15084_/Y _25003_/Q _15085_/Y VGND VGND VPWR VPWR _15086_/X sky130_fd_sc_hd__a2bb2o_4
X_19963_ _19962_/Y VGND VGND VPWR VPWR _19963_/X sky130_fd_sc_hd__buf_2
XFILLER_180_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22938__B1 _22924_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14037_ _13997_/X VGND VGND VPWR VPWR _14038_/D sky130_fd_sc_hd__inv_2
X_18914_ _18909_/Y _18913_/X _17415_/X _18913_/X VGND VGND VPWR VPWR _23922_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19894_ _19893_/Y _19891_/X _19620_/X _19891_/X VGND VGND VPWR VPWR _23580_/D sky130_fd_sc_hd__a2bb2o_4
X_18845_ _18841_/X _18842_/X _18845_/C _18844_/X VGND VGND VPWR VPWR _18845_/X sky130_fd_sc_hd__or4_4
XFILLER_67_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18776_ _18778_/B VGND VGND VPWR VPWR _18777_/B sky130_fd_sc_hd__inv_2
XFILLER_209_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21990__B _21867_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15988_ _15988_/A VGND VGND VPWR VPWR _15988_/X sky130_fd_sc_hd__buf_2
XFILLER_209_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12103__B1 _11775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14643__A2 _14630_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17727_ _17726_/X VGND VGND VPWR VPWR _17727_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23263__A _24475_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14939_ _24415_/Q VGND VGND VPWR VPWR _14939_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23958__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14885__A _14885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_41_0_HCLK clkbuf_6_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17658_ _17660_/B VGND VGND VPWR VPWR _17659_/B sky130_fd_sc_hd__inv_2
XFILLER_50_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16609_ _16608_/Y _16606_/X _16525_/X _16606_/X VGND VGND VPWR VPWR _24520_/D sky130_fd_sc_hd__a2bb2o_4
X_17589_ _17491_/A _17589_/B VGND VGND VPWR VPWR _17589_/X sky130_fd_sc_hd__or2_4
XFILLER_196_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19328_ _19326_/Y _19322_/X _19282_/X _19327_/X VGND VGND VPWR VPWR _19328_/X sky130_fd_sc_hd__a2bb2o_4
X_19259_ _19253_/Y VGND VGND VPWR VPWR _19259_/X sky130_fd_sc_hd__buf_2
XFILLER_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16605__A _16605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22270_ _21274_/X _22250_/X _22265_/X _22268_/Y _22269_/X VGND VGND VPWR VPWR _22270_/X
+ sky130_fd_sc_hd__o32a_4
X_21221_ _13768_/X _21219_/X _21178_/A _21220_/X VGND VGND VPWR VPWR _21222_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24746__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21152_ _12111_/Y _21151_/A _21574_/B _21151_/Y VGND VGND VPWR VPWR _21152_/X sky130_fd_sc_hd__a211o_4
XFILLER_132_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20103_ _20101_/Y _20096_/X _20102_/X _20096_/X VGND VGND VPWR VPWR _23502_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21083_ _21519_/A VGND VGND VPWR VPWR _22840_/A sky130_fd_sc_hd__buf_2
XFILLER_160_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20034_ _20034_/A VGND VGND VPWR VPWR _20034_/X sky130_fd_sc_hd__buf_2
X_24911_ _24910_/CLK _24911_/D HRESETn VGND VGND VPWR VPWR _15588_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_123_0_HCLK clkbuf_6_61_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_247_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__24506__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24842_ _25341_/CLK _24842_/D HRESETn VGND VGND VPWR VPWR _24842_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15831__B2 _15786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24773_ _25380_/CLK _15938_/X HRESETn VGND VGND VPWR VPWR _23101_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _21981_/Y _21982_/X _21983_/X _21984_/X VGND VGND VPWR VPWR _21985_/X sky130_fd_sc_hd__a211o_4
XPHY_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25534__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ _23427_/CLK _23724_/D VGND VGND VPWR VPWR _23724_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _24060_/Q _24059_/Q _20932_/B VGND VGND VPWR VPWR _20941_/B sky130_fd_sc_hd__or3_4
XFILLER_242_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _20866_/Y _20862_/X _13647_/B VGND VGND VPWR VPWR _20867_/X sky130_fd_sc_hd__o21a_4
X_23655_ _23665_/CLK _19681_/X VGND VGND VPWR VPWR _13304_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22606_ _21121_/A _22604_/X _22111_/X _22605_/X VGND VGND VPWR VPWR _22607_/B sky130_fd_sc_hd__o22a_4
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20798_ _20796_/Y _20793_/Y _20797_/X VGND VGND VPWR VPWR _20798_/X sky130_fd_sc_hd__o21a_4
X_23586_ _23559_/CLK _19880_/X VGND VGND VPWR VPWR _19876_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_139_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25325_ _25325_/CLK _25325_/D HRESETn VGND VGND VPWR VPWR _25325_/Q sky130_fd_sc_hd__dfrtp_4
X_22537_ _15018_/A _22534_/X _22536_/X VGND VGND VPWR VPWR _22537_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_8_61_0_HCLK clkbuf_7_30_0_HCLK/X VGND VGND VPWR VPWR _24341_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_155_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13270_ _13227_/X _13270_/B VGND VGND VPWR VPWR _13270_/X sky130_fd_sc_hd__or2_4
X_25256_ _25260_/CLK _25256_/D HRESETn VGND VGND VPWR VPWR _25256_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22468_ _22468_/A _22468_/B VGND VGND VPWR VPWR _22472_/C sky130_fd_sc_hd__nor2_4
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12221_ _12268_/A _12219_/Y _12217_/A _12220_/Y VGND VGND VPWR VPWR _12228_/B sky130_fd_sc_hd__a2bb2o_4
X_24207_ _24208_/CLK _24207_/D HRESETn VGND VGND VPWR VPWR _19208_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__11659__A _11659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22093__B1 _21339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24487__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21419_ _21419_/A _21419_/B _21419_/C _21418_/Y VGND VGND VPWR VPWR _21419_/X sky130_fd_sc_hd__or4_4
XFILLER_170_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18836__A1 _16494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22399_ _22399_/A VGND VGND VPWR VPWR _22399_/Y sky130_fd_sc_hd__inv_2
X_25187_ _25249_/CLK _14260_/X HRESETn VGND VGND VPWR VPWR _25187_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18836__B2 _18692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12152_ _18372_/A _20971_/B _12151_/X VGND VGND VPWR VPWR _25468_/D sky130_fd_sc_hd__a21o_4
XANTENNA__24416__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24138_ _24139_/CLK _24138_/D HRESETn VGND VGND VPWR VPWR _24138_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21840__B1 _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_2_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12083_ _12083_/A VGND VGND VPWR VPWR _12084_/A sky130_fd_sc_hd__inv_2
X_16960_ _16955_/X _16956_/X _16960_/C _16959_/X VGND VGND VPWR VPWR _16987_/A sky130_fd_sc_hd__or4_4
X_24069_ _25346_/CLK _24069_/D HRESETn VGND VGND VPWR VPWR _24069_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15911_ _14764_/A _15690_/A _15908_/X _15910_/Y VGND VGND VPWR VPWR _15911_/X sky130_fd_sc_hd__a211o_4
XFILLER_150_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16891_ _16101_/Y _24283_/Q _16101_/Y _24283_/Q VGND VGND VPWR VPWR _16891_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20946__A2 _20846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18630_ _24155_/Q VGND VGND VPWR VPWR _18707_/A sky130_fd_sc_hd__inv_2
XFILLER_77_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15842_ _15665_/X _15700_/X _15838_/X _12968_/A _15841_/X VGND VGND VPWR VPWR _24817_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22148__A1 _24721_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18561_ _18589_/A _18420_/Y _18561_/C _18587_/B VGND VGND VPWR VPWR _18562_/B sky130_fd_sc_hd__or4_4
X_15773_ _15773_/A _15773_/B VGND VGND VPWR VPWR _15773_/X sky130_fd_sc_hd__or2_4
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12985_ _12340_/Y _12985_/B _12984_/X VGND VGND VPWR VPWR _12985_/X sky130_fd_sc_hd__or3_4
XFILLER_218_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13833__B1 _13788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22699__A2 _22697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15016__D _15015_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17512_ _11687_/A _24315_/Q _11687_/Y _17511_/Y VGND VGND VPWR VPWR _17512_/X sky130_fd_sc_hd__o22a_4
X_14724_ _22044_/A _14735_/B VGND VGND VPWR VPWR _14724_/Y sky130_fd_sc_hd__nand2_4
XFILLER_205_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_28_0_HCLK clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_11936_ _17443_/A VGND VGND VPWR VPWR _11938_/A sky130_fd_sc_hd__buf_2
X_18492_ _16441_/X _18483_/D VGND VGND VPWR VPWR _18493_/B sky130_fd_sc_hd__or2_4
XFILLER_73_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21371__A2 _14182_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17443_ _17443_/A _18902_/D VGND VGND VPWR VPWR _17443_/X sky130_fd_sc_hd__or2_4
XFILLER_232_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14655_ _19341_/A _14648_/X _14654_/X VGND VGND VPWR VPWR _14655_/Y sky130_fd_sc_hd__a21oi_4
X_11867_ _11796_/A _11865_/Y _11864_/B _11866_/X VGND VGND VPWR VPWR _25518_/D sky130_fd_sc_hd__o22a_4
XPHY_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13606_ _13606_/A _13606_/B VGND VGND VPWR VPWR _14647_/B sky130_fd_sc_hd__or2_4
XPHY_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17374_ _17242_/B _17374_/B VGND VGND VPWR VPWR _17374_/X sky130_fd_sc_hd__or2_4
XFILLER_60_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14586_ _14555_/X _14575_/X _14585_/Y _14579_/X _14548_/A VGND VGND VPWR VPWR _25090_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11798_ _25515_/Q VGND VGND VPWR VPWR _11799_/A sky130_fd_sc_hd__inv_2
XANTENNA__22427__A _22394_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19113_ _19113_/A VGND VGND VPWR VPWR _19113_/Y sky130_fd_sc_hd__inv_2
X_16325_ _16344_/A VGND VGND VPWR VPWR _16325_/X sky130_fd_sc_hd__buf_2
X_13537_ _13538_/A _14554_/A _13536_/Y _13569_/A VGND VGND VPWR VPWR _13537_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_229_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19044_ _23875_/Q VGND VGND VPWR VPWR _19044_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16256_ _21842_/A VGND VGND VPWR VPWR _16256_/Y sky130_fd_sc_hd__inv_2
X_13468_ _13468_/A VGND VGND VPWR VPWR _13468_/Y sky130_fd_sc_hd__inv_2
X_15207_ _15207_/A _15207_/B VGND VGND VPWR VPWR _15207_/X sky130_fd_sc_hd__or2_4
X_12419_ _12443_/A _12226_/X _12418_/X VGND VGND VPWR VPWR _12428_/D sky130_fd_sc_hd__or3_4
X_16187_ _23297_/A VGND VGND VPWR VPWR _16187_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22623__A2 _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18827__B2 _18769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13399_ _13431_/A _13399_/B VGND VGND VPWR VPWR _13399_/X sky130_fd_sc_hd__or2_4
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16838__B1 _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24157__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15138_ _15137_/Y _24602_/Q _15295_/A _15081_/Y VGND VGND VPWR VPWR _15138_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17256__A _17175_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15069_ _15068_/Y _24591_/Q _15068_/Y _24591_/Q VGND VGND VPWR VPWR _15077_/A sky130_fd_sc_hd__a2bb2o_4
X_19946_ _19946_/A VGND VGND VPWR VPWR _19946_/X sky130_fd_sc_hd__buf_2
XFILLER_141_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19877_ _19597_/A _18279_/X _19455_/X VGND VGND VPWR VPWR _19878_/A sky130_fd_sc_hd__or3_4
XFILLER_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18828_ _16534_/Y _18641_/A _24552_/Q _18804_/A VGND VGND VPWR VPWR _18828_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22139__A1 _22716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14616__A2 _14610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18759_ _18755_/B _18758_/X VGND VGND VPWR VPWR _18764_/B sky130_fd_sc_hd__or2_4
XANTENNA__20410__A _20409_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21770_ _22381_/A _21770_/B VGND VGND VPWR VPWR _21772_/B sky130_fd_sc_hd__or2_4
XFILLER_24_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23351__A3 HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20721_ _20720_/X VGND VGND VPWR VPWR _24010_/D sky130_fd_sc_hd__inv_2
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15577__B1 _11691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20652_ _17392_/A _17392_/B VGND VGND VPWR VPWR _20652_/Y sky130_fd_sc_hd__nand2_4
X_23440_ _23441_/CLK _20270_/X VGND VGND VPWR VPWR _23440_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24998__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22311__A1 _14917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21241__A _22069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23371_ _23371_/A VGND VGND VPWR VPWR IRQ[27] sky130_fd_sc_hd__buf_2
XANTENNA__24927__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20583_ _20583_/A VGND VGND VPWR VPWR _20583_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25110_ _23958_/CLK _14504_/X HRESETn VGND VGND VPWR VPWR _14490_/B sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_48_0_HCLK clkbuf_6_24_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_48_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22322_ _21832_/A _22321_/X VGND VGND VPWR VPWR _22322_/X sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_5_19_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22253_ _21674_/X _22253_/B _22252_/X VGND VGND VPWR VPWR _22253_/X sky130_fd_sc_hd__and3_4
X_25041_ _25056_/CLK _14878_/Y HRESETn VGND VGND VPWR VPWR _14859_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_164_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24580__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19646__A _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21204_ _21204_/A VGND VGND VPWR VPWR _21207_/A sky130_fd_sc_hd__buf_2
X_22184_ _14249_/Y _14245_/A _17417_/Y _17411_/X VGND VGND VPWR VPWR _22184_/X sky130_fd_sc_hd__o22a_4
XFILLER_144_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22090__A3 _22055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21135_ _25102_/Q _21346_/A VGND VGND VPWR VPWR _21135_/Y sky130_fd_sc_hd__nand2_4
XFILLER_99_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21066_ _21066_/A _16270_/A VGND VGND VPWR VPWR _21066_/X sky130_fd_sc_hd__and2_4
XFILLER_235_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22800__A _16404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20017_ _20017_/A VGND VGND VPWR VPWR _22016_/B sky130_fd_sc_hd__inv_2
XFILLER_247_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14607__A2 _14610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24825_ _25428_/CLK _24825_/D HRESETn VGND VGND VPWR VPWR _24825_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21416__A _21178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13815__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12770_ _12770_/A VGND VGND VPWR VPWR _12770_/Y sky130_fd_sc_hd__inv_2
X_24756_ _24766_/CLK _24756_/D HRESETn VGND VGND VPWR VPWR _24756_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21135__B _21346_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21968_ _21968_/A _19585_/X VGND VGND VPWR VPWR _21968_/X sky130_fd_sc_hd__and2_4
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22550__A1 _24525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ HWDATA[17] VGND VGND VPWR VPWR _11721_/X sky130_fd_sc_hd__buf_2
X_23707_ _23691_/CLK _23707_/D VGND VGND VPWR VPWR _23707_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ _20919_/A VGND VGND VPWR VPWR _20919_/X sky130_fd_sc_hd__buf_2
XANTENNA__15568__B1 _15567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24687_ _24686_/CLK _16151_/X HRESETn VGND VGND VPWR VPWR _22191_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_203_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ _21896_/X _21899_/B _21899_/C VGND VGND VPWR VPWR _21899_/X sky130_fd_sc_hd__and3_4
XFILLER_120_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14171_/Y _14437_/X _14389_/X _14431_/A VGND VGND VPWR VPWR _25130_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _13807_/B VGND VGND VPWR VPWR _17703_/B sky130_fd_sc_hd__inv_2
X_23638_ _23627_/CLK _23638_/D VGND VGND VPWR VPWR _19727_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_80_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23350__B _25170_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22302__A1 _25374_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24668__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _14370_/B _14369_/X _14370_/Y VGND VGND VPWR VPWR _14371_/X sky130_fd_sc_hd__a21o_4
XFILLER_128_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23569_ _25070_/CLK _19923_/X VGND VGND VPWR VPWR _19922_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23318__A1_N _22543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16110_ _22980_/A VGND VGND VPWR VPWR _16110_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _13186_/X _13321_/X _25330_/Q _13245_/X VGND VGND VPWR VPWR _25330_/D sky130_fd_sc_hd__o22a_4
X_25308_ _25308_/CLK _13502_/X HRESETn VGND VGND VPWR VPWR _25308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_156_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17090_ _17004_/Y _17090_/B VGND VGND VPWR VPWR _17091_/A sky130_fd_sc_hd__or2_4
XFILLER_183_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16041_ _16040_/Y _16038_/X _11739_/X _16038_/X VGND VGND VPWR VPWR _24729_/D sky130_fd_sc_hd__a2bb2o_4
X_13253_ _13200_/A _20226_/A VGND VGND VPWR VPWR _13253_/X sky130_fd_sc_hd__or2_4
X_25239_ _25238_/CLK _14063_/X HRESETn VGND VGND VPWR VPWR _13990_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15740__B1 _24870_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12204_ _12204_/A VGND VGND VPWR VPWR _12204_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24250__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_5_0_HCLK clkbuf_5_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13184_ _13184_/A VGND VGND VPWR VPWR _13186_/A sky130_fd_sc_hd__inv_2
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19800_ _13446_/B VGND VGND VPWR VPWR _19800_/Y sky130_fd_sc_hd__inv_2
X_12135_ _12135_/A _12116_/X VGND VGND VPWR VPWR _12135_/X sky130_fd_sc_hd__and2_4
X_17992_ _18182_/A _17992_/B VGND VGND VPWR VPWR _17992_/X sky130_fd_sc_hd__or2_4
XFILLER_111_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23228__D _23228_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16943_ _16157_/Y _24261_/Q _21435_/A _17880_/A VGND VGND VPWR VPWR _16943_/X sky130_fd_sc_hd__a2bb2o_4
X_19731_ _19723_/A VGND VGND VPWR VPWR _19731_/X sky130_fd_sc_hd__buf_2
XFILLER_238_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12066_ _12064_/Y _12060_/X _11770_/X _12065_/X VGND VGND VPWR VPWR _12066_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23030__A2 _22559_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14212__B _14212_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16874_ _16872_/Y _16865_/X _16873_/X _16865_/X VGND VGND VPWR VPWR _24409_/D sky130_fd_sc_hd__a2bb2o_4
X_19662_ _19661_/Y _19657_/X _19587_/X _19657_/X VGND VGND VPWR VPWR _23662_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15825_ _12312_/Y _15823_/X _15616_/X _15823_/X VGND VGND VPWR VPWR _15825_/X sky130_fd_sc_hd__a2bb2o_4
X_18613_ _18613_/A VGND VGND VPWR VPWR _18613_/X sky130_fd_sc_hd__buf_2
XANTENNA__21326__A _15662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19593_ _19592_/Y _19590_/X _19543_/X _19590_/X VGND VGND VPWR VPWR _19593_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_231_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11852__A _11934_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15756_ _12524_/Y _15750_/X _15754_/X _15755_/X VGND VGND VPWR VPWR _24863_/D sky130_fd_sc_hd__a2bb2o_4
X_18544_ _18466_/B _18538_/B VGND VGND VPWR VPWR _18545_/C sky130_fd_sc_hd__nand2_4
X_12968_ _12968_/A VGND VGND VPWR VPWR _12968_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13282__A1 _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14707_ _22205_/A VGND VGND VPWR VPWR _14707_/X sky130_fd_sc_hd__buf_2
XFILLER_73_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11919_ _11897_/X VGND VGND VPWR VPWR _11919_/X sky130_fd_sc_hd__buf_2
X_18475_ _24162_/Q VGND VGND VPWR VPWR _18562_/A sky130_fd_sc_hd__inv_2
X_15687_ _15687_/A VGND VGND VPWR VPWR _15687_/Y sky130_fd_sc_hd__inv_2
X_12899_ _12899_/A VGND VGND VPWR VPWR _12899_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17426_ _17426_/A VGND VGND VPWR VPWR _21722_/A sky130_fd_sc_hd__inv_2
X_14638_ _13590_/A VGND VGND VPWR VPWR _14639_/A sky130_fd_sc_hd__inv_2
XANTENNA__23097__A2 _23095_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17357_ _24350_/Q _17357_/B VGND VGND VPWR VPWR _17359_/B sky130_fd_sc_hd__or2_4
XFILLER_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14569_ _14569_/A VGND VGND VPWR VPWR _14570_/B sky130_fd_sc_hd__inv_2
XFILLER_147_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16308_ _22944_/A VGND VGND VPWR VPWR _16308_/Y sky130_fd_sc_hd__inv_2
X_17288_ _17219_/Y _17253_/X _17343_/B VGND VGND VPWR VPWR _17288_/X sky130_fd_sc_hd__or3_4
X_19027_ _19026_/X VGND VGND VPWR VPWR _19028_/A sky130_fd_sc_hd__buf_2
XFILLER_173_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16239_ _16239_/A VGND VGND VPWR VPWR _16239_/X sky130_fd_sc_hd__buf_2
XANTENNA__20607__A1 _20601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14403__A _14403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19929_ _19929_/A VGND VGND VPWR VPWR _19929_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18833__A1_N _16530_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13019__A _13028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22940_ _16485_/A _22817_/B _23075_/C VGND VGND VPWR VPWR _22940_/X sky130_fd_sc_hd__and3_4
XFILLER_84_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25126__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22871_ _11681_/B _22870_/X _22495_/X _11717_/A _15983_/X VGND VGND VPWR VPWR _22871_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21106__A1_N _21736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24610_ _24597_/CLK _24610_/D HRESETn VGND VGND VPWR VPWR _24610_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_225_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21822_ _21822_/A _21649_/X VGND VGND VPWR VPWR _21827_/B sky130_fd_sc_hd__or2_4
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24541_ _24540_/CLK _24541_/D HRESETn VGND VGND VPWR VPWR _16554_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_11_0_HCLK clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21753_ _21771_/A _19242_/Y VGND VGND VPWR VPWR _21753_/X sky130_fd_sc_hd__or2_4
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20704_ _20704_/A VGND VGND VPWR VPWR _20704_/Y sky130_fd_sc_hd__inv_2
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24472_ _25028_/CLK _24472_/D HRESETn VGND VGND VPWR VPWR _15046_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21684_ _21817_/A _21684_/B VGND VGND VPWR VPWR _21684_/X sky130_fd_sc_hd__or2_4
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22067__A _22365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23423_ _23706_/CLK _23423_/D VGND VGND VPWR VPWR _22003_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24761__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20635_ _17389_/B _20634_/Y _20621_/C VGND VGND VPWR VPWR _20635_/X sky130_fd_sc_hd__and3_4
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16065__A _15988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15970__B1 _15616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12593__A _12592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19161__B1 _19138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24079__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20566_ _20543_/A VGND VGND VPWR VPWR _20566_/X sky130_fd_sc_hd__buf_2
X_23354_ VGND VGND VPWR VPWR _23354_/HI IRQ[30] sky130_fd_sc_hd__conb_1
XFILLER_166_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24008__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22305_ _24654_/Q _22932_/A VGND VGND VPWR VPWR _22308_/B sky130_fd_sc_hd__or2_4
XFILLER_180_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20497_ _20485_/X _20497_/B VGND VGND VPWR VPWR _20497_/X sky130_fd_sc_hd__or2_4
X_23285_ _22552_/X _23284_/X _22135_/C _24113_/Q _22555_/X VGND VGND VPWR VPWR _23285_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_106_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25024_ _25028_/CLK _25024_/D HRESETn VGND VGND VPWR VPWR _14892_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22236_ _22015_/A _22236_/B VGND VGND VPWR VPWR _22236_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_135_0_HCLK clkbuf_7_67_0_HCLK/X VGND VGND VPWR VPWR _23452_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_161_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_198_0_HCLK clkbuf_7_99_0_HCLK/X VGND VGND VPWR VPWR _24594_/CLK sky130_fd_sc_hd__clkbuf_1
X_22167_ _14375_/Y _21849_/X VGND VGND VPWR VPWR _22174_/A sky130_fd_sc_hd__nor2_4
X_21118_ _21832_/A VGND VGND VPWR VPWR _21118_/X sky130_fd_sc_hd__buf_2
X_22098_ _22928_/A VGND VGND VPWR VPWR _22098_/X sky130_fd_sc_hd__buf_2
X_13940_ _13940_/A VGND VGND VPWR VPWR _13941_/D sky130_fd_sc_hd__inv_2
X_21049_ _21016_/A _21048_/Y VGND VGND VPWR VPWR _21049_/X sky130_fd_sc_hd__and2_4
XFILLER_247_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16053__A1_N _16052_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13871_ _25244_/Q _13849_/X _23442_/Q _13844_/X VGND VGND VPWR VPWR _13871_/X sky130_fd_sc_hd__o22a_4
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17343__B _17343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15610_ _24902_/Q VGND VGND VPWR VPWR _15610_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12822_ _12948_/A _22295_/A _12816_/Y _24788_/Q VGND VGND VPWR VPWR _12823_/D sky130_fd_sc_hd__a2bb2o_4
X_24808_ _24834_/CLK _24808_/D HRESETn VGND VGND VPWR VPWR _24808_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_216_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15144__A _24602_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16590_ _16589_/Y _16585_/X _16236_/X _16585_/X VGND VGND VPWR VPWR _16590_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15541_ _15541_/A _14177_/B VGND VGND VPWR VPWR _15636_/D sky130_fd_sc_hd__or2_4
XFILLER_243_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23361__A _23348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24849__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12753_ _22861_/A VGND VGND VPWR VPWR _12753_/Y sky130_fd_sc_hd__inv_2
X_24739_ _25538_/CLK _16015_/X HRESETn VGND VGND VPWR VPWR _16014_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18455__A _18774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11704_/A VGND VGND VPWR VPWR _22807_/A sky130_fd_sc_hd__buf_2
X_18260_ _11830_/Y _18236_/A _16787_/X _18236_/A VGND VGND VPWR VPWR _24227_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15472_/A VGND VGND VPWR VPWR _15472_/X sky130_fd_sc_hd__buf_2
XFILLER_15_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12684_/A _12684_/B VGND VGND VPWR VPWR _12686_/B sky130_fd_sc_hd__or2_4
XFILLER_42_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _16315_/Y _17200_/A _24633_/Q _17249_/C VGND VGND VPWR VPWR _17211_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _21365_/A VGND VGND VPWR VPWR _22327_/B sky130_fd_sc_hd__buf_2
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18191_ _18094_/A _18191_/B _18190_/X VGND VGND VPWR VPWR _18195_/B sky130_fd_sc_hd__and3_4
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15961__B1 _24761_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19152__B1 _19057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17142_ _17142_/A _17129_/X _17141_/Y VGND VGND VPWR VPWR _24380_/D sky130_fd_sc_hd__and3_4
XANTENNA__24431__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14354_ _14344_/X _14353_/X _25483_/Q _14349_/X VGND VGND VPWR VPWR _25158_/D sky130_fd_sc_hd__o22a_4
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13305_ _13219_/X _13303_/X _13304_/X VGND VGND VPWR VPWR _13305_/X sky130_fd_sc_hd__and3_4
XFILLER_128_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_31_0_HCLK clkbuf_7_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17073_ _17073_/A VGND VGND VPWR VPWR _17073_/Y sky130_fd_sc_hd__inv_2
X_14285_ _14285_/A _14296_/A VGND VGND VPWR VPWR _14285_/X sky130_fd_sc_hd__or2_4
XANTENNA__16703__A _24484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_94_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_94_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_16024_ _24735_/Q VGND VGND VPWR VPWR _16024_/Y sky130_fd_sc_hd__inv_2
X_13236_ _13231_/X _13233_/X _13235_/X VGND VGND VPWR VPWR _13236_/X sky130_fd_sc_hd__and3_4
XFILLER_156_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13167_ _13167_/A _19046_/A VGND VGND VPWR VPWR _13169_/B sky130_fd_sc_hd__or2_4
XFILLER_124_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12118_ _24105_/Q _12129_/A _12117_/Y VGND VGND VPWR VPWR _12119_/B sky130_fd_sc_hd__o21a_4
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13098_ _13098_/A _13098_/B _13091_/C VGND VGND VPWR VPWR _25338_/D sky130_fd_sc_hd__and3_4
X_17975_ _13597_/A VGND VGND VPWR VPWR _17999_/A sky130_fd_sc_hd__buf_2
XANTENNA__25290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_HCLK clkbuf_3_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19714_ _19713_/Y _19707_/X _19646_/X _19694_/A VGND VGND VPWR VPWR _19714_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12049_ _12049_/A VGND VGND VPWR VPWR _12049_/Y sky130_fd_sc_hd__inv_2
X_16926_ _21435_/A _17880_/A _22153_/A _16925_/Y VGND VGND VPWR VPWR _16929_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19645_ _13439_/B VGND VGND VPWR VPWR _19645_/Y sky130_fd_sc_hd__inv_2
X_16857_ _16855_/Y _16856_/X RsRx_S0 _16856_/X VGND VGND VPWR VPWR _16857_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15808_ _12325_/Y _15806_/X _11718_/X _15806_/X VGND VGND VPWR VPWR _15808_/X sky130_fd_sc_hd__a2bb2o_4
X_16788_ _16786_/Y _16726_/A _16787_/X _16726_/A VGND VGND VPWR VPWR _16788_/X sky130_fd_sc_hd__a2bb2o_4
X_19576_ _19576_/A VGND VGND VPWR VPWR _19576_/X sky130_fd_sc_hd__buf_2
XFILLER_225_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15739_ HWDATA[15] VGND VGND VPWR VPWR _15739_/X sky130_fd_sc_hd__buf_2
X_18527_ _18526_/X VGND VGND VPWR VPWR _18528_/B sky130_fd_sc_hd__inv_2
XANTENNA__15989__A _15988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15204__D _15242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24519__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18458_ _18440_/Y _18505_/A VGND VGND VPWR VPWR _18493_/A sky130_fd_sc_hd__or2_4
XFILLER_178_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14204__B1 _13798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17409_ _20628_/A VGND VGND VPWR VPWR _20672_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_3_5_0_HCLK_A clkbuf_3_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18389_ _18388_/Y _18386_/X _24191_/Q _18386_/X VGND VGND VPWR VPWR _18389_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15952__B1 _15951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20420_ _21762_/B _20415_/X _19820_/A _20415_/X VGND VGND VPWR VPWR _23380_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24172__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24101__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20351_ _22357_/B _20350_/X _19600_/A _20350_/X VGND VGND VPWR VPWR _23409_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17709__A _17709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23070_ _16810_/A _22807_/X _23001_/X _23069_/X VGND VGND VPWR VPWR _23071_/C sky130_fd_sc_hd__a211o_4
X_20282_ _20281_/Y _20279_/X _19984_/X _20279_/X VGND VGND VPWR VPWR _20282_/X sky130_fd_sc_hd__a2bb2o_4
X_22021_ _22021_/A _22019_/X _22020_/X VGND VGND VPWR VPWR _22021_/X sky130_fd_sc_hd__and3_4
XANTENNA__25378__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11757__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_208_0_HCLK clkbuf_7_104_0_HCLK/X VGND VGND VPWR VPWR _24049_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_170_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25307__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22350__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17444__A _13584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23972_ _23972_/CLK _23972_/D HRESETn VGND VGND VPWR VPWR _23972_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_68_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22923_ _22786_/X _22921_/X _22789_/X _22922_/X VGND VGND VPWR VPWR _22924_/B sky130_fd_sc_hd__o22a_4
XFILLER_84_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22854_ _23328_/A VGND VGND VPWR VPWR _22854_/X sky130_fd_sc_hd__buf_2
XFILLER_232_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21805_ _21453_/X _21797_/X _21805_/C VGND VGND VPWR VPWR _21805_/X sky130_fd_sc_hd__or3_4
XANTENNA__24942__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22785_ _22686_/A VGND VGND VPWR VPWR _23060_/A sky130_fd_sc_hd__buf_2
XFILLER_197_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24524_ _24555_/CLK _16599_/X HRESETn VGND VGND VPWR VPWR _24524_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21736_ _21736_/A VGND VGND VPWR VPWR _22928_/A sky130_fd_sc_hd__buf_2
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16196__B1 _16004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24455_ _24443_/CLK _16770_/X HRESETn VGND VGND VPWR VPWR _15008_/A sky130_fd_sc_hd__dfrtp_4
X_21667_ _21663_/X _21666_/X _18301_/X VGND VGND VPWR VPWR _21668_/C sky130_fd_sc_hd__o21a_4
XFILLER_212_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15943__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19134__B1 _19063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23406_ _23406_/CLK _20358_/X VGND VGND VPWR VPWR _20357_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__13212__A _13334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20618_ _20618_/A VGND VGND VPWR VPWR _20618_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24386_ _24377_/CLK _24386_/D HRESETn VGND VGND VPWR VPWR _24386_/Q sky130_fd_sc_hd__dfrtp_4
X_21598_ _21598_/A VGND VGND VPWR VPWR _21598_/X sky130_fd_sc_hd__buf_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22525__A _22525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23337_ _23128_/A _23337_/B _23337_/C _23337_/D VGND VGND VPWR VPWR _23337_/X sky130_fd_sc_hd__or4_4
Xclkbuf_6_18_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20549_ _18872_/X _20547_/Y _20553_/C VGND VGND VPWR VPWR _20549_/X sky130_fd_sc_hd__and3_4
XFILLER_152_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14070_ _14054_/A VGND VGND VPWR VPWR _14070_/X sky130_fd_sc_hd__buf_2
X_23268_ _23268_/A _23267_/X VGND VGND VPWR VPWR _23268_/Y sky130_fd_sc_hd__nor2_4
XFILLER_153_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13021_ _12287_/Y _13018_/X _13020_/Y VGND VGND VPWR VPWR _13021_/X sky130_fd_sc_hd__o21a_4
X_25007_ _25204_/CLK _25007_/D HRESETn VGND VGND VPWR VPWR _15070_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14439__A1_N _14166_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22219_ _22219_/A _22217_/X _22219_/C VGND VGND VPWR VPWR _22219_/X sky130_fd_sc_hd__and3_4
XANTENNA__13585__C _25057_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23199_ _23197_/X _23198_/X _22140_/A VGND VGND VPWR VPWR _23199_/X sky130_fd_sc_hd__or3_4
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25048__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14972_ _25038_/Q VGND VGND VPWR VPWR _14972_/Y sky130_fd_sc_hd__inv_2
X_17760_ _24274_/Q VGND VGND VPWR VPWR _17760_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23075__B _23075_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13923_ _13927_/B _13914_/X _13879_/C _13923_/D VGND VGND VPWR VPWR _13937_/A sky130_fd_sc_hd__or4_4
X_16711_ _24481_/Q VGND VGND VPWR VPWR _16711_/Y sky130_fd_sc_hd__inv_2
X_17691_ _17580_/C _17665_/D VGND VGND VPWR VPWR _17696_/B sky130_fd_sc_hd__or2_4
XFILLER_207_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16642_ _16692_/A VGND VGND VPWR VPWR _16655_/A sky130_fd_sc_hd__buf_2
X_19430_ _18207_/B VGND VGND VPWR VPWR _19430_/Y sky130_fd_sc_hd__inv_2
X_13854_ _13841_/X _13853_/X VGND VGND VPWR VPWR _13854_/X sky130_fd_sc_hd__or2_4
XFILLER_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14434__B1 _14380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12805_ _12804_/Y _24807_/Q _25378_/Q _12743_/Y VGND VGND VPWR VPWR _12805_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24683__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16573_ _16571_/Y _16567_/X _16397_/X _16572_/X VGND VGND VPWR VPWR _16573_/X sky130_fd_sc_hd__a2bb2o_4
X_19361_ _19359_/Y _19356_/X _19360_/X _19356_/X VGND VGND VPWR VPWR _23764_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21604__A _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13785_ _14380_/A VGND VGND VPWR VPWR _13785_/X sky130_fd_sc_hd__buf_2
XFILLER_222_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19373__B1 _19282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15524_ _15530_/A VGND VGND VPWR VPWR _15524_/X sky130_fd_sc_hd__buf_2
X_18312_ _21665_/A _18292_/X _18305_/X VGND VGND VPWR VPWR _18312_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_43_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24612__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12736_ _25374_/Q _12734_/Y _12735_/Y _23187_/A VGND VGND VPWR VPWR _12736_/X sky130_fd_sc_hd__a2bb2o_4
X_19292_ _23788_/Q VGND VGND VPWR VPWR _19292_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18243_ _11844_/Y _18236_/X _15743_/X _18236_/X VGND VGND VPWR VPWR _24239_/D sky130_fd_sc_hd__a2bb2o_4
X_15455_ _14269_/X _24075_/Q _15436_/Y _14232_/C _15436_/B VGND VGND VPWR VPWR _24959_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22138__C _22138_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12667_ _12664_/C _12663_/X VGND VGND VPWR VPWR _12668_/B sky130_fd_sc_hd__or2_4
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15934__B1 _15560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12748__B1 _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ HWDATA[5] VGND VGND VPWR VPWR _14407_/A sky130_fd_sc_hd__buf_2
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18174_ _18027_/A _19405_/A VGND VGND VPWR VPWR _18174_/X sky130_fd_sc_hd__or2_4
X_15386_ _15294_/D _15385_/X VGND VGND VPWR VPWR _15386_/X sky130_fd_sc_hd__or2_4
X_12598_ _12664_/A _12671_/A _12598_/C VGND VGND VPWR VPWR _12598_/X sky130_fd_sc_hd__or3_4
XFILLER_184_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22435__A _22435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17125_ _17125_/A _16982_/Y _17041_/C _17124_/X VGND VGND VPWR VPWR _17126_/B sky130_fd_sc_hd__or4_4
XFILLER_7_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14337_ _14337_/A VGND VGND VPWR VPWR _14338_/B sky130_fd_sc_hd__inv_2
XFILLER_237_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17056_ _17062_/A _17056_/B VGND VGND VPWR VPWR _17069_/B sky130_fd_sc_hd__or2_4
XANTENNA__25070__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14268_ _15451_/A VGND VGND VPWR VPWR _15432_/A sky130_fd_sc_hd__buf_2
X_16007_ _15998_/A VGND VGND VPWR VPWR _16007_/X sky130_fd_sc_hd__buf_2
XFILLER_98_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13173__B1 _13150_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13219_ _13422_/A VGND VGND VPWR VPWR _13219_/X sky130_fd_sc_hd__buf_2
XFILLER_131_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14199_ _20667_/A _14187_/B VGND VGND VPWR VPWR _14199_/X sky130_fd_sc_hd__or2_4
XFILLER_171_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25400__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_181_0_HCLK clkbuf_7_90_0_HCLK/X VGND VGND VPWR VPWR _25146_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_97_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17264__A _17343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_38_0_HCLK clkbuf_8_39_0_HCLK/A VGND VGND VPWR VPWR _24199_/CLK sky130_fd_sc_hd__clkbuf_1
X_17958_ _17940_/A _17958_/B VGND VGND VPWR VPWR _17958_/X sky130_fd_sc_hd__or2_4
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16909_ _22405_/A _24265_/Q _16147_/Y _16908_/Y VGND VGND VPWR VPWR _16909_/X sky130_fd_sc_hd__o22a_4
X_17889_ _17810_/A _17850_/X _17889_/C VGND VGND VPWR VPWR _17889_/X sky130_fd_sc_hd__and3_4
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19628_ _19624_/Y _19627_/X _19414_/X _19627_/X VGND VGND VPWR VPWR _23674_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15768__A3 _15643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19559_ _23694_/Q VGND VGND VPWR VPWR _21816_/B sky130_fd_sc_hd__inv_2
XFILLER_53_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18095__A _18095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16608__A _24520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24353__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15512__A _15530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22570_ _21055_/X _22565_/X _21832_/X _22569_/Y VGND VGND VPWR VPWR _22570_/X sky130_fd_sc_hd__a211o_4
XFILLER_222_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21521_ _21521_/A _23002_/A VGND VGND VPWR VPWR _21521_/X sky130_fd_sc_hd__or2_4
XFILLER_194_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24240_ _25091_/CLK _24240_/D HRESETn VGND VGND VPWR VPWR _22696_/A sky130_fd_sc_hd__dfrtp_4
X_21452_ _21452_/A VGND VGND VPWR VPWR _21518_/C sky130_fd_sc_hd__inv_2
XFILLER_119_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20403_ _13395_/B VGND VGND VPWR VPWR _20403_/Y sky130_fd_sc_hd__inv_2
X_21383_ _13525_/Y _21281_/B _21177_/A VGND VGND VPWR VPWR _21383_/X sky130_fd_sc_hd__o21a_4
X_24171_ _24654_/CLK _24171_/D HRESETn VGND VGND VPWR VPWR _24171_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17439__A _13797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16343__A _24618_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23122_ _16654_/Y _23291_/B VGND VGND VPWR VPWR _23122_/X sky130_fd_sc_hd__and2_4
X_20334_ _20328_/Y VGND VGND VPWR VPWR _20334_/X sky130_fd_sc_hd__buf_2
X_20265_ _19939_/A _19960_/X _18284_/X VGND VGND VPWR VPWR _20266_/A sky130_fd_sc_hd__or3_4
X_23053_ _23160_/A _23039_/X _23053_/C _23053_/D VGND VGND VPWR VPWR _23053_/X sky130_fd_sc_hd__or4_4
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22004_ _20374_/Y _22001_/Y _22395_/A _22003_/Y VGND VGND VPWR VPWR _22004_/X sky130_fd_sc_hd__a211o_4
XFILLER_131_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16102__B1 _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20196_ _20196_/A VGND VGND VPWR VPWR _21245_/B sky130_fd_sc_hd__inv_2
XANTENNA__22080__A _22379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23955_ _25100_/CLK _23955_/D HRESETn VGND VGND VPWR VPWR _14523_/A sky130_fd_sc_hd__dfstp_4
XFILLER_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_9_0_HCLK clkbuf_5_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22906_ _22486_/X _22905_/X _22489_/X _24735_/Q _22865_/X VGND VGND VPWR VPWR _22907_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_217_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23886_ _23887_/CLK _23886_/D VGND VGND VPWR VPWR _18118_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14416__B1 _14384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21424__A _22451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22837_ _24597_/Q _23022_/B VGND VGND VPWR VPWR _22837_/X sky130_fd_sc_hd__or2_4
XANTENNA__16518__A _14400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11950__A _11950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24094__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13570_ _22540_/A _25093_/Q _13536_/A _14552_/A VGND VGND VPWR VPWR _13570_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22768_ _22474_/X _22767_/X _22477_/X _24836_/Q _22478_/X VGND VGND VPWR VPWR _22768_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_241_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _12521_/A VGND VGND VPWR VPWR _12521_/Y sky130_fd_sc_hd__inv_2
X_24507_ _24032_/CLK _16649_/X HRESETn VGND VGND VPWR VPWR _24507_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24023__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21719_ _21719_/A _21716_/Y _21719_/C _21719_/D VGND VGND VPWR VPWR _21719_/X sky130_fd_sc_hd__and4_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25487_ _25325_/CLK _25487_/D HRESETn VGND VGND VPWR VPWR _23350_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_13_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22699_ _22521_/B _22697_/X _22468_/A _22698_/X VGND VGND VPWR VPWR _22700_/A sky130_fd_sc_hd__o22a_4
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19107__B1 _19106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A VGND VGND VPWR VPWR _15240_/Y sky130_fd_sc_hd__inv_2
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12452_ _12434_/A _12452_/B _12452_/C VGND VGND VPWR VPWR _25446_/D sky130_fd_sc_hd__and3_4
X_24438_ _25021_/CLK _16809_/X HRESETn VGND VGND VPWR VPWR _24438_/Q sky130_fd_sc_hd__dfrtp_4
X_15171_ _15171_/A VGND VGND VPWR VPWR _15171_/Y sky130_fd_sc_hd__inv_2
X_12383_ _12254_/Y _12380_/X _12374_/Y _12382_/X VGND VGND VPWR VPWR _12384_/A sky130_fd_sc_hd__a211o_4
X_24369_ _24641_/CLK _17278_/Y HRESETn VGND VGND VPWR VPWR _24369_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14122_ _25223_/Q _14106_/X _14108_/A _14108_/B VGND VGND VPWR VPWR _14122_/X sky130_fd_sc_hd__o22a_4
XFILLER_181_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25143__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14053_ _14053_/A VGND VGND VPWR VPWR _14054_/A sky130_fd_sc_hd__buf_2
X_18930_ _18929_/Y _18925_/X _17440_/X _18925_/A VGND VGND VPWR VPWR _18930_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22414__B1 _22946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13004_ _12970_/X _13002_/X _13003_/X VGND VGND VPWR VPWR _25364_/D sky130_fd_sc_hd__and3_4
XANTENNA__22702__B _21843_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18861_ _18861_/A _18861_/B _18859_/X _18861_/D VGND VGND VPWR VPWR _18861_/X sky130_fd_sc_hd__or4_4
XANTENNA__20503__A _20503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19830__B2 _19805_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_254_0_HCLK clkbuf_8_255_0_HCLK/A VGND VGND VPWR VPWR _25243_/CLK sky130_fd_sc_hd__clkbuf_1
X_17812_ _17757_/Y _17758_/Y _17833_/B VGND VGND VPWR VPWR _17813_/B sky130_fd_sc_hd__or3_4
XFILLER_121_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18792_ _18679_/Y _18789_/X VGND VGND VPWR VPWR _18792_/X sky130_fd_sc_hd__or2_4
XFILLER_121_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14955_ _15228_/A VGND VGND VPWR VPWR _15061_/A sky130_fd_sc_hd__inv_2
X_17743_ _24284_/Q VGND VGND VPWR VPWR _17743_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24864__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22193__A2 _22417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13906_ _13883_/Y _13901_/X _14239_/A VGND VGND VPWR VPWR _13954_/A sky130_fd_sc_hd__a21o_4
XFILLER_235_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14886_ _14886_/A VGND VGND VPWR VPWR _15182_/A sky130_fd_sc_hd__inv_2
X_17674_ _17577_/C _17676_/B _17673_/Y VGND VGND VPWR VPWR _24302_/D sky130_fd_sc_hd__o21a_4
XFILLER_208_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18617__A1_N _16619_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19413_ _19426_/A VGND VGND VPWR VPWR _19413_/X sky130_fd_sc_hd__buf_2
X_13837_ _25255_/Q VGND VGND VPWR VPWR _13837_/Y sky130_fd_sc_hd__inv_2
X_16625_ _14765_/A _14762_/C _16621_/X _13727_/A _16624_/X VGND VGND VPWR VPWR _24514_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_223_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19346__B1 _19279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16556_ _16554_/Y _16555_/X _16382_/X _16555_/X VGND VGND VPWR VPWR _24541_/D sky130_fd_sc_hd__a2bb2o_4
X_19344_ _19340_/Y _19343_/X _19301_/X _19343_/X VGND VGND VPWR VPWR _19344_/X sky130_fd_sc_hd__a2bb2o_4
X_13768_ _13768_/A VGND VGND VPWR VPWR _13768_/X sky130_fd_sc_hd__buf_2
XFILLER_204_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12719_ _12584_/X _12722_/A VGND VGND VPWR VPWR _12719_/X sky130_fd_sc_hd__or2_4
X_15507_ _15505_/Y _15506_/X HADDR[14] _15506_/X VGND VGND VPWR VPWR _15507_/X sky130_fd_sc_hd__a2bb2o_4
X_16487_ _24566_/Q VGND VGND VPWR VPWR _16487_/Y sky130_fd_sc_hd__inv_2
X_19275_ _19274_/X VGND VGND VPWR VPWR _19290_/A sky130_fd_sc_hd__inv_2
X_13699_ _13676_/A _13676_/B VGND VGND VPWR VPWR _13699_/Y sky130_fd_sc_hd__nand2_4
XFILLER_248_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15438_ _13931_/A _15432_/X _15427_/X _13914_/X _15433_/X VGND VGND VPWR VPWR _24971_/D
+ sky130_fd_sc_hd__a32o_4
X_18226_ _18098_/A _18224_/X _18225_/X VGND VGND VPWR VPWR _18227_/C sky130_fd_sc_hd__and3_4
X_15369_ _15369_/A _15369_/B VGND VGND VPWR VPWR _15370_/C sky130_fd_sc_hd__or2_4
X_18157_ _18125_/A _23845_/Q VGND VGND VPWR VPWR _18159_/B sky130_fd_sc_hd__or2_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12691__A _12569_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16163__A _21064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17108_ _17099_/C _17099_/D VGND VGND VPWR VPWR _17108_/Y sky130_fd_sc_hd__nand2_4
X_18088_ _18123_/A _18088_/B _18087_/X VGND VGND VPWR VPWR _18089_/C sky130_fd_sc_hd__and3_4
XANTENNA__15135__B2 _24595_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17039_ _17039_/A VGND VGND VPWR VPWR _17039_/Y sky130_fd_sc_hd__inv_2
X_20050_ _23523_/Q VGND VGND VPWR VPWR _20050_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21509__A _21178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22184__A2 _14245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23740_ _23747_/CLK _19429_/X VGND VGND VPWR VPWR _18175_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15536__A2_N _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24534__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _20953_/A VGND VGND VPWR VPWR _20952_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16399__B1 _16397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23671_ _23665_/CLK _23671_/D VGND VGND VPWR VPWR _13307_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _24048_/Q VGND VGND VPWR VPWR _20883_/Y sky130_fd_sc_hd__inv_2
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19337__B1 _19203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25410_ _25409_/CLK _25410_/D HRESETn VGND VGND VPWR VPWR _25410_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11770__A _13829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22622_ _24047_/Q _21303_/X _13120_/A _21317_/X VGND VGND VPWR VPWR _22622_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25341_ _25341_/CLK _25341_/D HRESETn VGND VGND VPWR VPWR _25341_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_210_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22553_ _22553_/A _22630_/B VGND VGND VPWR VPWR _22553_/X sky130_fd_sc_hd__or2_4
XFILLER_222_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21504_ _21504_/A _21278_/X VGND VGND VPWR VPWR _21504_/X sky130_fd_sc_hd__or2_4
X_25272_ _25272_/CLK _13795_/X HRESETn VGND VGND VPWR VPWR _25272_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22484_ _22298_/A _22484_/B VGND VGND VPWR VPWR _22498_/C sky130_fd_sc_hd__and2_4
XFILLER_6_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25393__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24223_ _23398_/CLK _24223_/D HRESETn VGND VGND VPWR VPWR _18268_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21435_ _21435_/A _23002_/A VGND VGND VPWR VPWR _21435_/X sky130_fd_sc_hd__or2_4
XFILLER_135_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22644__B1 _21832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16073__A _24716_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25322__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24154_ _24148_/CLK _24154_/D HRESETn VGND VGND VPWR VPWR _24154_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21366_ _14871_/Y _21365_/X _14227_/Y _14209_/X VGND VGND VPWR VPWR _21372_/B sky130_fd_sc_hd__o22a_4
XANTENNA__16323__B1 _16226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18401__A2_N _18400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23105_ _24810_/Q _23040_/X VGND VGND VPWR VPWR _23105_/X sky130_fd_sc_hd__or2_4
X_20317_ _21974_/A _20316_/X _15762_/X _20316_/X VGND VGND VPWR VPWR _23422_/D sky130_fd_sc_hd__a2bb2o_4
X_24085_ _25226_/CLK _20468_/X HRESETn VGND VGND VPWR VPWR _20444_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_104_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21297_ _21588_/A VGND VGND VPWR VPWR _21297_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22947__A1 _12813_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22522__B _22522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23036_ _23036_/A _22897_/X VGND VGND VPWR VPWR _23036_/X sky130_fd_sc_hd__or2_4
XFILLER_107_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20248_ _20243_/A VGND VGND VPWR VPWR _20248_/X sky130_fd_sc_hd__buf_2
XANTENNA__22411__A3 _22138_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20179_ _20178_/X VGND VGND VPWR VPWR _20180_/A sky130_fd_sc_hd__inv_2
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11664__B _11664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_HCLK_A clkbuf_3_4_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_21_0_HCLK clkbuf_8_21_0_HCLK/A VGND VGND VPWR VPWR _24377_/CLK sky130_fd_sc_hd__clkbuf_1
X_24987_ _24976_/CLK _15392_/X HRESETn VGND VGND VPWR VPWR _24987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_84_0_HCLK clkbuf_8_85_0_HCLK/A VGND VGND VPWR VPWR _25387_/CLK sky130_fd_sc_hd__clkbuf_1
X_14740_ _14739_/X VGND VGND VPWR VPWR _14740_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24275__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11952_ _11945_/Y _18902_/B _11951_/X VGND VGND VPWR VPWR _11952_/X sky130_fd_sc_hd__o21a_4
X_23938_ _23938_/CLK _20551_/Y HRESETn VGND VGND VPWR VPWR _18872_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21383__B1 _21177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24204__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14671_ _22069_/A _22367_/A VGND VGND VPWR VPWR _14671_/X sky130_fd_sc_hd__and2_4
X_11883_ _11883_/A VGND VGND VPWR VPWR _11883_/Y sky130_fd_sc_hd__inv_2
X_23869_ _23853_/CLK _23869_/D VGND VGND VPWR VPWR _19061_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_60_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19328__B1 _19282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16410_ _22701_/A VGND VGND VPWR VPWR _16410_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11680__A _22136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13622_ _13621_/Y _13586_/A VGND VGND VPWR VPWR _13622_/X sky130_fd_sc_hd__or2_4
XFILLER_199_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17390_ _20643_/A _20640_/A VGND VGND VPWR VPWR _20645_/A sky130_fd_sc_hd__or2_4
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16341_ _24619_/Q VGND VGND VPWR VPWR _16341_/Y sky130_fd_sc_hd__inv_2
X_13553_ _25085_/Q VGND VGND VPWR VPWR _14550_/A sky130_fd_sc_hd__inv_2
X_25539_ _25538_/CLK _25539_/D HRESETn VGND VGND VPWR VPWR _25539_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12504_ _25407_/Q _12502_/Y _12503_/Y _12515_/A VGND VGND VPWR VPWR _12507_/C sky130_fd_sc_hd__a2bb2o_4
X_19060_ _19059_/Y _19054_/X _18965_/X _19054_/X VGND VGND VPWR VPWR _23870_/D sky130_fd_sc_hd__a2bb2o_4
X_16272_ _22890_/B VGND VGND VPWR VPWR _16272_/X sky130_fd_sc_hd__buf_2
X_13484_ _13484_/A VGND VGND VPWR VPWR _13499_/A sky130_fd_sc_hd__inv_2
XFILLER_157_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15223_ _15203_/X _15223_/B _15222_/X VGND VGND VPWR VPWR _25025_/D sky130_fd_sc_hd__and3_4
X_18011_ _18057_/A VGND VGND VPWR VPWR _18053_/A sky130_fd_sc_hd__buf_2
XANTENNA__21438__A1 _16637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12435_ _12431_/X VGND VGND VPWR VPWR _12436_/B sky130_fd_sc_hd__inv_2
XANTENNA__21438__B2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25063__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15154_ _15148_/Y VGND VGND VPWR VPWR _15296_/A sky130_fd_sc_hd__buf_2
X_12366_ _12360_/Y VGND VGND VPWR VPWR _13097_/A sky130_fd_sc_hd__buf_2
XANTENNA__16314__B1 _15951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22713__A _22713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14105_ _14105_/A _14105_/B _14091_/A VGND VGND VPWR VPWR _14106_/B sky130_fd_sc_hd__or3_4
XFILLER_181_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15085_ _15085_/A VGND VGND VPWR VPWR _15085_/Y sky130_fd_sc_hd__inv_2
X_19962_ _19962_/A VGND VGND VPWR VPWR _19962_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12297_ _24847_/Q VGND VGND VPWR VPWR _12297_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14036_ _13990_/C VGND VGND VPWR VPWR _14038_/B sky130_fd_sc_hd__inv_2
X_18913_ _18925_/A VGND VGND VPWR VPWR _18913_/X sky130_fd_sc_hd__buf_2
XANTENNA__21329__A _21582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19893_ _19893_/A VGND VGND VPWR VPWR _19893_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18844_ _24560_/Q _24139_/Q _16503_/Y _18778_/A VGND VGND VPWR VPWR _18844_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18775_ _18694_/B _18774_/X VGND VGND VPWR VPWR _18778_/B sky130_fd_sc_hd__or2_4
X_15987_ _15983_/X _15986_/Y VGND VGND VPWR VPWR _15988_/A sky130_fd_sc_hd__and2_4
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17726_ _18279_/A _17726_/B VGND VGND VPWR VPWR _17726_/X sky130_fd_sc_hd__and2_4
X_14938_ _25025_/Q _14936_/Y _15261_/A _14940_/A VGND VGND VPWR VPWR _14946_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_180_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21064__A _21064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17657_ _17582_/B _17656_/X VGND VGND VPWR VPWR _17660_/B sky130_fd_sc_hd__or2_4
XANTENNA__16896__A2_N _16895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14869_ _14863_/Y _14805_/X _14806_/X _14868_/X VGND VGND VPWR VPWR _14869_/X sky130_fd_sc_hd__o22a_4
X_16608_ _24520_/Q VGND VGND VPWR VPWR _16608_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21999__A _13772_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17588_ _17587_/X VGND VGND VPWR VPWR _17589_/B sky130_fd_sc_hd__inv_2
XANTENNA__23998__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19327_ _19327_/A VGND VGND VPWR VPWR _19327_/X sky130_fd_sc_hd__buf_2
XANTENNA__15997__A _15988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16539_ _16539_/A VGND VGND VPWR VPWR _16792_/A sky130_fd_sc_hd__buf_2
XANTENNA__22874__B1 _24276_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23927__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19258_ _23800_/Q VGND VGND VPWR VPWR _22066_/B sky130_fd_sc_hd__inv_2
XANTENNA__16553__B1 _16467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18209_ _18113_/A _18209_/B VGND VGND VPWR VPWR _18209_/X sky130_fd_sc_hd__or2_4
X_19189_ _19188_/Y _19186_/X _19122_/X _19186_/X VGND VGND VPWR VPWR _23825_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14406__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13310__A _13433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21220_ _21220_/A _13769_/Y VGND VGND VPWR VPWR _21220_/X sky130_fd_sc_hd__and2_4
XFILLER_145_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21151_ _21151_/A _21150_/X VGND VGND VPWR VPWR _21151_/Y sky130_fd_sc_hd__nor2_4
XFILLER_160_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20102_ _20102_/A VGND VGND VPWR VPWR _20102_/X sky130_fd_sc_hd__buf_2
XFILLER_171_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21082_ _22523_/B VGND VGND VPWR VPWR _21082_/X sky130_fd_sc_hd__buf_2
XANTENNA__24786__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20143__A _20137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20033_ _20032_/X VGND VGND VPWR VPWR _20034_/A sky130_fd_sc_hd__inv_2
X_24910_ _24910_/CLK _24910_/D HRESETn VGND VGND VPWR VPWR _24910_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24715__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24841_ _24809_/CLK _24841_/D HRESETn VGND VGND VPWR VPWR _12296_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_74_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24772_ _24766_/CLK _15940_/X HRESETn VGND VGND VPWR VPWR _24772_/Q sky130_fd_sc_hd__dfrtp_4
X_21984_ _22400_/A _22266_/A _22003_/A _21984_/D VGND VGND VPWR VPWR _21984_/X sky130_fd_sc_hd__or4_4
XPHY_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23723_ _23691_/CLK _23723_/D VGND VGND VPWR VPWR _23723_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _24060_/Q VGND VGND VPWR VPWR _20935_/Y sky130_fd_sc_hd__inv_2
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _23665_/CLK _19683_/X VGND VGND VPWR VPWR _13340_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _24044_/Q VGND VGND VPWR VPWR _20866_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22605_ _16689_/Y _22641_/B VGND VGND VPWR VPWR _22605_/X sky130_fd_sc_hd__and2_4
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23585_ _23559_/CLK _23585_/D VGND VGND VPWR VPWR _19881_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20797_ _20796_/A _20793_/A _20793_/B VGND VGND VPWR VPWR _20797_/X sky130_fd_sc_hd__or3_4
XANTENNA__18283__A _17704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25503__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25324_ _23887_/CLK _13465_/X HRESETn VGND VGND VPWR VPWR _25324_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22517__B _22696_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22536_ _22535_/X VGND VGND VPWR VPWR _22536_/X sky130_fd_sc_hd__buf_2
XFILLER_194_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15898__A2 _15887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25255_ _25260_/CLK _13838_/X HRESETn VGND VGND VPWR VPWR _25255_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22467_ _20862_/C _23129_/A _16696_/Y _22279_/X VGND VGND VPWR VPWR _22468_/B sky130_fd_sc_hd__o22a_4
XFILLER_167_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12220_ _22150_/A VGND VGND VPWR VPWR _12220_/Y sky130_fd_sc_hd__inv_2
X_24206_ _23391_/CLK _18343_/X HRESETn VGND VGND VPWR VPWR _13284_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13220__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21418_ _21418_/A VGND VGND VPWR VPWR _21418_/Y sky130_fd_sc_hd__inv_2
X_25186_ _25249_/CLK _14263_/X HRESETn VGND VGND VPWR VPWR _25186_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18836__A2 _24142_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22398_ _22395_/Y _22396_/X _22397_/X _13544_/A _22051_/X VGND VGND VPWR VPWR _22399_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_136_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12151_ _12149_/X _12150_/Y VGND VGND VPWR VPWR _12151_/X sky130_fd_sc_hd__and2_4
X_24137_ _24139_/CLK _18793_/X HRESETn VGND VGND VPWR VPWR _24137_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21840__A1 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12581__B2 _24885_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21349_ _21349_/A VGND VGND VPWR VPWR _21364_/B sky130_fd_sc_hd__inv_2
XANTENNA__21840__B2 _21839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12082_ _12082_/A VGND VGND VPWR VPWR _13483_/A sky130_fd_sc_hd__buf_2
X_24068_ _25346_/CLK _24068_/D HRESETn VGND VGND VPWR VPWR _24068_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17346__B _17366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23042__B1 _24878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23067__C _23066_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11675__A _16446_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19797__B1 _19708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15910_ _15910_/A VGND VGND VPWR VPWR _15910_/Y sky130_fd_sc_hd__inv_2
X_23019_ _16663_/Y _22829_/X _15578_/Y _22832_/X VGND VGND VPWR VPWR _23019_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24456__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16890_ _22191_/A _16889_/Y _16096_/Y _24285_/Q VGND VGND VPWR VPWR _16890_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23364__A _23364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15841_ _15670_/X _15836_/B VGND VGND VPWR VPWR _15841_/X sky130_fd_sc_hd__or2_4
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16989__A1_N _24733_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22148__A2 _22282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18560_ _18560_/A _18477_/D VGND VGND VPWR VPWR _18587_/B sky130_fd_sc_hd__or2_4
XFILLER_58_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12984_ _12984_/A _12981_/X _12983_/X VGND VGND VPWR VPWR _12984_/X sky130_fd_sc_hd__or3_4
X_15772_ _15544_/Y _15642_/X _15770_/X _21017_/B _15771_/X VGND VGND VPWR VPWR _15772_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_76_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17511_ _24315_/Q VGND VGND VPWR VPWR _17511_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11935_ _11948_/B _17442_/B VGND VGND VPWR VPWR _11935_/X sky130_fd_sc_hd__or2_4
X_14723_ _14722_/Y _14701_/Y _22043_/A _14701_/A VGND VGND VPWR VPWR _14735_/B sky130_fd_sc_hd__o22a_4
X_18491_ _18491_/A VGND VGND VPWR VPWR _18491_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14654_ _14654_/A VGND VGND VPWR VPWR _14654_/X sky130_fd_sc_hd__buf_2
X_17442_ _11947_/A _17442_/B VGND VGND VPWR VPWR _18902_/D sky130_fd_sc_hd__or2_4
X_11866_ _11802_/Y _11860_/Y VGND VGND VPWR VPWR _11866_/X sky130_fd_sc_hd__and2_4
XFILLER_178_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21108__B1 _21047_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13605_ _13600_/A VGND VGND VPWR VPWR _13606_/B sky130_fd_sc_hd__inv_2
XPHY_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14585_ _14548_/Y _14554_/X VGND VGND VPWR VPWR _14585_/Y sky130_fd_sc_hd__nand2_4
X_17373_ _17203_/X _17344_/B VGND VGND VPWR VPWR _17374_/B sky130_fd_sc_hd__or2_4
XPHY_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11797_ _11797_/A VGND VGND VPWR VPWR _11797_/Y sky130_fd_sc_hd__inv_2
XPHY_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19112_ _19111_/Y _19109_/X _19067_/X _19109_/X VGND VGND VPWR VPWR _19112_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22427__B _22409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13536_ _13536_/A VGND VGND VPWR VPWR _13536_/Y sky130_fd_sc_hd__inv_2
X_16324_ _22710_/A VGND VGND VPWR VPWR _16324_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16535__B1 _16358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16927__A1_N _16133_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16255_ _16254_/Y _16252_/X _16062_/X _16252_/X VGND VGND VPWR VPWR _24652_/D sky130_fd_sc_hd__a2bb2o_4
X_19043_ _19042_/Y _19040_/X _18951_/X _19040_/X VGND VGND VPWR VPWR _19043_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22608__B1 _21832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13467_ _13466_/Y _13464_/X _11765_/X _13464_/X VGND VGND VPWR VPWR _25323_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15206_ _15062_/X _15214_/D VGND VGND VPWR VPWR _15207_/B sky130_fd_sc_hd__or2_4
X_12418_ _12418_/A _12418_/B _12271_/X _12370_/X VGND VGND VPWR VPWR _12418_/X sky130_fd_sc_hd__or4_4
X_16186_ _16177_/Y _16185_/X _15991_/X _16185_/X VGND VGND VPWR VPWR _16186_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13398_ _13252_/A _18927_/A VGND VGND VPWR VPWR _13400_/B sky130_fd_sc_hd__or2_4
XFILLER_127_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15137_ _24998_/Q VGND VGND VPWR VPWR _15137_/Y sky130_fd_sc_hd__inv_2
X_12349_ _25357_/Q VGND VGND VPWR VPWR _12349_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16441__A _18560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21831__B2 _11706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15068_ _24987_/Q VGND VGND VPWR VPWR _15068_/Y sky130_fd_sc_hd__inv_2
X_19945_ _19945_/A VGND VGND VPWR VPWR _19945_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21059__A _21059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14313__A2 _25170_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14019_ _14017_/Y _14018_/X _14019_/C _14019_/D VGND VGND VPWR VPWR _14020_/A sky130_fd_sc_hd__or4_4
XANTENNA__24197__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19876_ _19876_/A VGND VGND VPWR VPWR _19876_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24126__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18827_ _16498_/Y _18769_/A _16498_/Y _18769_/A VGND VGND VPWR VPWR _18830_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23274__A _23251_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18758_ _18692_/Y _18746_/X VGND VGND VPWR VPWR _18758_/X sky130_fd_sc_hd__or2_4
XFILLER_215_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17703__C _21177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17709_ _17709_/A VGND VGND VPWR VPWR _21475_/A sky130_fd_sc_hd__buf_2
XFILLER_209_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18689_ _18689_/A VGND VGND VPWR VPWR _18689_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20720_ _15615_/Y _20708_/X _20716_/X _20719_/Y VGND VGND VPWR VPWR _20720_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22618__A _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20651_ _20651_/A VGND VGND VPWR VPWR _20651_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22847__B1 _12329_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22311__A2 _21325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19712__B1 _19711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23370_ _21017_/X VGND VGND VPWR VPWR IRQ[26] sky130_fd_sc_hd__buf_2
X_20582_ _14414_/Y _20566_/X _20556_/X _20581_/X VGND VGND VPWR VPWR _20583_/A sky130_fd_sc_hd__a211o_4
XFILLER_139_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16526__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20138__A _20137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22321_ _17346_/A _22429_/A _12197_/A _21075_/Y VGND VGND VPWR VPWR _22321_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25040_ _25015_/CLK _15052_/Y HRESETn VGND VGND VPWR VPWR pwm_S6 sky130_fd_sc_hd__dfrtp_4
XFILLER_180_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22252_ _22255_/A _19993_/Y VGND VGND VPWR VPWR _22252_/X sky130_fd_sc_hd__or2_4
XFILLER_118_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24967__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22353__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21203_ _21199_/X _21202_/X _22257_/A VGND VGND VPWR VPWR _21203_/X sky130_fd_sc_hd__o21a_4
XFILLER_145_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22183_ _22183_/A VGND VGND VPWR VPWR _22183_/Y sky130_fd_sc_hd__inv_2
X_21134_ _21159_/A VGND VGND VPWR VPWR _21346_/A sky130_fd_sc_hd__inv_2
XANTENNA__23024__B1 _22098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21065_ _15661_/A VGND VGND VPWR VPWR _21736_/A sky130_fd_sc_hd__buf_2
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20016_ _22262_/B _20013_/X _19967_/X _20013_/X VGND VGND VPWR VPWR _23537_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20601__A _20601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23327__B2 _21315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24824_ _24855_/CLK _24824_/D HRESETn VGND VGND VPWR VPWR _24824_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12079__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12618__A2 _12626_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24755_ _25369_/CLK _24755_/D HRESETn VGND VGND VPWR VPWR _22410_/A sky130_fd_sc_hd__dfrtp_4
X_21967_ _21968_/A _19585_/X _14602_/Y _23685_/Q VGND VGND VPWR VPWR _21967_/X sky130_fd_sc_hd__o22a_4
XFILLER_27_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _25537_/Q VGND VGND VPWR VPWR _11720_/Y sky130_fd_sc_hd__inv_2
X_23706_ _23706_/CLK _19527_/X VGND VGND VPWR VPWR _23706_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13215__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22550__A2 _21098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ _20892_/X _20917_/Y _24499_/Q _20896_/X VGND VGND VPWR VPWR _24055_/D sky130_fd_sc_hd__a2bb2o_4
X_24686_ _24686_/CLK _24686_/D HRESETn VGND VGND VPWR VPWR _22153_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_54_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ _22386_/A _21898_/B VGND VGND VPWR VPWR _21899_/C sky130_fd_sc_hd__or2_4
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_158_0_HCLK clkbuf_7_79_0_HCLK/X VGND VGND VPWR VPWR _25109_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21432__A _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _14664_/A VGND VGND VPWR VPWR _11651_/Y sky130_fd_sc_hd__inv_2
X_23637_ _23644_/CLK _23637_/D VGND VGND VPWR VPWR _13379_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ _16703_/Y _20846_/X _20834_/X _20848_/X VGND VGND VPWR VPWR _20850_/A sky130_fd_sc_hd__o22a_4
XFILLER_120_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19703__B1 _19702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _14096_/A _14370_/B VGND VGND VPWR VPWR _14370_/Y sky130_fd_sc_hd__nor2_4
XFILLER_23_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23568_ _25070_/CLK _19926_/X VGND VGND VPWR VPWR _19924_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_211_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _11951_/X _13302_/X _13320_/X _25331_/Q _13243_/X VGND VGND VPWR VPWR _13321_/X
+ sky130_fd_sc_hd__o32a_4
X_25307_ _25466_/CLK _25307_/D HRESETn VGND VGND VPWR VPWR _13503_/A sky130_fd_sc_hd__dfrtp_4
X_22519_ _21178_/A _13771_/A _21377_/X VGND VGND VPWR VPWR _22520_/A sky130_fd_sc_hd__or3_4
XFILLER_10_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23499_ _23499_/CLK _20112_/X VGND VGND VPWR VPWR _23499_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16040_ _16040_/A VGND VGND VPWR VPWR _16040_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13252_ _13252_/A _23816_/Q VGND VGND VPWR VPWR _13254_/B sky130_fd_sc_hd__or2_4
X_25238_ _25238_/CLK _14064_/X HRESETn VGND VGND VPWR VPWR _13978_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_129_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12203_ _12201_/A _22898_/A _12201_/Y _12202_/Y VGND VGND VPWR VPWR _12203_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12554__B2 _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13183_ _11970_/Y _13182_/Y _11962_/A VGND VGND VPWR VPWR _13184_/A sky130_fd_sc_hd__o21a_4
X_25169_ _25164_/CLK _25169_/D HRESETn VGND VGND VPWR VPWR _25169_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24637__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23078__B _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12134_ _12119_/A _12119_/B _12119_/Y _12133_/X VGND VGND VPWR VPWR _12145_/A sky130_fd_sc_hd__a211o_4
XFILLER_97_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17991_ _17999_/A VGND VGND VPWR VPWR _18182_/A sky130_fd_sc_hd__buf_2
XFILLER_145_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19730_ _13379_/B VGND VGND VPWR VPWR _19730_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24290__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12065_ _12060_/A VGND VGND VPWR VPWR _12065_/X sky130_fd_sc_hd__buf_2
X_16942_ _16942_/A _16937_/X _16942_/C _16942_/D VGND VGND VPWR VPWR _16949_/C sky130_fd_sc_hd__or4_4
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23030__A3 _22849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22710__B _21864_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19661_ _13339_/B VGND VGND VPWR VPWR _19661_/Y sky130_fd_sc_hd__inv_2
X_16873_ _16867_/X VGND VGND VPWR VPWR _16873_/X sky130_fd_sc_hd__buf_2
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18612_ _24147_/Q VGND VGND VPWR VPWR _18613_/A sky130_fd_sc_hd__inv_2
X_15824_ _12306_/Y _15820_/X _15754_/X _15823_/X VGND VGND VPWR VPWR _24828_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19592_ _19592_/A VGND VGND VPWR VPWR _19592_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25496__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18543_ _18523_/X _18540_/B _18542_/Y VGND VGND VPWR VPWR _18543_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_54_0_HCLK clkbuf_7_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12967_ _12967_/A _12958_/B _12967_/C VGND VGND VPWR VPWR _25368_/D sky130_fd_sc_hd__and3_4
X_15755_ _15759_/A VGND VGND VPWR VPWR _15755_/X sky130_fd_sc_hd__buf_2
XFILLER_206_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11918_ _19617_/A VGND VGND VPWR VPWR _11918_/Y sky130_fd_sc_hd__inv_2
X_14706_ _14706_/A VGND VGND VPWR VPWR _22205_/A sky130_fd_sc_hd__buf_2
XFILLER_205_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18474_ _18589_/A _18420_/Y _18473_/Y _18400_/Y VGND VGND VPWR VPWR _18478_/B sky130_fd_sc_hd__or4_4
X_12898_ _12813_/Y _12892_/X _12862_/X _12894_/Y VGND VGND VPWR VPWR _12899_/A sky130_fd_sc_hd__a211o_4
X_15686_ _15686_/A _15686_/B VGND VGND VPWR VPWR _15687_/A sky130_fd_sc_hd__or2_4
XFILLER_221_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16756__B1 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17425_ _17424_/Y _17422_/X _16778_/X _17422_/X VGND VGND VPWR VPWR _24330_/D sky130_fd_sc_hd__a2bb2o_4
X_11849_ _11849_/A _11849_/B VGND VGND VPWR VPWR _11856_/B sky130_fd_sc_hd__and2_4
X_14637_ _18123_/A VGND VGND VPWR VPWR _17942_/A sky130_fd_sc_hd__buf_2
XFILLER_221_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14568_ _14563_/A _14563_/B VGND VGND VPWR VPWR _14569_/A sky130_fd_sc_hd__and2_4
X_17356_ _17358_/B VGND VGND VPWR VPWR _17357_/B sky130_fd_sc_hd__inv_2
XANTENNA__13779__B _14243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16307_ _16305_/Y _16306_/X _16020_/X _16306_/X VGND VGND VPWR VPWR _16307_/X sky130_fd_sc_hd__a2bb2o_4
X_13519_ _13462_/C _13456_/X _12160_/C _13483_/A VGND VGND VPWR VPWR _13520_/A sky130_fd_sc_hd__or4_4
XFILLER_147_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19747__A _19740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14499_ _23958_/Q VGND VGND VPWR VPWR _14499_/X sky130_fd_sc_hd__buf_2
X_17287_ _17286_/X VGND VGND VPWR VPWR _24367_/D sky130_fd_sc_hd__inv_2
XFILLER_174_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19026_ _19341_/A _19163_/B _19026_/C _19026_/D VGND VGND VPWR VPWR _19026_/X sky130_fd_sc_hd__and4_4
X_16238_ _22590_/A VGND VGND VPWR VPWR _16238_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23254__B1 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24378__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16169_ _16166_/X VGND VGND VPWR VPWR _16170_/B sky130_fd_sc_hd__buf_2
XFILLER_114_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24307__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15495__B1 HADDR[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19928_ _19927_/Y _19925_/X _19610_/X _19925_/X VGND VGND VPWR VPWR _19928_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12204__A _12204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22620__B _22696_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19859_ _19859_/A VGND VGND VPWR VPWR _19859_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22870_ _22870_/A _22909_/B VGND VGND VPWR VPWR _22870_/X sky130_fd_sc_hd__or2_4
X_21821_ _21805_/X _21820_/X _21501_/X VGND VGND VPWR VPWR _21821_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_237_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23942__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19933__B1 _19617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24540_ _24540_/CLK _24540_/D HRESETn VGND VGND VPWR VPWR _16557_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_221_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21752_ _21775_/A _21752_/B VGND VGND VPWR VPWR _21754_/B sky130_fd_sc_hd__or2_4
XFILLER_240_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16747__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21740__B1 _21582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20703_ _20702_/X VGND VGND VPWR VPWR _24006_/D sky130_fd_sc_hd__inv_2
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24471_ _25021_/CLK _16738_/X HRESETn VGND VGND VPWR VPWR _16737_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21683_ _21657_/A _21683_/B VGND VGND VPWR VPWR _21685_/B sky130_fd_sc_hd__or2_4
XFILLER_197_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12874__A _12804_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16346__A _24617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23422_ _23425_/CLK _23422_/D VGND VGND VPWR VPWR _21984_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_196_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20634_ _17388_/A _17388_/B VGND VGND VPWR VPWR _20634_/Y sky130_fd_sc_hd__nand2_4
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23353_ VGND VGND VPWR VPWR _23353_/HI IRQ[29] sky130_fd_sc_hd__conb_1
X_20565_ _20565_/A VGND VGND VPWR VPWR _23941_/D sky130_fd_sc_hd__inv_2
XFILLER_164_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22304_ _22195_/X _22272_/Y _22285_/Y _22304_/D VGND VGND VPWR VPWR HRDATA[6] sky130_fd_sc_hd__or4_4
XFILLER_192_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23284_ _24711_/Q _23156_/X VGND VGND VPWR VPWR _23284_/X sky130_fd_sc_hd__or2_4
XFILLER_166_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15722__A1 _15540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20496_ _20496_/A _20486_/Y _24076_/Q VGND VGND VPWR VPWR _20497_/B sky130_fd_sc_hd__and3_4
XFILLER_180_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25023_ _25028_/CLK _25023_/D HRESETn VGND VGND VPWR VPWR _15228_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_118_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22235_ _22251_/A _22235_/B VGND VGND VPWR VPWR _22235_/X sky130_fd_sc_hd__or2_4
XANTENNA__11712__A1_N _11710_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24730__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18267__A3 _18257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24048__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22166_ _21845_/A _22163_/X _22166_/C VGND VGND VPWR VPWR _22195_/B sky130_fd_sc_hd__and3_4
XFILLER_133_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21117_ _13110_/B VGND VGND VPWR VPWR _21117_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19392__A _18981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22097_ _22097_/A _23088_/B VGND VGND VPWR VPWR _22097_/X sky130_fd_sc_hd__or2_4
XFILLER_120_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21048_ _21128_/B VGND VGND VPWR VPWR _21048_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21427__A _21427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13870_ _13860_/X _13869_/X _25186_/Q _13845_/Y VGND VGND VPWR VPWR _13870_/X sky130_fd_sc_hd__o22a_4
XFILLER_247_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12821_ _25374_/Q VGND VGND VPWR VPWR _12948_/A sky130_fd_sc_hd__inv_2
XFILLER_74_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24807_ _24804_/CLK _24807_/D HRESETn VGND VGND VPWR VPWR _24807_/Q sky130_fd_sc_hd__dfrtp_4
X_22999_ _23209_/A _22996_/X _22998_/X VGND VGND VPWR VPWR _23006_/C sky130_fd_sc_hd__and3_4
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12752_ _25386_/Q VGND VGND VPWR VPWR _12838_/A sky130_fd_sc_hd__inv_2
X_15540_ _15724_/A VGND VGND VPWR VPWR _15540_/X sky130_fd_sc_hd__buf_2
XFILLER_199_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24738_ _24737_/CLK _24738_/D HRESETn VGND VGND VPWR VPWR _24738_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16738__B1 _15721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _15981_/A VGND VGND VPWR VPWR _11704_/A sky130_fd_sc_hd__buf_2
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _15458_/A VGND VGND VPWR VPWR _15471_/X sky130_fd_sc_hd__buf_2
X_12683_ _12682_/X VGND VGND VPWR VPWR _12684_/B sky130_fd_sc_hd__inv_2
X_24669_ _24675_/CLK _16208_/X HRESETn VGND VGND VPWR VPWR _16207_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14422_/A VGND VGND VPWR VPWR _21365_/A sky130_fd_sc_hd__buf_2
X_17210_ _16300_/Y _17298_/A _16300_/Y _17298_/A VGND VGND VPWR VPWR _17210_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18190_ _18126_/A _19158_/A VGND VGND VPWR VPWR _18190_/X sky130_fd_sc_hd__or2_4
XANTENNA__24889__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14353_ _25158_/Q _14340_/X _25157_/Q _14345_/X VGND VGND VPWR VPWR _14353_/X sky130_fd_sc_hd__o22a_4
X_17141_ _16975_/Y _17128_/X VGND VGND VPWR VPWR _17141_/Y sky130_fd_sc_hd__nand2_4
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24818__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13304_ _13443_/A _13304_/B VGND VGND VPWR VPWR _13304_/X sky130_fd_sc_hd__or2_4
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17072_ _17381_/B _17072_/B _17071_/X VGND VGND VPWR VPWR _17073_/A sky130_fd_sc_hd__or3_4
XFILLER_10_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22039__A1 _21954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14284_ _14288_/A VGND VGND VPWR VPWR _14296_/A sky130_fd_sc_hd__buf_2
XFILLER_115_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13235_ _13234_/X _13235_/B VGND VGND VPWR VPWR _13235_/X sky130_fd_sc_hd__or2_4
X_16023_ _16022_/Y _16019_/X _15946_/X _16019_/X VGND VGND VPWR VPWR _16023_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24471__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18258__A3 _18257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16269__A2 _15986_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24400__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13166_ _13385_/A VGND VGND VPWR VPWR _13353_/A sky130_fd_sc_hd__buf_2
XFILLER_3_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18663__B1 _24516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12117_ _12116_/X VGND VGND VPWR VPWR _12117_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13097_ _13097_/A _13097_/B VGND VGND VPWR VPWR _13098_/B sky130_fd_sc_hd__or2_4
X_17974_ _18090_/A VGND VGND VPWR VPWR _17981_/A sky130_fd_sc_hd__buf_2
XFILLER_69_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16618__A2_N _16541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19713_ _13442_/B VGND VGND VPWR VPWR _19713_/Y sky130_fd_sc_hd__inv_2
X_12048_ _12032_/Y _12047_/Y _11793_/X _12047_/Y VGND VGND VPWR VPWR _25487_/D sky130_fd_sc_hd__a2bb2o_4
X_16925_ _16925_/A VGND VGND VPWR VPWR _16925_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19644_ _19643_/Y _19641_/X _19543_/X _19641_/X VGND VGND VPWR VPWR _19644_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16856_ _14777_/X VGND VGND VPWR VPWR _16856_/X sky130_fd_sc_hd__buf_2
XANTENNA__16790__A1_N _16789_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15807_ _12303_/Y _15803_/X _11715_/X _15806_/X VGND VGND VPWR VPWR _24839_/D sky130_fd_sc_hd__a2bb2o_4
X_19575_ _19575_/A VGND VGND VPWR VPWR _19576_/A sky130_fd_sc_hd__buf_2
XFILLER_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16787_ _18951_/A VGND VGND VPWR VPWR _16787_/X sky130_fd_sc_hd__buf_2
X_13999_ _13995_/A _13990_/C _13999_/C VGND VGND VPWR VPWR _13999_/X sky130_fd_sc_hd__or3_4
X_18526_ _18442_/Y _18526_/B VGND VGND VPWR VPWR _18526_/X sky130_fd_sc_hd__or2_4
X_15738_ _15699_/Y VGND VGND VPWR VPWR _15738_/X sky130_fd_sc_hd__buf_2
XFILLER_18_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18457_ _24188_/Q VGND VGND VPWR VPWR _18457_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15669_ _22890_/B VGND VGND VPWR VPWR _16368_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_141_0_HCLK clkbuf_7_70_0_HCLK/X VGND VGND VPWR VPWR _23853_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_221_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17408_ _24074_/Q _13956_/Y _24334_/Q _13956_/A VGND VGND VPWR VPWR _24334_/D sky130_fd_sc_hd__o22a_4
X_18388_ _24192_/Q VGND VGND VPWR VPWR _18388_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17339_ _17246_/Y _17333_/X _17284_/X _17335_/Y VGND VGND VPWR VPWR _17340_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24559__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20350_ _20349_/Y VGND VGND VPWR VPWR _20350_/X sky130_fd_sc_hd__buf_2
XFILLER_174_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19009_ _19008_/Y _19004_/X _18981_/X _19004_/X VGND VGND VPWR VPWR _19009_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12518__B2 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20281_ _23435_/Q VGND VGND VPWR VPWR _20281_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22020_ _22020_/A _22020_/B VGND VGND VPWR VPWR _22020_/X sky130_fd_sc_hd__or2_4
XANTENNA__20056__A3 _11760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24141__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14140__B1 _25138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23971_ _24340_/CLK _21001_/X HRESETn VGND VGND VPWR VPWR _14790_/A sky130_fd_sc_hd__dfstp_4
XFILLER_229_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11773__A HWDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25347__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22922_ _22922_/A _22989_/B VGND VGND VPWR VPWR _22922_/X sky130_fd_sc_hd__and2_4
XFILLER_216_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22853_ _22853_/A VGND VGND VPWR VPWR _22853_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21804_ _21800_/X _21803_/X _18301_/X VGND VGND VPWR VPWR _21805_/C sky130_fd_sc_hd__o21a_4
X_22784_ _22782_/X _22784_/B _22876_/C VGND VGND VPWR VPWR _22784_/X sky130_fd_sc_hd__or3_4
XFILLER_225_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22078__A _21622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24523_ _24539_/CLK _16602_/X HRESETn VGND VGND VPWR VPWR _16600_/A sky130_fd_sc_hd__dfrtp_4
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21735_ _21556_/Y _21728_/X _21730_/X _21734_/Y VGND VGND VPWR VPWR _21735_/X sky130_fd_sc_hd__a211o_4
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24454_ _24073_/CLK _16771_/X HRESETn VGND VGND VPWR VPWR _24454_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12206__B1 _12204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21666_ _21475_/A _21666_/B _21665_/X VGND VGND VPWR VPWR _21666_/X sky130_fd_sc_hd__and3_4
XANTENNA__24982__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23405_ _23437_/CLK _23405_/D VGND VGND VPWR VPWR _20359_/A sky130_fd_sc_hd__dfxtp_4
X_20617_ _14863_/Y _20615_/X _20672_/A _20616_/X VGND VGND VPWR VPWR _20618_/A sky130_fd_sc_hd__a211o_4
X_24385_ _24377_/CLK _24385_/D HRESETn VGND VGND VPWR VPWR _17034_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24911__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21597_ _21597_/A VGND VGND VPWR VPWR _21597_/X sky130_fd_sc_hd__buf_2
XFILLER_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22525__B _21748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23336_ _23213_/A _23333_/X _23336_/C VGND VGND VPWR VPWR _23337_/D sky130_fd_sc_hd__and3_4
XANTENNA__24229__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20548_ _18886_/X VGND VGND VPWR VPWR _20553_/C sky130_fd_sc_hd__buf_2
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23267_ _12205_/Y _22718_/X _22719_/X _12316_/Y _22846_/X VGND VGND VPWR VPWR _23267_/X
+ sky130_fd_sc_hd__o32a_4
X_20479_ _20479_/A _20479_/B VGND VGND VPWR VPWR _20525_/C sky130_fd_sc_hd__or2_4
XFILLER_152_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13020_ _12287_/Y _13018_/X _13019_/X VGND VGND VPWR VPWR _13020_/Y sky130_fd_sc_hd__a21oi_4
X_25006_ _25204_/CLK _15314_/Y HRESETn VGND VGND VPWR VPWR _15150_/A sky130_fd_sc_hd__dfrtp_4
X_22218_ _22210_/A _22218_/B VGND VGND VPWR VPWR _22219_/C sky130_fd_sc_hd__or2_4
XFILLER_133_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18645__B1 _16589_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23198_ _17175_/Y _22485_/X _12735_/A _22444_/X VGND VGND VPWR VPWR _23198_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15459__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13585__D _13584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22149_ _22840_/A VGND VGND VPWR VPWR _22149_/X sky130_fd_sc_hd__buf_2
XFILLER_86_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14971_ _14970_/Y _16847_/A _25009_/Q _14939_/Y VGND VGND VPWR VPWR _14978_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20061__A _11785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23075__C _23075_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20204__B1 _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16710_ _16708_/Y _16704_/X _16353_/X _16709_/X VGND VGND VPWR VPWR _16710_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11683__A _11682_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25088__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13922_ _13922_/A VGND VGND VPWR VPWR _13927_/B sky130_fd_sc_hd__buf_2
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19070__B1 _18998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17690_ _17690_/A VGND VGND VPWR VPWR _24295_/D sky130_fd_sc_hd__inv_2
XANTENNA__16959__B1 _16009_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25017__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16641_ _16660_/A VGND VGND VPWR VPWR _16692_/A sky130_fd_sc_hd__buf_2
XFILLER_207_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13853_ _20476_/B _13850_/X _13851_/Y _13852_/X VGND VGND VPWR VPWR _13853_/X sky130_fd_sc_hd__o22a_4
XFILLER_223_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15631__B1 _15472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12804_ _25390_/Q VGND VGND VPWR VPWR _12804_/Y sky130_fd_sc_hd__inv_2
X_19360_ _19360_/A VGND VGND VPWR VPWR _19360_/X sky130_fd_sc_hd__buf_2
X_16572_ _16548_/A VGND VGND VPWR VPWR _16572_/X sky130_fd_sc_hd__buf_2
XANTENNA__12445__B1 _12390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13784_ _13792_/A VGND VGND VPWR VPWR _13784_/X sky130_fd_sc_hd__buf_2
XFILLER_16_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18311_ _22262_/A VGND VGND VPWR VPWR _21665_/A sky130_fd_sc_hd__buf_2
XFILLER_204_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15523_ _21133_/A VGND VGND VPWR VPWR _15523_/Y sky130_fd_sc_hd__inv_2
X_12735_ _12735_/A VGND VGND VPWR VPWR _12735_/Y sky130_fd_sc_hd__inv_2
X_19291_ _19289_/Y _19290_/X _19200_/X _19290_/X VGND VGND VPWR VPWR _19291_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18242_ _18238_/X _18240_/X _16229_/A _22696_/A _18241_/X VGND VGND VPWR VPWR _24240_/D
+ sky130_fd_sc_hd__a32o_4
X_12666_ _12597_/A _12670_/B _12665_/Y VGND VGND VPWR VPWR _12666_/X sky130_fd_sc_hd__o21a_4
X_15454_ _14232_/C _15451_/X _15426_/X _13902_/A _15436_/B VGND VGND VPWR VPWR _15454_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_214_0_HCLK clkbuf_8_214_0_HCLK/A VGND VGND VPWR VPWR _24460_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22716__A _22716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ _20592_/A VGND VGND VPWR VPWR _14405_/Y sky130_fd_sc_hd__inv_2
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18832__A1_N _16536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18173_ _18044_/A _18173_/B _18172_/X VGND VGND VPWR VPWR _18173_/X sky130_fd_sc_hd__or3_4
XANTENNA__24652__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12597_/A _12664_/C _12564_/Y _12555_/Y VGND VGND VPWR VPWR _12598_/C sky130_fd_sc_hd__or4_4
X_15385_ _15298_/A _15384_/X VGND VGND VPWR VPWR _15385_/X sky130_fd_sc_hd__or2_4
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ _17020_/Y _17040_/Y VGND VGND VPWR VPWR _17124_/X sky130_fd_sc_hd__or2_4
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14336_ _14329_/A _14339_/B _14335_/Y VGND VGND VPWR VPWR _25164_/D sky130_fd_sc_hd__o21a_4
XFILLER_116_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14267_ _14266_/Y VGND VGND VPWR VPWR _15451_/A sky130_fd_sc_hd__buf_2
X_17055_ _17054_/X VGND VGND VPWR VPWR _24403_/D sky130_fd_sc_hd__inv_2
XFILLER_116_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18847__A1_N _24552_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13218_ _13187_/A VGND VGND VPWR VPWR _13345_/A sky130_fd_sc_hd__buf_2
X_16006_ _16006_/A VGND VGND VPWR VPWR _16006_/Y sky130_fd_sc_hd__inv_2
X_14198_ _25205_/Q VGND VGND VPWR VPWR _14198_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22451__A _22451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13149_ _13187_/A VGND VGND VPWR VPWR _13433_/A sky130_fd_sc_hd__inv_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17957_ _17942_/A _17955_/X _17956_/X VGND VGND VPWR VPWR _17957_/X sky130_fd_sc_hd__and3_4
XFILLER_39_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16908_ _24265_/Q VGND VGND VPWR VPWR _16908_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17888_ _21059_/A _17625_/A VGND VGND VPWR VPWR _17889_/C sky130_fd_sc_hd__or2_4
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19627_ _19641_/A VGND VGND VPWR VPWR _19627_/X sky130_fd_sc_hd__buf_2
XFILLER_66_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16839_ _14911_/Y _16837_/X _16601_/X _16837_/X VGND VGND VPWR VPWR _16839_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19558_ _21950_/B _19555_/X _11915_/X _19555_/X VGND VGND VPWR VPWR _23695_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_24_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_24_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18509_ _18509_/A VGND VGND VPWR VPWR _18509_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19489_ _23719_/Q VGND VGND VPWR VPWR _21919_/B sky130_fd_sc_hd__inv_2
XANTENNA__17375__B1 _17268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21520_ _21843_/B VGND VGND VPWR VPWR _21520_/X sky130_fd_sc_hd__buf_2
XFILLER_210_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21530__A _22716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18823__B _18823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21451_ _23328_/A _21430_/Y _21444_/Y _21445_/X _21450_/X VGND VGND VPWR VPWR _21452_/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24393__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20402_ _20400_/Y _20401_/X _20061_/X _20401_/X VGND VGND VPWR VPWR _20402_/X sky130_fd_sc_hd__a2bb2o_4
X_24170_ _24159_/CLK _18559_/Y HRESETn VGND VGND VPWR VPWR _18470_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24322__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21382_ _21962_/A _21380_/X _13771_/A _21381_/X VGND VGND VPWR VPWR _21382_/X sky130_fd_sc_hd__a211o_4
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23121_ _22730_/A VGND VGND VPWR VPWR _23291_/B sky130_fd_sc_hd__buf_2
XFILLER_135_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20333_ _20333_/A VGND VGND VPWR VPWR _20333_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11768__A _25525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23052_ _22774_/X _23048_/Y _22868_/X _23051_/X VGND VGND VPWR VPWR _23053_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22999__C _22998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20264_ _20264_/A VGND VGND VPWR VPWR _22337_/B sky130_fd_sc_hd__inv_2
XFILLER_115_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22003_ _22003_/A _22396_/B VGND VGND VPWR VPWR _22003_/Y sky130_fd_sc_hd__nor2_4
XFILLER_143_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25528__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20195_ _21389_/B _20192_/X _20109_/X _20192_/X VGND VGND VPWR VPWR _23468_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20959__A1_N _20828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22187__B1 _21556_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19052__B1 _18981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_106_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_106_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23954_ _23951_/CLK _23954_/D HRESETn VGND VGND VPWR VPWR _23954_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11934__C _11934_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25110__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22905_ _24631_/Q _22904_/X VGND VGND VPWR VPWR _22905_/X sky130_fd_sc_hd__or2_4
X_23885_ _23887_/CLK _19019_/X VGND VGND VPWR VPWR _18150_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16620__A1_N _16619_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22836_ _22530_/A VGND VGND VPWR VPWR _23022_/B sky130_fd_sc_hd__buf_2
XFILLER_71_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22767_ _24764_/Q _23278_/B VGND VGND VPWR VPWR _22767_/X sky130_fd_sc_hd__or2_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12520_ _25420_/Q VGND VGND VPWR VPWR _12597_/A sky130_fd_sc_hd__inv_2
XFILLER_201_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21718_ _14391_/Y _14183_/X _14452_/Y _17412_/X VGND VGND VPWR VPWR _21719_/D sky130_fd_sc_hd__o22a_4
X_24506_ _24032_/CLK _16651_/X HRESETn VGND VGND VPWR VPWR _24506_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25486_ _23938_/CLK _25486_/D HRESETn VGND VGND VPWR VPWR _12049_/A sky130_fd_sc_hd__dfrtp_4
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22698_ _20887_/Y _21596_/X _16682_/Y _22452_/X VGND VGND VPWR VPWR _22698_/X sky130_fd_sc_hd__o22a_4
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12418_/A _12448_/X VGND VGND VPWR VPWR _12452_/C sky130_fd_sc_hd__or2_4
XANTENNA__21440__A _21439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21649_ _13768_/X VGND VGND VPWR VPWR _21649_/X sky130_fd_sc_hd__buf_2
X_24437_ _24460_/CLK _16811_/X HRESETn VGND VGND VPWR VPWR _16810_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18646__A2_N _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16534__A _16534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15170_ _14972_/Y _15168_/X _15169_/X _15162_/Y VGND VGND VPWR VPWR _15171_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24063__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12382_ _12415_/A VGND VGND VPWR VPWR _12382_/X sky130_fd_sc_hd__buf_2
X_24368_ _24365_/CLK _24368_/D HRESETn VGND VGND VPWR VPWR _24368_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_44_0_HCLK clkbuf_8_45_0_HCLK/A VGND VGND VPWR VPWR _25081_/CLK sky130_fd_sc_hd__clkbuf_1
X_14121_ _14115_/X VGND VGND VPWR VPWR _23955_/D sky130_fd_sc_hd__buf_2
X_23319_ _22286_/X _23309_/X _23319_/C _23318_/X VGND VGND VPWR VPWR _23319_/X sky130_fd_sc_hd__or4_4
XANTENNA__11678__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24299_ _24947_/CLK _17680_/X HRESETn VGND VGND VPWR VPWR _17509_/A sky130_fd_sc_hd__dfrtp_4
X_14052_ _14052_/A VGND VGND VPWR VPWR _14053_/A sky130_fd_sc_hd__buf_2
XANTENNA__22414__A1 _21077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23367__A _21014_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13003_ _12315_/Y _13001_/A VGND VGND VPWR VPWR _13003_/X sky130_fd_sc_hd__or2_4
XANTENNA__12902__A1 _12766_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22702__C _21741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18860_ _24568_/Q _18613_/X _24574_/Q _18698_/A VGND VGND VPWR VPWR _18861_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19291__B1 _19200_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17811_ _17755_/Y _17756_/Y _17555_/X _17811_/D VGND VGND VPWR VPWR _17833_/B sky130_fd_sc_hd__or4_4
X_18791_ _18791_/A _18791_/B VGND VGND VPWR VPWR _18793_/B sky130_fd_sc_hd__or2_4
XFILLER_153_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17742_ _24288_/Q VGND VGND VPWR VPWR _17768_/C sky130_fd_sc_hd__inv_2
XANTENNA__19043__B1 _18951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14954_ _15214_/B _14936_/A _14898_/X _14899_/Y VGND VGND VPWR VPWR _14958_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17054__C1 _17053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13905_ _13904_/X VGND VGND VPWR VPWR _14239_/A sky130_fd_sc_hd__inv_2
XFILLER_75_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17673_ _17577_/C _17676_/B _17593_/X VGND VGND VPWR VPWR _17673_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_47_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14885_ _14885_/A VGND VGND VPWR VPWR _14885_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15604__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19412_ _19412_/A VGND VGND VPWR VPWR _19426_/A sky130_fd_sc_hd__inv_2
XFILLER_208_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16624_ _13729_/Y _16170_/B _16632_/B VGND VGND VPWR VPWR _16624_/X sky130_fd_sc_hd__a21o_4
X_13836_ _21381_/A _13832_/X _13521_/X _13832_/X VGND VGND VPWR VPWR _25256_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22403__A1_N _21284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15080__B2 _16404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19343_ _19343_/A VGND VGND VPWR VPWR _19343_/X sky130_fd_sc_hd__buf_2
X_16555_ _16548_/A VGND VGND VPWR VPWR _16555_/X sky130_fd_sc_hd__buf_2
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24833__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13767_ _19570_/A _14208_/A VGND VGND VPWR VPWR _13768_/A sky130_fd_sc_hd__or2_4
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15506_ _15489_/A VGND VGND VPWR VPWR _15506_/X sky130_fd_sc_hd__buf_2
XANTENNA__13133__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12718_ _12584_/X _12722_/A VGND VGND VPWR VPWR _12718_/Y sky130_fd_sc_hd__nand2_4
X_19274_ _20052_/A _19094_/B _20387_/C VGND VGND VPWR VPWR _19274_/X sky130_fd_sc_hd__or3_4
X_16486_ _16485_/Y _16482_/X _16395_/X _16482_/X VGND VGND VPWR VPWR _24567_/D sky130_fd_sc_hd__a2bb2o_4
X_13698_ _13678_/B _13694_/X _13697_/Y _13690_/X _11826_/A VGND VGND VPWR VPWR _13698_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_231_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12180__A2_N _12178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22446__A _21439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18225_ _18193_/A _23819_/Q VGND VGND VPWR VPWR _18225_/X sky130_fd_sc_hd__or2_4
X_15437_ _14269_/X _24073_/Q _15436_/Y _13927_/B _15433_/X VGND VGND VPWR VPWR _15437_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12649_ _12607_/X _12626_/D _12638_/C VGND VGND VPWR VPWR _12649_/X sky130_fd_sc_hd__o21a_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18156_ _18124_/A _18156_/B _18155_/X VGND VGND VPWR VPWR _18156_/X sky130_fd_sc_hd__or3_4
XANTENNA__18857__B1 _16507_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15368_ _15355_/X VGND VGND VPWR VPWR _15369_/B sky130_fd_sc_hd__inv_2
X_17107_ _17105_/A _17103_/X _17106_/Y VGND VGND VPWR VPWR _17107_/X sky130_fd_sc_hd__and3_4
X_14319_ _14318_/X VGND VGND VPWR VPWR _14349_/A sky130_fd_sc_hd__buf_2
XFILLER_156_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18087_ _18193_/A _23895_/Q VGND VGND VPWR VPWR _18087_/X sky130_fd_sc_hd__or2_4
X_15299_ _15294_/X _15299_/B _15298_/X VGND VGND VPWR VPWR _15300_/C sky130_fd_sc_hd__or3_4
X_17038_ _17125_/A _16982_/Y _17038_/C _17038_/D VGND VGND VPWR VPWR _17038_/X sky130_fd_sc_hd__or4_4
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18989_ _18988_/Y _18986_/X _18942_/X _18986_/X VGND VGND VPWR VPWR _18989_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19034__B1 _18985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20951_ _20828_/X _20950_/Y _24507_/Q _20874_/X VGND VGND VPWR VPWR _20951_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23670_ _23665_/CLK _23670_/D VGND VGND VPWR VPWR _13343_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12409__B1 _12390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20882_ _20870_/X _20881_/Y _24491_/Q _20875_/X VGND VGND VPWR VPWR _20882_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11880__A1 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15071__B2 _16363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22621_ _22515_/X _22619_/X _21956_/X _22620_/Y VGND VGND VPWR VPWR _22621_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15242__B _15242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24574__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14438__A1_N _14158_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25340_ _25341_/CLK _25340_/D HRESETn VGND VGND VPWR VPWR _25340_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22552_ _22132_/B VGND VGND VPWR VPWR _22552_/X sky130_fd_sc_hd__buf_2
XFILLER_179_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24503__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21503_ _21642_/A VGND VGND VPWR VPWR _21503_/X sky130_fd_sc_hd__buf_2
X_25271_ _25325_/CLK _25271_/D HRESETn VGND VGND VPWR VPWR _25271_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22483_ _21424_/X _22482_/X _21427_/X _24864_/Q _21428_/X VGND VGND VPWR VPWR _22484_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_22_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24222_ _23398_/CLK _24222_/D HRESETn VGND VGND VPWR VPWR _21504_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_166_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21434_ _21533_/A VGND VGND VPWR VPWR _23002_/A sky130_fd_sc_hd__buf_2
XFILLER_108_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18848__B1 _24568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_3_0_HCLK clkbuf_8_3_0_HCLK/A VGND VGND VPWR VPWR _23499_/CLK sky130_fd_sc_hd__clkbuf_1
X_24153_ _24148_/CLK _24153_/D HRESETn VGND VGND VPWR VPWR _24153_/Q sky130_fd_sc_hd__dfrtp_4
X_21365_ _21365_/A VGND VGND VPWR VPWR _21365_/X sky130_fd_sc_hd__buf_2
XFILLER_162_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23104_ _21423_/A VGND VGND VPWR VPWR _23280_/A sky130_fd_sc_hd__buf_2
X_20316_ _20315_/Y VGND VGND VPWR VPWR _20316_/X sky130_fd_sc_hd__buf_2
XFILLER_135_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24084_ _25113_/CLK _24084_/D HRESETn VGND VGND VPWR VPWR _20605_/A sky130_fd_sc_hd__dfrtp_4
X_21296_ _21296_/A _15649_/Y _15660_/A _21048_/Y VGND VGND VPWR VPWR _21588_/A sky130_fd_sc_hd__or4_4
X_23035_ _21537_/X VGND VGND VPWR VPWR _23035_/X sky130_fd_sc_hd__buf_2
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25362__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20247_ _20247_/A VGND VGND VPWR VPWR _22075_/B sky130_fd_sc_hd__inv_2
XFILLER_1_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16087__B1 _15991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20178_ _14683_/A _13737_/X _19072_/C _20157_/D VGND VGND VPWR VPWR _20178_/X sky130_fd_sc_hd__or4_4
XFILLER_131_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15834__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24986_ _24976_/CLK _15394_/X HRESETn VGND VGND VPWR VPWR _15295_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_217_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21435__A _21435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11951_ _11951_/A VGND VGND VPWR VPWR _11951_/X sky130_fd_sc_hd__buf_2
X_23937_ _25211_/CLK _23937_/D HRESETn VGND VGND VPWR VPWR _20544_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21383__A1 _13525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11882_ _25515_/Q _11934_/C _11874_/X _11881_/Y VGND VGND VPWR VPWR _11883_/A sky130_fd_sc_hd__a211o_4
X_14670_ _21622_/A VGND VGND VPWR VPWR _22367_/A sky130_fd_sc_hd__buf_2
XFILLER_244_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23868_ _25171_/CLK _19068_/X VGND VGND VPWR VPWR _23868_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_205_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13621_ _13579_/X VGND VGND VPWR VPWR _13621_/Y sky130_fd_sc_hd__inv_2
X_22819_ _23251_/A _22819_/B _22818_/X VGND VGND VPWR VPWR _22819_/X sky130_fd_sc_hd__and3_4
XANTENNA__17339__B1 _17284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23799_ _23808_/CLK _19262_/X VGND VGND VPWR VPWR _19261_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__22332__B1 _14207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16340_ _16339_/Y _16337_/X _16145_/X _16337_/X VGND VGND VPWR VPWR _24620_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_213_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24244__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13552_ _13552_/A VGND VGND VPWR VPWR _13552_/Y sky130_fd_sc_hd__inv_2
X_25538_ _25538_/CLK _25538_/D HRESETn VGND VGND VPWR VPWR _11717_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_158_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21170__A _16852_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12503_ _12503_/A VGND VGND VPWR VPWR _12503_/Y sky130_fd_sc_hd__inv_2
X_13483_ _13483_/A _12086_/X _12058_/C _13483_/D VGND VGND VPWR VPWR _13484_/A sky130_fd_sc_hd__or4_4
X_16271_ _15651_/X _15986_/Y _16267_/X _24645_/Q _16270_/X VGND VGND VPWR VPWR _24645_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_157_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25469_ _25471_/CLK _25469_/D HRESETn VGND VGND VPWR VPWR _25469_/Q sky130_fd_sc_hd__dfrtp_4
X_18010_ _18090_/A VGND VGND VPWR VPWR _18056_/A sky130_fd_sc_hd__buf_2
X_12434_ _12434_/A _12428_/X _12433_/Y VGND VGND VPWR VPWR _12434_/X sky130_fd_sc_hd__and3_4
X_15222_ _25025_/Q _15221_/Y VGND VGND VPWR VPWR _15222_/X sky130_fd_sc_hd__or2_4
XFILLER_145_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12365_ _25341_/Q VGND VGND VPWR VPWR _12979_/D sky130_fd_sc_hd__inv_2
X_15153_ _15153_/A VGND VGND VPWR VPWR _15294_/D sky130_fd_sc_hd__inv_2
XFILLER_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14104_ _14089_/C _14103_/X _14090_/A VGND VGND VPWR VPWR _14105_/B sky130_fd_sc_hd__or3_4
XFILLER_5_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15084_ _15084_/A VGND VGND VPWR VPWR _15084_/Y sky130_fd_sc_hd__inv_2
X_19961_ _19455_/A _18288_/X _18276_/X _19960_/X VGND VGND VPWR VPWR _19962_/A sky130_fd_sc_hd__or4_4
XFILLER_180_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12296_ _12296_/A VGND VGND VPWR VPWR _12296_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14035_ _14034_/X VGND VGND VPWR VPWR _14039_/C sky130_fd_sc_hd__inv_2
X_18912_ _18911_/X VGND VGND VPWR VPWR _18925_/A sky130_fd_sc_hd__inv_2
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19892_ _21676_/B _19891_/X _19617_/X _19891_/X VGND VGND VPWR VPWR _19892_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16078__B1 _24714_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21071__B1 _21047_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25032__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18843_ _16456_/A _24156_/Q _16456_/Y _18700_/C VGND VGND VPWR VPWR _18845_/C sky130_fd_sc_hd__o22a_4
XFILLER_68_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15825__B1 _15616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19016__B1 _18965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18774_ _18774_/A _18745_/D VGND VGND VPWR VPWR _18774_/X sky130_fd_sc_hd__or2_4
X_15986_ _16270_/B VGND VGND VPWR VPWR _15986_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21990__D _21990_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17725_ _17725_/A VGND VGND VPWR VPWR _17725_/X sky130_fd_sc_hd__buf_2
XFILLER_209_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14937_ _25013_/Q VGND VGND VPWR VPWR _15261_/A sky130_fd_sc_hd__inv_2
XFILLER_236_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21374__A1 _21345_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12967__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15343__A _15282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17656_ _17614_/A _17581_/X VGND VGND VPWR VPWR _17656_/X sky130_fd_sc_hd__or2_4
XANTENNA__21064__B _21064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14868_ _14864_/Y _14867_/Y _14859_/X VGND VGND VPWR VPWR _14868_/X sky130_fd_sc_hd__o21a_4
XFILLER_208_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16250__B1 _16055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16607_ _16605_/Y _16606_/X _16522_/X _16606_/X VGND VGND VPWR VPWR _24521_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_224_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13819_ _22540_/A _13817_/X _13818_/X _13817_/X VGND VGND VPWR VPWR _25265_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17587_ _17587_/A _17586_/X VGND VGND VPWR VPWR _17587_/X sky130_fd_sc_hd__or2_4
X_14799_ _14798_/X VGND VGND VPWR VPWR _14799_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21126__B2 _15661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19326_ _18048_/B VGND VGND VPWR VPWR _19326_/Y sky130_fd_sc_hd__inv_2
X_16538_ _24546_/Q VGND VGND VPWR VPWR _16538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12811__B1 _25388_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22874__B2 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16002__B1 _16001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19257_ _22214_/B _19254_/X _16864_/X _19254_/X VGND VGND VPWR VPWR _23801_/D sky130_fd_sc_hd__a2bb2o_4
X_16469_ _16469_/A VGND VGND VPWR VPWR _16469_/Y sky130_fd_sc_hd__inv_2
X_18208_ _14636_/A _18208_/B _18207_/X VGND VGND VPWR VPWR _18208_/X sky130_fd_sc_hd__and3_4
X_19188_ _18018_/B VGND VGND VPWR VPWR _19188_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23967__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18139_ _17979_/X _18139_/B VGND VGND VPWR VPWR _18139_/X sky130_fd_sc_hd__or2_4
XFILLER_144_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16902__A _24276_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21150_ _12081_/A _24191_/Q _25170_/Q _13457_/D VGND VGND VPWR VPWR _21150_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_90_0_HCLK clkbuf_8_91_0_HCLK/A VGND VGND VPWR VPWR _25369_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_172_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20101_ _23502_/Q VGND VGND VPWR VPWR _20101_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21081_ _21080_/X VGND VGND VPWR VPWR _22523_/B sky130_fd_sc_hd__buf_2
XANTENNA__14422__A _14422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20032_ _20157_/C _13744_/X _13753_/X _13754_/X VGND VGND VPWR VPWR _20032_/X sky130_fd_sc_hd__or4_4
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15816__B1 _24833_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19007__B1 _19006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24840_ _24809_/CLK _24840_/D HRESETn VGND VGND VPWR VPWR _24840_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18663__A1_N _16613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21255__A _22199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15831__A3 _15830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21983_ _21983_/A _20318_/X VGND VGND VPWR VPWR _21983_/X sky130_fd_sc_hd__and2_4
X_24771_ _25380_/CLK _24771_/D HRESETn VGND VGND VPWR VPWR _23036_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24755__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16349__A _14380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22562__B1 _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11781__A _14392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20934_ _20919_/X _20933_/Y _24503_/Q _20923_/X VGND VGND VPWR VPWR _20934_/X sky130_fd_sc_hd__a2bb2o_4
X_23722_ _23406_/CLK _23722_/D VGND VGND VPWR VPWR _19477_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_226_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16241__B1 _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15044__B2 _24477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20865_ _20864_/X VGND VGND VPWR VPWR _24043_/D sky130_fd_sc_hd__inv_2
X_23653_ _23665_/CLK _19686_/X VGND VGND VPWR VPWR _13372_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_53_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22604_ _15605_/Y _22756_/B VGND VGND VPWR VPWR _22604_/X sky130_fd_sc_hd__and2_4
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23584_ _23559_/CLK _23584_/D VGND VGND VPWR VPWR _19883_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_223_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12802__B1 _12801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20796_ _20796_/A VGND VGND VPWR VPWR _20796_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22535_ _23178_/A VGND VGND VPWR VPWR _22535_/X sky130_fd_sc_hd__buf_2
X_25323_ _23887_/CLK _25323_/D HRESETn VGND VGND VPWR VPWR _13466_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22466_ _22466_/A VGND VGND VPWR VPWR _23129_/A sky130_fd_sc_hd__buf_2
X_25254_ _24958_/CLK _13843_/X HRESETn VGND VGND VPWR VPWR _25254_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15898__A3 _15830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22814__A _22814_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16941__A2_N _16940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21417_ _21382_/X _21383_/X _22515_/A _21416_/X VGND VGND VPWR VPWR _21418_/A sky130_fd_sc_hd__a211o_4
X_24205_ _23391_/CLK _18345_/X HRESETn VGND VGND VPWR VPWR _13187_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25543__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25185_ _25249_/CLK _14265_/X HRESETn VGND VGND VPWR VPWR _14264_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22093__A2 _22420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19395__A _18985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22397_ _23706_/Q _22397_/B VGND VGND VPWR VPWR _22397_/X sky130_fd_sc_hd__or2_4
X_12150_ _18372_/D VGND VGND VPWR VPWR _12150_/Y sky130_fd_sc_hd__inv_2
X_24136_ _24139_/CLK _18796_/Y HRESETn VGND VGND VPWR VPWR _24136_/Q sky130_fd_sc_hd__dfrtp_4
X_21348_ _21348_/A VGND VGND VPWR VPWR _21349_/A sky130_fd_sc_hd__buf_2
XFILLER_162_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_118_0_HCLK clkbuf_7_59_0_HCLK/X VGND VGND VPWR VPWR _24834_/CLK sky130_fd_sc_hd__clkbuf_1
X_12081_ _12081_/A VGND VGND VPWR VPWR _12082_/A sky130_fd_sc_hd__buf_2
X_24067_ _25346_/CLK _23339_/X HRESETn VGND VGND VPWR VPWR _24067_/Q sky130_fd_sc_hd__dfrtp_4
X_21279_ _21379_/B _21277_/X _25271_/Q _21278_/X VGND VGND VPWR VPWR _21279_/X sky130_fd_sc_hd__o22a_4
X_23018_ _24057_/Q _21303_/A _13108_/C _21598_/X VGND VGND VPWR VPWR _23018_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15807__B1 _11715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15840_ _15651_/X _15761_/X _15838_/X _12592_/A _15839_/X VGND VGND VPWR VPWR _15840_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16480__B1 _16391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21165__A _16619_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15771_ _15773_/A _15771_/B VGND VGND VPWR VPWR _15771_/X sky130_fd_sc_hd__or2_4
XANTENNA__24496__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12983_ _12330_/Y _13069_/A _13068_/C _12983_/D VGND VGND VPWR VPWR _12983_/X sky130_fd_sc_hd__or4_4
X_24969_ _24959_/CLK _15442_/X HRESETn VGND VGND VPWR VPWR _13878_/B sky130_fd_sc_hd__dfrtp_4
X_17510_ _25528_/Q _17509_/A _11755_/Y _17670_/A VGND VGND VPWR VPWR _17515_/B sky130_fd_sc_hd__o22a_4
XANTENNA__11691__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14722_ _22043_/A VGND VGND VPWR VPWR _14722_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11934_ _11934_/A _11934_/B _11934_/C VGND VGND VPWR VPWR _17442_/B sky130_fd_sc_hd__or3_4
X_18490_ _18457_/Y _18483_/X _18484_/Y _18489_/X VGND VGND VPWR VPWR _18491_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24425__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17441_ _17435_/Y _17438_/Y _17440_/X _17438_/Y VGND VGND VPWR VPWR _17441_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14653_ _14652_/X VGND VGND VPWR VPWR _14654_/A sky130_fd_sc_hd__buf_2
XFILLER_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11865_ _11864_/X VGND VGND VPWR VPWR _11865_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _19116_/A VGND VGND VPWR VPWR _13606_/A sky130_fd_sc_hd__inv_2
XPHY_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17372_ _17372_/A VGND VGND VPWR VPWR _24345_/D sky130_fd_sc_hd__inv_2
XPHY_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11796_ _11796_/A _11796_/B VGND VGND VPWR VPWR _11860_/A sky130_fd_sc_hd__and2_4
X_14584_ _14557_/B _14575_/X _14583_/Y _14579_/X _13563_/A VGND VGND VPWR VPWR _14584_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_41_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19111_ _23852_/Q VGND VGND VPWR VPWR _19111_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15520__A2_N _15519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16323_ _16322_/Y _16319_/X _16226_/X _16319_/X VGND VGND VPWR VPWR _24627_/D sky130_fd_sc_hd__a2bb2o_4
X_13535_ _13535_/A VGND VGND VPWR VPWR _14554_/A sky130_fd_sc_hd__inv_2
XFILLER_158_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19042_ _23876_/Q VGND VGND VPWR VPWR _19042_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16254_ _22097_/A VGND VGND VPWR VPWR _16254_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13466_ _13466_/A VGND VGND VPWR VPWR _13466_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15205_ _15229_/A _15039_/X _15205_/C VGND VGND VPWR VPWR _15214_/D sky130_fd_sc_hd__or3_4
XANTENNA__25284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12417_ _12263_/A VGND VGND VPWR VPWR _12434_/A sky130_fd_sc_hd__buf_2
XFILLER_127_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16185_ _16184_/X VGND VGND VPWR VPWR _16185_/X sky130_fd_sc_hd__buf_2
X_13397_ _13397_/A _13395_/X _13397_/C VGND VGND VPWR VPWR _13397_/X sky130_fd_sc_hd__and3_4
XANTENNA__16299__B1 _15939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_14_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__25213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15136_ _15129_/X _15136_/B _15136_/C _15136_/D VGND VGND VPWR VPWR _15136_/X sky130_fd_sc_hd__or4_4
X_12348_ _12341_/X _12343_/X _12348_/C _12347_/X VGND VGND VPWR VPWR _12369_/B sky130_fd_sc_hd__or4_4
Xclkbuf_7_77_0_HCLK clkbuf_7_77_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_77_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22162__C _22161_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21350__A2_N _22327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12279_ _12279_/A _12279_/B VGND VGND VPWR VPWR _12379_/A sky130_fd_sc_hd__or2_4
X_15067_ _15182_/A _15067_/B VGND VGND VPWR VPWR _15160_/A sky130_fd_sc_hd__or2_4
X_19944_ _19943_/Y _19941_/X _19603_/X _19941_/X VGND VGND VPWR VPWR _19944_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14018_ _13986_/X _13987_/X _13979_/C _25234_/Q VGND VGND VPWR VPWR _14018_/X sky130_fd_sc_hd__a211o_4
XFILLER_110_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19875_ _21200_/B _19869_/X _19874_/X _19856_/Y VGND VGND VPWR VPWR _23587_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_229_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12795__A1_N _22667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18826_ _16490_/Y _24144_/Q _16490_/Y _24144_/Q VGND VGND VPWR VPWR _18826_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16471__B1 _16382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21075__A _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18757_ _18693_/C _18755_/X _18756_/Y VGND VGND VPWR VPWR _18757_/X sky130_fd_sc_hd__o21a_4
X_15969_ _12192_/Y _15964_/X _15754_/X _15968_/X VGND VGND VPWR VPWR _24756_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17703__D _21176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17708_ _17707_/X VGND VGND VPWR VPWR _17709_/A sky130_fd_sc_hd__buf_2
XFILLER_36_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24166__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18688_ _24138_/Q VGND VGND VPWR VPWR _18694_/B sky130_fd_sc_hd__inv_2
XFILLER_224_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23290__A _23288_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17639_ _17523_/Y _17646_/A _17648_/A _17648_/B VGND VGND VPWR VPWR _17645_/B sky130_fd_sc_hd__or4_4
XFILLER_224_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20650_ _14227_/Y _20638_/X _20629_/X _20649_/X VGND VGND VPWR VPWR _20651_/A sky130_fd_sc_hd__a211o_4
XFILLER_223_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22847__B2 _22846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19309_ _19308_/Y _19306_/X _19194_/X _19306_/X VGND VGND VPWR VPWR _19309_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20581_ _18880_/B _20580_/Y _20572_/X VGND VGND VPWR VPWR _20581_/X sky130_fd_sc_hd__and3_4
XFILLER_177_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22320_ _22313_/Y _22315_/Y _22316_/X _22320_/D VGND VGND VPWR VPWR _22320_/X sky130_fd_sc_hd__or4_4
XFILLER_149_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22251_ _22251_/A _22251_/B VGND VGND VPWR VPWR _22253_/B sky130_fd_sc_hd__or2_4
XFILLER_180_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12748__A1_N _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21202_ _21204_/A _21202_/B _21202_/C VGND VGND VPWR VPWR _21202_/X sky130_fd_sc_hd__and3_4
XFILLER_191_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22182_ _15460_/Y _21365_/X _14215_/Y _21351_/X VGND VGND VPWR VPWR _22183_/A sky130_fd_sc_hd__o22a_4
XFILLER_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17447__B _21177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11771__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21318__A2_N _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21133_ _21133_/A _21133_/B _13807_/A _17703_/B VGND VGND VPWR VPWR _21343_/B sky130_fd_sc_hd__or4_4
XFILLER_120_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21064_ _21064_/A _21064_/B VGND VGND VPWR VPWR _21064_/X sky130_fd_sc_hd__or2_4
XFILLER_120_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24936__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22783__B1 _12740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20015_ _23537_/Q VGND VGND VPWR VPWR _22262_/B sky130_fd_sc_hd__inv_2
XFILLER_48_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23184__B _22658_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_28_0_HCLK_A clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16462__B1 _16459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23327__A2 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24823_ _24855_/CLK _24823_/D HRESETn VGND VGND VPWR VPWR _24823_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24754_ _25369_/CLK _24754_/D HRESETn VGND VGND VPWR VPWR _22276_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_64_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21966_ _21963_/X _21964_/X _21965_/X VGND VGND VPWR VPWR _21966_/Y sky130_fd_sc_hd__o21ai_4
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ _23706_/CLK _23705_/D VGND VGND VPWR VPWR _19528_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21713__A _21711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _24055_/Q _20911_/A _20916_/X VGND VGND VPWR VPWR _20917_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21897_ _22083_/A _21897_/B VGND VGND VPWR VPWR _21899_/B sky130_fd_sc_hd__or2_4
X_24685_ _24704_/CLK _24685_/D HRESETn VGND VGND VPWR VPWR _16154_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_214_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/A VGND VGND VPWR VPWR _11650_/Y sky130_fd_sc_hd__inv_2
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _20847_/Y _20842_/Y _13644_/X VGND VGND VPWR VPWR _20848_/X sky130_fd_sc_hd__o21a_4
X_23636_ _23644_/CLK _23636_/D VGND VGND VPWR VPWR _13411_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ _20753_/X _20778_/Y _15583_/A _20757_/X VGND VGND VPWR VPWR _24023_/D sky130_fd_sc_hd__a2bb2o_4
X_23567_ _25070_/CLK _19928_/X VGND VGND VPWR VPWR _23567_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13231__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _13353_/A _13309_/X _13319_/X VGND VGND VPWR VPWR _13320_/X sky130_fd_sc_hd__and3_4
X_25306_ _25308_/CLK _25306_/D HRESETn VGND VGND VPWR VPWR _12013_/C sky130_fd_sc_hd__dfrtp_4
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22518_ _22515_/X _22516_/X _21956_/A _22517_/Y VGND VGND VPWR VPWR _22518_/X sky130_fd_sc_hd__o22a_4
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23498_ _24199_/CLK _23498_/D VGND VGND VPWR VPWR _23498_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17190__B2 _17251_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13251_ _13390_/A _13251_/B _13251_/C VGND VGND VPWR VPWR _13255_/B sky130_fd_sc_hd__and3_4
X_22449_ _22445_/X _22447_/X _22876_/C VGND VGND VPWR VPWR _22449_/X sky130_fd_sc_hd__or3_4
X_25237_ _23976_/CLK _14066_/X HRESETn VGND VGND VPWR VPWR _25237_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16542__A _16541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12202_ _22898_/A VGND VGND VPWR VPWR _12202_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13182_ _11950_/A _11961_/C VGND VGND VPWR VPWR _13182_/Y sky130_fd_sc_hd__nor2_4
X_25168_ _25479_/CLK _25168_/D HRESETn VGND VGND VPWR VPWR _25168_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11762__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12133_ _12133_/A _12133_/B _12128_/X _12132_/X VGND VGND VPWR VPWR _12133_/X sky130_fd_sc_hd__or4_4
X_24119_ _25224_/CLK _18894_/X HRESETn VGND VGND VPWR VPWR _20982_/B sky130_fd_sc_hd__dfstp_4
XANTENNA__19219__B1 _19194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17990_ _18095_/A VGND VGND VPWR VPWR _17990_/X sky130_fd_sc_hd__buf_2
X_25099_ _25100_/CLK _25099_/D HRESETn VGND VGND VPWR VPWR _25099_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12064_ _25484_/Q VGND VGND VPWR VPWR _12064_/Y sky130_fd_sc_hd__inv_2
X_16941_ _24703_/Q _16940_/Y _16113_/Y _24278_/Q VGND VGND VPWR VPWR _16942_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24677__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19660_ _19659_/Y _19657_/X _19534_/X _19657_/X VGND VGND VPWR VPWR _23663_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22710__C _21864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17373__A _17203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16872_ _19820_/A VGND VGND VPWR VPWR _16872_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24606__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18611_ _24525_/Q _18789_/C _16554_/Y _24152_/Q VGND VGND VPWR VPWR _18618_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15823_ _15820_/A VGND VGND VPWR VPWR _15823_/X sky130_fd_sc_hd__buf_2
XFILLER_77_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19591_ _19589_/Y _19590_/X _19540_/X _19590_/X VGND VGND VPWR VPWR _23685_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18542_ _18467_/B _18538_/X VGND VGND VPWR VPWR _18542_/Y sky130_fd_sc_hd__nand2_4
X_15754_ HWDATA[8] VGND VGND VPWR VPWR _15754_/X sky130_fd_sc_hd__buf_2
X_12966_ _21027_/A _12650_/A VGND VGND VPWR VPWR _12967_/C sky130_fd_sc_hd__or2_4
XFILLER_205_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14705_ _14705_/A VGND VGND VPWR VPWR _14706_/A sky130_fd_sc_hd__inv_2
XANTENNA__21623__A _22381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11917_ _19981_/A VGND VGND VPWR VPWR _19617_/A sky130_fd_sc_hd__buf_2
X_18473_ _18473_/A VGND VGND VPWR VPWR _18473_/Y sky130_fd_sc_hd__inv_2
X_15685_ _15684_/X VGND VGND VPWR VPWR _24889_/D sky130_fd_sc_hd__inv_2
X_12897_ _12889_/X _12897_/B _12897_/C VGND VGND VPWR VPWR _25389_/D sky130_fd_sc_hd__and3_4
XFILLER_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17424_ _24330_/Q VGND VGND VPWR VPWR _17424_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15621__A _24898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14636_ _14636_/A VGND VGND VPWR VPWR _18123_/A sky130_fd_sc_hd__buf_2
XFILLER_220_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11848_ _11848_/A _11848_/B VGND VGND VPWR VPWR _11849_/B sky130_fd_sc_hd__and2_4
XFILLER_20_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17352_/B _17352_/C VGND VGND VPWR VPWR _17358_/B sky130_fd_sc_hd__or2_4
XFILLER_158_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14567_ _25097_/Q _14566_/X _14564_/Y VGND VGND VPWR VPWR _14567_/X sky130_fd_sc_hd__o21a_4
XFILLER_20_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11779_ HWDATA[3] VGND VGND VPWR VPWR _11780_/A sky130_fd_sc_hd__buf_2
XFILLER_147_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16306_ _16284_/X VGND VGND VPWR VPWR _16306_/X sky130_fd_sc_hd__buf_2
XANTENNA__13141__A _13168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13518_ _25304_/Q VGND VGND VPWR VPWR SSn_S2 sky130_fd_sc_hd__inv_2
XFILLER_186_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17286_ _17284_/X _17280_/Y _17285_/X VGND VGND VPWR VPWR _17286_/X sky130_fd_sc_hd__or3_4
X_14498_ _25111_/Q _14496_/X _14491_/X _14497_/Y VGND VGND VPWR VPWR _14498_/X sky130_fd_sc_hd__a211o_4
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19025_ _13613_/A VGND VGND VPWR VPWR _19163_/B sky130_fd_sc_hd__buf_2
X_16237_ _16235_/Y _16230_/X _16236_/X _16230_/X VGND VGND VPWR VPWR _24659_/D sky130_fd_sc_hd__a2bb2o_4
X_13449_ _13385_/A _13441_/X _13448_/X VGND VGND VPWR VPWR _13449_/X sky130_fd_sc_hd__and3_4
XFILLER_173_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23254__A1 _24745_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16452__A _16724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21265__B1 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16168_ RsRx_S0 _16167_/Y _14763_/Y VGND VGND VPWR VPWR _16168_/X sky130_fd_sc_hd__a21o_4
XFILLER_114_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15119_ _15132_/A _15117_/Y _15298_/A _15121_/A VGND VGND VPWR VPWR _15127_/A sky130_fd_sc_hd__a2bb2o_4
X_16099_ _16111_/A VGND VGND VPWR VPWR _16099_/X sky130_fd_sc_hd__buf_2
XFILLER_141_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19927_ _23567_/Q VGND VGND VPWR VPWR _19927_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_101_0_HCLK clkbuf_7_50_0_HCLK/X VGND VGND VPWR VPWR _24762_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_164_0_HCLK clkbuf_7_82_0_HCLK/X VGND VGND VPWR VPWR _23875_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_68_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24347__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_7_0_HCLK clkbuf_7_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19858_ _22339_/B _19857_/X _19600_/X _19857_/X VGND VGND VPWR VPWR _19858_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_229_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18809_ _18793_/A _18809_/B _18808_/Y VGND VGND VPWR VPWR _24132_/D sky130_fd_sc_hd__and3_4
XFILLER_244_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19789_ _19784_/A VGND VGND VPWR VPWR _19789_/X sky130_fd_sc_hd__buf_2
XANTENNA__15798__A2 _15789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20791__A2 _20708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21820_ _21954_/A _21812_/X _21819_/X VGND VGND VPWR VPWR _21820_/X sky130_fd_sc_hd__or3_4
XANTENNA__12220__A _22150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21751_ _21720_/Y _21735_/X _21751_/C _21750_/X VGND VGND VPWR VPWR _21751_/X sky130_fd_sc_hd__or4_4
XFILLER_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20702_ _21746_/A _20687_/X _20696_/X _20701_/X VGND VGND VPWR VPWR _20702_/X sky130_fd_sc_hd__o22a_4
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21682_ _21484_/X _21680_/X _21682_/C VGND VGND VPWR VPWR _21682_/X sky130_fd_sc_hd__and3_4
X_24470_ _24460_/CLK _24470_/D HRESETn VGND VGND VPWR VPWR _15037_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_196_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23982__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20633_ _20632_/X VGND VGND VPWR VPWR _23978_/D sky130_fd_sc_hd__inv_2
X_23421_ _23425_/CLK _23421_/D VGND VGND VPWR VPWR _23421_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23352_ VGND VGND VPWR VPWR _23352_/HI IRQ[28] sky130_fd_sc_hd__conb_1
X_20564_ _14428_/Y _20543_/X _20557_/X _20563_/X VGND VGND VPWR VPWR _20565_/A sky130_fd_sc_hd__a211o_4
XFILLER_164_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22303_ _22286_/X _22293_/Y _22298_/X _22140_/A _22302_/X VGND VGND VPWR VPWR _22304_/D
+ sky130_fd_sc_hd__o32a_4
X_23283_ _23282_/X VGND VGND VPWR VPWR _23283_/Y sky130_fd_sc_hd__inv_2
X_20495_ _14266_/Y _20502_/B _20495_/C VGND VGND VPWR VPWR _20495_/X sky130_fd_sc_hd__and3_4
XFILLER_118_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12890__A _22667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22234_ _21208_/A VGND VGND VPWR VPWR _22251_/A sky130_fd_sc_hd__buf_2
X_25022_ _25028_/CLK _25022_/D HRESETn VGND VGND VPWR VPWR _25022_/Q sky130_fd_sc_hd__dfrtp_4
X_22165_ _16605_/A _21325_/X _15663_/A _22164_/X VGND VGND VPWR VPWR _22166_/C sky130_fd_sc_hd__a211o_4
XFILLER_246_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_60_0_HCLK clkbuf_7_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21116_ _21077_/X _21078_/X _21097_/X _21110_/X _21115_/X VGND VGND VPWR VPWR _21288_/C
+ sky130_fd_sc_hd__a32o_4
XFILLER_132_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16683__B1 _15741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21708__A _21080_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22096_ _22995_/A VGND VGND VPWR VPWR _22708_/A sky130_fd_sc_hd__buf_2
XANTENNA__24770__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13497__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21047_ _21579_/B VGND VGND VPWR VPWR _21047_/X sky130_fd_sc_hd__buf_2
XANTENNA__19621__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14610__A _14610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24017__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16926__A1_N _21435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12820_ _12828_/A _12808_/Y _12807_/X _24789_/Q VGND VGND VPWR VPWR _12820_/X sky130_fd_sc_hd__a2bb2o_4
X_24806_ _24804_/CLK _15873_/X HRESETn VGND VGND VPWR VPWR _22972_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22998_ _16566_/A _22884_/X _22928_/X _22997_/X VGND VGND VPWR VPWR _22998_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22539__A _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12751_ _12742_/X _12745_/X _12751_/C _12751_/D VGND VGND VPWR VPWR _12751_/X sky130_fd_sc_hd__or4_4
X_24737_ _24737_/CLK _16021_/X HRESETn VGND VGND VPWR VPWR _24737_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ _21462_/A _21949_/B _21948_/X VGND VGND VPWR VPWR _21949_/X sky130_fd_sc_hd__and3_4
XFILLER_215_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11701_/X VGND VGND VPWR VPWR _15981_/A sky130_fd_sc_hd__buf_2
XFILLER_188_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15468_/Y _15463_/X _15469_/X _15463_/X VGND VGND VPWR VPWR _15470_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12553_/Y _12681_/X VGND VGND VPWR VPWR _12682_/X sky130_fd_sc_hd__or2_4
X_24668_ _24662_/CLK _16211_/X HRESETn VGND VGND VPWR VPWR _22996_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_203_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _25137_/Q VGND VGND VPWR VPWR _14421_/Y sky130_fd_sc_hd__inv_2
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ _23859_/CLK _23619_/D VGND VGND VPWR VPWR _23619_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15160__B _15311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19688__B1 _19543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12224__B2 _24760_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24599_ _24551_/CLK _24599_/D HRESETn VGND VGND VPWR VPWR _15091_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17140_ _17142_/A _17140_/B _17140_/C VGND VGND VPWR VPWR _24381_/D sky130_fd_sc_hd__and3_4
XANTENNA__14193__A1_N _20510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14352_ _14344_/X _14351_/X _25484_/Q _14349_/X VGND VGND VPWR VPWR _14352_/X sky130_fd_sc_hd__o22a_4
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22274__A _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _13264_/X _13303_/B VGND VGND VPWR VPWR _13303_/X sky130_fd_sc_hd__or2_4
XFILLER_7_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17071_ _17045_/X _17062_/X _17023_/Y VGND VGND VPWR VPWR _17071_/X sky130_fd_sc_hd__o21a_4
XFILLER_156_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14283_ _14283_/A _14283_/B VGND VGND VPWR VPWR _14288_/A sky130_fd_sc_hd__or2_4
XFILLER_109_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16022_ _24736_/Q VGND VGND VPWR VPWR _16022_/Y sky130_fd_sc_hd__inv_2
X_13234_ _13421_/A VGND VGND VPWR VPWR _13234_/X sky130_fd_sc_hd__buf_2
XFILLER_170_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24858__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16269__A3 _16267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13165_ _13284_/A VGND VGND VPWR VPWR _13385_/A sky130_fd_sc_hd__inv_2
XFILLER_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16674__B1 _16400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12116_ _24105_/Q _12129_/A VGND VGND VPWR VPWR _12116_/X sky130_fd_sc_hd__and2_4
XFILLER_2_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13096_ _13097_/A _13097_/B VGND VGND VPWR VPWR _13098_/A sky130_fd_sc_hd__nand2_4
X_17973_ _17968_/X _17973_/B _17973_/C VGND VGND VPWR VPWR _17973_/X sky130_fd_sc_hd__and3_4
X_12047_ _12047_/A VGND VGND VPWR VPWR _12047_/Y sky130_fd_sc_hd__inv_2
X_16924_ _17752_/C VGND VGND VPWR VPWR _17880_/A sky130_fd_sc_hd__buf_2
X_19712_ _19710_/Y _19707_/X _19711_/X _19707_/X VGND VGND VPWR VPWR _19712_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15616__A _14400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24440__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_237_0_HCLK clkbuf_8_237_0_HCLK/A VGND VGND VPWR VPWR _25056_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16855_ _16854_/X VGND VGND VPWR VPWR _16855_/Y sky130_fd_sc_hd__inv_2
X_19643_ _13407_/B VGND VGND VPWR VPWR _19643_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15806_ _15792_/X VGND VGND VPWR VPWR _15806_/X sky130_fd_sc_hd__buf_2
X_19574_ _13807_/A _13807_/B _13763_/X _19573_/X VGND VGND VPWR VPWR _19575_/A sky130_fd_sc_hd__and4_4
X_16786_ _16786_/A VGND VGND VPWR VPWR _16786_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12040__A _21574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13998_ _13989_/X _13997_/X VGND VGND VPWR VPWR _13999_/C sky130_fd_sc_hd__or2_4
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18525_ _18468_/C _18524_/X VGND VGND VPWR VPWR _18526_/B sky130_fd_sc_hd__or2_4
X_15737_ _15724_/X _15709_/X _15735_/X _24871_/Q _15736_/X VGND VGND VPWR VPWR _15737_/X
+ sky130_fd_sc_hd__a32o_4
X_12949_ _12762_/Y _12952_/B _12854_/X VGND VGND VPWR VPWR _12949_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_80_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18456_ _18580_/A VGND VGND VPWR VPWR _18497_/A sky130_fd_sc_hd__buf_2
XFILLER_34_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15668_ _22530_/A VGND VGND VPWR VPWR _22890_/B sky130_fd_sc_hd__buf_2
XFILLER_233_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17407_ _17384_/A _17398_/A _23990_/Q _21000_/B _17401_/A VGND VGND VPWR VPWR _17407_/X
+ sky130_fd_sc_hd__a32o_4
X_14619_ _14619_/A _14607_/Y VGND VGND VPWR VPWR _14619_/Y sky130_fd_sc_hd__nor2_4
XFILLER_194_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18387_ _18385_/Y _18386_/X _24192_/Q _18386_/X VGND VGND VPWR VPWR _18387_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15599_ _15598_/Y _15596_/X _11735_/X _15596_/X VGND VGND VPWR VPWR _15599_/X sky130_fd_sc_hd__a2bb2o_4
X_17338_ _17338_/A _17338_/B _17337_/X VGND VGND VPWR VPWR _17338_/X sky130_fd_sc_hd__and3_4
XFILLER_174_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17269_ _17232_/Y _17266_/X _17260_/B _17268_/X VGND VGND VPWR VPWR _17270_/A sky130_fd_sc_hd__a211o_4
XFILLER_162_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19008_ _19008_/A VGND VGND VPWR VPWR _19008_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20280_ _21655_/B _20279_/X _19981_/X _20279_/X VGND VGND VPWR VPWR _20280_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24599__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22986__B1 _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17011__A1_N _24744_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24528__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_47_0_HCLK clkbuf_6_46_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22738__B1 _22737_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24181__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23970_ _25243_/CLK _21007_/Y HRESETn VGND VGND VPWR VPWR _21008_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_229_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22921_ _16670_/Y _22921_/B VGND VGND VPWR VPWR _22921_/X sky130_fd_sc_hd__and2_4
XANTENNA__24110__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22852_ _22761_/X _22850_/X _22437_/A _22851_/X VGND VGND VPWR VPWR _22853_/A sky130_fd_sc_hd__o22a_4
XFILLER_25_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22359__A _21936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21803_ _21803_/A _21803_/B _21803_/C VGND VGND VPWR VPWR _21803_/X sky130_fd_sc_hd__and3_4
XANTENNA__25387__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22783_ _17314_/C _22430_/X _12740_/A _22299_/X VGND VGND VPWR VPWR _22784_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15261__A _15261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24522_ _24539_/CLK _16604_/X HRESETn VGND VGND VPWR VPWR _24522_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21734_ _21733_/X VGND VGND VPWR VPWR _21734_/Y sky130_fd_sc_hd__inv_2
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12206__A1 _12204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24453_ _24073_/CLK _16773_/X HRESETn VGND VGND VPWR VPWR _24453_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21665_ _21665_/A _21665_/B VGND VGND VPWR VPWR _21665_/X sky130_fd_sc_hd__or2_4
XFILLER_101_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23404_ _23675_/CLK _20363_/X VGND VGND VPWR VPWR _20361_/A sky130_fd_sc_hd__dfxtp_4
X_20616_ _17385_/B _17401_/A VGND VGND VPWR VPWR _20616_/X sky130_fd_sc_hd__and2_4
X_21596_ _22466_/A VGND VGND VPWR VPWR _21596_/X sky130_fd_sc_hd__buf_2
X_24384_ _24377_/CLK _24384_/D HRESETn VGND VGND VPWR VPWR _24384_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20547_ _18872_/A _20544_/A VGND VGND VPWR VPWR _20547_/Y sky130_fd_sc_hd__nand2_4
X_23335_ _24445_/Q _22282_/A _22801_/X _23334_/X VGND VGND VPWR VPWR _23336_/C sky130_fd_sc_hd__a211o_4
XFILLER_153_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20478_ _20477_/X VGND VGND VPWR VPWR _20478_/Y sky130_fd_sc_hd__inv_2
X_23266_ _22824_/X _23257_/Y _23261_/Y _23265_/X VGND VGND VPWR VPWR _23266_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16850__A1_N _14932_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25005_ _25005_/CLK _25005_/D HRESETn VGND VGND VPWR VPWR _25005_/Q sky130_fd_sc_hd__dfrtp_4
X_22217_ _22221_/A _22217_/B VGND VGND VPWR VPWR _22217_/X sky130_fd_sc_hd__or2_4
XFILLER_180_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23197_ _12279_/A _22984_/X _24285_/Q _22493_/X VGND VGND VPWR VPWR _23197_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18645__B2 _24138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24269__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16656__B1 _16295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22148_ _24721_/Q _22282_/A _22525_/A _22147_/X VGND VGND VPWR VPWR _22148_/X sky130_fd_sc_hd__a211o_4
XFILLER_0_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14970_ _25011_/Q VGND VGND VPWR VPWR _14970_/Y sky130_fd_sc_hd__inv_2
X_22079_ _22378_/A _20120_/Y VGND VGND VPWR VPWR _22079_/X sky130_fd_sc_hd__or2_4
XFILLER_121_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13921_ _24974_/Q VGND VGND VPWR VPWR _13938_/B sky130_fd_sc_hd__inv_2
XFILLER_48_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20996__B _14185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16640_ _16640_/A VGND VGND VPWR VPWR _16660_/A sky130_fd_sc_hd__inv_2
X_13852_ _13840_/C VGND VGND VPWR VPWR _13852_/X sky130_fd_sc_hd__buf_2
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_67_0_HCLK clkbuf_8_67_0_HCLK/A VGND VGND VPWR VPWR _24686_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12803_ _12803_/A _12797_/X _12799_/X _12802_/X VGND VGND VPWR VPWR _12824_/B sky130_fd_sc_hd__or4_4
XFILLER_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16571_ _16571_/A VGND VGND VPWR VPWR _16571_/Y sky130_fd_sc_hd__inv_2
X_13783_ _16721_/A _16721_/B _13772_/C _13783_/D VGND VGND VPWR VPWR _13792_/A sky130_fd_sc_hd__and4_4
XFILLER_204_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16267__A _13797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18310_ _21920_/A VGND VGND VPWR VPWR _22262_/A sky130_fd_sc_hd__buf_2
X_15522_ _15640_/A _15519_/X HADDR[8] _15519_/X VGND VGND VPWR VPWR _24933_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25057__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12734_ _22295_/A VGND VGND VPWR VPWR _12734_/Y sky130_fd_sc_hd__inv_2
X_19290_ _19290_/A VGND VGND VPWR VPWR _19290_/X sky130_fd_sc_hd__buf_2
XFILLER_16_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18241_ _18241_/A VGND VGND VPWR VPWR _18241_/X sky130_fd_sc_hd__buf_2
XFILLER_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15453_ _14269_/X _14239_/A _15426_/X _13907_/B _15447_/X VGND VGND VPWR VPWR _15453_/X
+ sky130_fd_sc_hd__a32o_4
X_12665_ _12597_/A _12670_/B _12641_/X VGND VGND VPWR VPWR _12665_/Y sky130_fd_sc_hd__a21oi_4
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14117_/Y _14398_/X _14403_/X _14398_/X VGND VGND VPWR VPWR _14404_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18172_ _17984_/X _18170_/X _18171_/X VGND VGND VPWR VPWR _18172_/X sky130_fd_sc_hd__and3_4
XFILLER_187_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ _15139_/Y _15383_/X VGND VGND VPWR VPWR _15384_/X sky130_fd_sc_hd__or2_4
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _12657_/A VGND VGND VPWR VPWR _12596_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20517__A _20517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17123_ _17123_/A VGND VGND VPWR VPWR _24385_/D sky130_fd_sc_hd__inv_2
X_14335_ _14329_/A _14339_/B _14314_/X VGND VGND VPWR VPWR _14335_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_117_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17054_ _17019_/Y _17047_/X _17050_/B _17053_/X VGND VGND VPWR VPWR _17054_/X sky130_fd_sc_hd__a211o_4
X_14266_ _23967_/Q VGND VGND VPWR VPWR _14266_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20691__B2 _20690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24692__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16005_ _16003_/Y _15998_/X _16004_/X _15998_/X VGND VGND VPWR VPWR _16005_/X sky130_fd_sc_hd__a2bb2o_4
X_13217_ _13263_/A _13217_/B _13217_/C VGND VGND VPWR VPWR _13217_/X sky130_fd_sc_hd__and3_4
XANTENNA__24621__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14197_ _20517_/B _14188_/X _13785_/X _14190_/X VGND VGND VPWR VPWR _14197_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13148_ _13172_/A _13148_/B _13147_/X VGND VGND VPWR VPWR _13148_/X sky130_fd_sc_hd__and3_4
XANTENNA__21348__A _21348_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15346__A _15331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11874__A RsRx_S1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13079_ _13085_/A _13079_/B _13078_/Y VGND VGND VPWR VPWR _25345_/D sky130_fd_sc_hd__and3_4
X_17956_ _17944_/A _17956_/B VGND VGND VPWR VPWR _17956_/X sky130_fd_sc_hd__or2_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12689__B _12592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16907_ _24705_/Q _16906_/A _16103_/Y _16906_/Y VGND VGND VPWR VPWR _16910_/C sky130_fd_sc_hd__o22a_4
XFILLER_239_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17887_ _17810_/A _17880_/X _17886_/Y VGND VGND VPWR VPWR _24259_/D sky130_fd_sc_hd__and3_4
XFILLER_65_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19626_ _19626_/A VGND VGND VPWR VPWR _19641_/A sky130_fd_sc_hd__inv_2
XFILLER_238_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16838_ _14929_/Y _16834_/X _16597_/X _16837_/X VGND VGND VPWR VPWR _16838_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21083__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25480__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16769_ _16766_/A VGND VGND VPWR VPWR _16769_/X sky130_fd_sc_hd__buf_2
X_19557_ _23695_/Q VGND VGND VPWR VPWR _21950_/B sky130_fd_sc_hd__inv_2
XFILLER_179_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18508_ _18823_/B _18504_/B _18507_/X VGND VGND VPWR VPWR _18509_/A sky130_fd_sc_hd__or3_4
X_19488_ _22010_/B _19482_/X _11911_/X _19487_/X VGND VGND VPWR VPWR _23720_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17375__A1 _17241_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18439_ _16207_/Y _24180_/Q _22548_/A _18400_/Y VGND VGND VPWR VPWR _18439_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21450_ _12833_/C _21446_/X _21449_/X VGND VGND VPWR VPWR _21450_/X sky130_fd_sc_hd__o21a_4
X_20401_ _20389_/A VGND VGND VPWR VPWR _20401_/X sky130_fd_sc_hd__buf_2
XFILLER_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21381_ _21381_/A _22582_/A VGND VGND VPWR VPWR _21381_/X sky130_fd_sc_hd__and2_4
XFILLER_193_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24709__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14425__A _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20332_ _22251_/B _20329_/X _19603_/A _20329_/X VGND VGND VPWR VPWR _23416_/D sky130_fd_sc_hd__a2bb2o_4
X_23120_ _22468_/A VGND VGND VPWR VPWR _23120_/X sky130_fd_sc_hd__buf_2
XFILLER_190_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23051_ _22908_/X _23049_/X _23050_/X _11690_/A _22910_/X VGND VGND VPWR VPWR _23051_/X
+ sky130_fd_sc_hd__a32o_4
X_20263_ _23442_/Q _20262_/Y _23972_/Q _20261_/X VGND VGND VPWR VPWR _20263_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24362__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22002_ _13780_/Y _13804_/Y VGND VGND VPWR VPWR _22395_/A sky130_fd_sc_hd__or2_4
XANTENNA__21258__A _22213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20194_ _23468_/Q VGND VGND VPWR VPWR _21389_/B sky130_fd_sc_hd__inv_2
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24509__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11784__A HWDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23953_ _23951_/CLK sda_i_S4 HRESETn VGND VGND VPWR VPWR _23954_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_229_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_220_0_HCLK clkbuf_7_110_0_HCLK/X VGND VGND VPWR VPWR _24462_/CLK sky130_fd_sc_hd__clkbuf_1
X_22904_ _21533_/A VGND VGND VPWR VPWR _22904_/X sky130_fd_sc_hd__buf_2
X_23884_ _23884_/CLK _23884_/D VGND VGND VPWR VPWR _19020_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22835_ _22835_/A VGND VGND VPWR VPWR _22835_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22766_ _22733_/X _22740_/Y _22766_/C _22766_/D VGND VGND VPWR VPWR HRDATA[15] sky130_fd_sc_hd__or4_4
XFILLER_198_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22817__A _16492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24505_ _24060_/CLK _16653_/X HRESETn VGND VGND VPWR VPWR _24505_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21717_ _14412_/Y _14212_/A _14435_/Y _15457_/A VGND VGND VPWR VPWR _21719_/C sky130_fd_sc_hd__o22a_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25485_ _23938_/CLK _12063_/X HRESETn VGND VGND VPWR VPWR _25485_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22697_ _22515_/X _22695_/X _21956_/A _22696_/Y VGND VGND VPWR VPWR _22697_/X sky130_fd_sc_hd__o22a_4
XFILLER_197_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17533__A1_N _11732_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12450_ _12229_/A _12450_/B VGND VGND VPWR VPWR _12452_/B sky130_fd_sc_hd__or2_4
X_24436_ _24460_/CLK _16812_/X HRESETn VGND VGND VPWR VPWR _14966_/A sky130_fd_sc_hd__dfrtp_4
X_21648_ _21642_/X _21647_/X _13552_/Y _21642_/X VGND VGND VPWR VPWR _21648_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12381_ _12261_/X VGND VGND VPWR VPWR _12415_/A sky130_fd_sc_hd__inv_2
X_24367_ _24365_/CLK _24367_/D HRESETn VGND VGND VPWR VPWR _24367_/Q sky130_fd_sc_hd__dfrtp_4
X_21579_ _15005_/Y _21579_/B VGND VGND VPWR VPWR _21579_/X sky130_fd_sc_hd__and2_4
XFILLER_165_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14120_ _14114_/X _14119_/X _14086_/A _14114_/X VGND VGND VPWR VPWR _25224_/D sky130_fd_sc_hd__a2bb2o_4
X_23318_ _22543_/X _23315_/Y _23155_/X _23317_/X VGND VGND VPWR VPWR _23318_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24298_ _24947_/CLK _17682_/X HRESETn VGND VGND VPWR VPWR _17513_/A sky130_fd_sc_hd__dfrtp_4
X_14051_ _13965_/X VGND VGND VPWR VPWR _14052_/A sky130_fd_sc_hd__inv_2
X_23249_ _24576_/Q _23075_/B _23075_/C VGND VGND VPWR VPWR _23249_/X sky130_fd_sc_hd__and3_4
X_13002_ _12315_/A _13001_/Y VGND VGND VPWR VPWR _13002_/X sky130_fd_sc_hd__or2_4
XANTENNA__21168__A _15666_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24032__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20072__A _20067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_30_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_61_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17810_ _17810_/A VGND VGND VPWR VPWR _17818_/A sky130_fd_sc_hd__buf_2
X_18790_ _18789_/X VGND VGND VPWR VPWR _18791_/B sky130_fd_sc_hd__inv_2
XFILLER_121_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17741_ _17810_/A VGND VGND VPWR VPWR _17790_/A sky130_fd_sc_hd__buf_2
X_14953_ _25025_/Q VGND VGND VPWR VPWR _15214_/B sky130_fd_sc_hd__inv_2
XFILLER_48_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13904_ _24975_/Q _14232_/B _14232_/C _14231_/A VGND VGND VPWR VPWR _13904_/X sky130_fd_sc_hd__or4_4
XANTENNA__17381__A _17239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17672_ _17499_/Y _17671_/X VGND VGND VPWR VPWR _17676_/B sky130_fd_sc_hd__or2_4
X_14884_ _14883_/Y _24445_/Q _14883_/Y _24445_/Q VGND VGND VPWR VPWR _14891_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16623_ RsRx_S0 _16170_/B _16622_/Y VGND VGND VPWR VPWR _16632_/B sky130_fd_sc_hd__o21a_4
X_19411_ _19411_/A _20199_/B _19387_/A _13613_/A VGND VGND VPWR VPWR _19412_/A sky130_fd_sc_hd__or4_4
XANTENNA__16801__B1 _16464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13835_ _25256_/Q VGND VGND VPWR VPWR _21381_/A sky130_fd_sc_hd__inv_2
XANTENNA__22335__D1 _22334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16554_ _16554_/A VGND VGND VPWR VPWR _16554_/Y sky130_fd_sc_hd__inv_2
X_19342_ _19342_/A VGND VGND VPWR VPWR _19343_/A sky130_fd_sc_hd__inv_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12969__A2 _12854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21689__B1 _21501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13766_ _11676_/A _14395_/A VGND VGND VPWR VPWR _14208_/A sky130_fd_sc_hd__or2_4
XFILLER_90_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15505_ _24939_/Q VGND VGND VPWR VPWR _15505_/Y sky130_fd_sc_hd__inv_2
X_12717_ _12717_/A _12721_/B VGND VGND VPWR VPWR _12722_/A sky130_fd_sc_hd__or2_4
X_19273_ _19273_/A VGND VGND VPWR VPWR _20052_/A sky130_fd_sc_hd__buf_2
XANTENNA__21631__A _22380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16485_ _16485_/A VGND VGND VPWR VPWR _16485_/Y sky130_fd_sc_hd__inv_2
X_13697_ _11826_/Y _13677_/B VGND VGND VPWR VPWR _13697_/Y sky130_fd_sc_hd__nand2_4
XFILLER_70_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18224_ _18004_/X _23827_/Q VGND VGND VPWR VPWR _18224_/X sky130_fd_sc_hd__or2_4
X_15436_ _15436_/A _15436_/B VGND VGND VPWR VPWR _15436_/Y sky130_fd_sc_hd__nor2_4
X_12648_ _12648_/A _12639_/X _12648_/C VGND VGND VPWR VPWR _12648_/X sky130_fd_sc_hd__and3_4
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24873__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16127__A1_N _16126_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18155_ _18056_/A _18155_/B _18155_/C VGND VGND VPWR VPWR _18155_/X sky130_fd_sc_hd__and3_4
XFILLER_175_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15367_ _15352_/A _15367_/B _15366_/Y VGND VGND VPWR VPWR _24992_/D sky130_fd_sc_hd__and3_4
XANTENNA__24802__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12579_ _12578_/Y _24858_/Q _12724_/A _12550_/Y VGND VGND VPWR VPWR _12586_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14245__A _14245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17106_ _17103_/A _17103_/B VGND VGND VPWR VPWR _17106_/Y sky130_fd_sc_hd__nand2_4
XFILLER_172_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14318_ _14318_/A _14339_/A VGND VGND VPWR VPWR _14318_/X sky130_fd_sc_hd__or2_4
XFILLER_8_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18086_ _18004_/X _23775_/Q VGND VGND VPWR VPWR _18088_/B sky130_fd_sc_hd__or2_4
X_15298_ _15298_/A _15139_/Y _15409_/A _15087_/Y VGND VGND VPWR VPWR _15298_/X sky130_fd_sc_hd__or4_4
XFILLER_183_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_112_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_112_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17037_ _24384_/Q VGND VGND VPWR VPWR _17038_/C sky130_fd_sc_hd__inv_2
XFILLER_172_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14249_ _25191_/Q VGND VGND VPWR VPWR _14249_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17556__A _17555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16460__A _16453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23277__B _23277_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22181__B _22181_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21078__A _21078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18490__C1 _18489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18988_ _23895_/Q VGND VGND VPWR VPWR _18988_/Y sky130_fd_sc_hd__inv_2
X_17939_ _17934_/X _17938_/X _18020_/A VGND VGND VPWR VPWR _17947_/B sky130_fd_sc_hd__o21a_4
XFILLER_239_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20950_ _20953_/B _13653_/X _20949_/X VGND VGND VPWR VPWR _20950_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19609_ _19609_/A VGND VGND VPWR VPWR _21951_/B sky130_fd_sc_hd__inv_2
XANTENNA__12409__A1 _12194_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20881_ _24047_/Q _13648_/X _20880_/Y VGND VGND VPWR VPWR _20881_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_50_0_HCLK clkbuf_8_51_0_HCLK/A VGND VGND VPWR VPWR _24227_/CLK sky130_fd_sc_hd__clkbuf_1
X_22620_ _22620_/A _22696_/B VGND VGND VPWR VPWR _22620_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13324__A _13388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22551_ _22629_/A _22548_/X _22550_/X VGND VGND VPWR VPWR _22577_/C sky130_fd_sc_hd__and3_4
XFILLER_195_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21502_ _21477_/X _21499_/X _21501_/X VGND VGND VPWR VPWR _21502_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_167_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15966__A1_N _12178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25270_ _24172_/CLK _25270_/D HRESETn VGND VGND VPWR VPWR _13542_/A sky130_fd_sc_hd__dfrtp_4
X_22482_ _22482_/A _22901_/B VGND VGND VPWR VPWR _22482_/X sky130_fd_sc_hd__or2_4
XFILLER_210_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24221_ _23398_/CLK _24221_/D HRESETn VGND VGND VPWR VPWR _23348_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11779__A HWDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21433_ _15851_/X VGND VGND VPWR VPWR _21533_/A sky130_fd_sc_hd__buf_2
XFILLER_148_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18848__B2 _18613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24543__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21364_ _23964_/Q _21364_/B VGND VGND VPWR VPWR _21372_/A sky130_fd_sc_hd__nand2_4
X_24152_ _24148_/CLK _24152_/D HRESETn VGND VGND VPWR VPWR _24152_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22372__A _22365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17520__A1 _25529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20315_ _20310_/X VGND VGND VPWR VPWR _20315_/Y sky130_fd_sc_hd__inv_2
X_23103_ _23103_/A _23102_/X VGND VGND VPWR VPWR _23103_/X sky130_fd_sc_hd__and2_4
XFILLER_162_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15531__B1 HADDR[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21295_ _24894_/Q _21294_/X VGND VGND VPWR VPWR _21295_/X sky130_fd_sc_hd__or2_4
X_24083_ _25113_/CLK _24083_/D HRESETn VGND VGND VPWR VPWR _20437_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20246_ _22198_/B _20243_/X _16858_/X _20243_/X VGND VGND VPWR VPWR _20246_/X sky130_fd_sc_hd__a2bb2o_4
X_23034_ _23011_/X _23015_/X _23034_/C _23033_/X VGND VGND VPWR VPWR HRDATA[22] sky130_fd_sc_hd__or4_4
XFILLER_162_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_17_0_HCLK clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20177_ _20177_/A VGND VGND VPWR VPWR _20177_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21138__D _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24985_ _24985_/CLK _24985_/D HRESETn VGND VGND VPWR VPWR _15106_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_245_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15714__A _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25331__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11950_ _11950_/A VGND VGND VPWR VPWR _11951_/A sky130_fd_sc_hd__inv_2
X_23936_ _23932_/CLK _20986_/A HRESETn VGND VGND VPWR VPWR _20987_/C sky130_fd_sc_hd__dfstp_4
XANTENNA__21435__B _23002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18728__C _18745_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22580__A1 _24425_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11881_ _11881_/A VGND VGND VPWR VPWR _11881_/Y sky130_fd_sc_hd__inv_2
X_23867_ _23853_/CLK _23867_/D VGND VGND VPWR VPWR _23867_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_232_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13620_ _13579_/X _13588_/X _13620_/C _13620_/D VGND VGND VPWR VPWR _13620_/X sky130_fd_sc_hd__or4_4
XFILLER_189_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13234__A _13421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22818_ _16576_/A _22730_/X _22533_/X _22817_/X VGND VGND VPWR VPWR _22818_/X sky130_fd_sc_hd__a211o_4
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23798_ _23806_/CLK _23798_/D VGND VGND VPWR VPWR _23798_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__22332__A1 _22331_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18536__B1 _18489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13551_ _13543_/X _13545_/X _13548_/X _13550_/X VGND VGND VPWR VPWR _13575_/B sky130_fd_sc_hd__or4_4
X_25537_ _24310_/CLK _25537_/D HRESETn VGND VGND VPWR VPWR _25537_/Q sky130_fd_sc_hd__dfrtp_4
X_22749_ _21294_/X _22748_/X _21300_/A _24835_/Q _22490_/X VGND VGND VPWR VPWR _22749_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_197_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12820__B2 _24789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12502_ _24861_/Q VGND VGND VPWR VPWR _12502_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16270_ _16270_/A _16270_/B VGND VGND VPWR VPWR _16270_/X sky130_fd_sc_hd__or2_4
XFILLER_186_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21170__B _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13482_ _16181_/A _13482_/B VGND VGND VPWR VPWR _13483_/D sky130_fd_sc_hd__or2_4
X_25468_ _25109_/CLK _25468_/D HRESETn VGND VGND VPWR VPWR _18372_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_9_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20067__A _20067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21601__D _21600_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15221_ _15221_/A VGND VGND VPWR VPWR _15221_/Y sky130_fd_sc_hd__inv_2
X_12433_ _12187_/Y _12433_/B VGND VGND VPWR VPWR _12433_/Y sky130_fd_sc_hd__nand2_4
X_24419_ _24419_/CLK _24419_/D HRESETn VGND VGND VPWR VPWR _14940_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24284__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25399_ _25397_/CLK _25399_/D HRESETn VGND VGND VPWR VPWR _25399_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18760__A _18760_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20646__A1 _14229_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15152_ _15288_/A _15140_/Y _15139_/Y _24584_/Q VGND VGND VPWR VPWR _15156_/C sky130_fd_sc_hd__a2bb2o_4
X_12364_ _25363_/Q _12352_/Y _13069_/A _24824_/Q VGND VGND VPWR VPWR _12364_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24213__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22282__A _22282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14103_ _14088_/C _14102_/X _14103_/C VGND VGND VPWR VPWR _14103_/X sky130_fd_sc_hd__or3_4
X_15083_ _15295_/A _15081_/Y _15082_/Y _24606_/Q VGND VGND VPWR VPWR _15089_/B sky130_fd_sc_hd__a2bb2o_4
X_19960_ _18279_/A VGND VGND VPWR VPWR _19960_/X sky130_fd_sc_hd__buf_2
XANTENNA__15522__B1 HADDR[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12295_ _12980_/A _12293_/Y _13005_/A _24846_/Q VGND VGND VPWR VPWR _12295_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_181_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14034_ _14034_/A _14033_/X _14034_/C _13981_/X VGND VGND VPWR VPWR _14034_/X sky130_fd_sc_hd__or4_4
X_18911_ _19209_/A _18911_/B _19047_/C VGND VGND VPWR VPWR _18911_/X sky130_fd_sc_hd__or3_4
X_19891_ _19878_/Y VGND VGND VPWR VPWR _19891_/X sky130_fd_sc_hd__buf_2
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18842_ _24574_/Q _18698_/A _16534_/Y _18641_/A VGND VGND VPWR VPWR _18842_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15985_ _16366_/A _15985_/B VGND VGND VPWR VPWR _16270_/B sky130_fd_sc_hd__or2_4
X_18773_ _18773_/A VGND VGND VPWR VPWR _24140_/D sky130_fd_sc_hd__inv_2
XFILLER_0_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13836__B1 _13521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25072__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14936_ _14936_/A VGND VGND VPWR VPWR _14936_/Y sky130_fd_sc_hd__inv_2
X_17724_ _22257_/A VGND VGND VPWR VPWR _17725_/A sky130_fd_sc_hd__buf_2
XFILLER_76_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21374__A2 _21356_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15135__A2_N _24595_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25001__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14867_ _14859_/B _14866_/X VGND VGND VPWR VPWR _14867_/Y sky130_fd_sc_hd__nor2_4
X_17655_ _17627_/A VGND VGND VPWR VPWR _17682_/A sky130_fd_sc_hd__buf_2
XANTENNA__16681__A1_N _16679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_37_0_HCLK clkbuf_7_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_74_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13818_ _15965_/A VGND VGND VPWR VPWR _13818_/X sky130_fd_sc_hd__buf_2
X_16606_ _16598_/A VGND VGND VPWR VPWR _16606_/X sky130_fd_sc_hd__buf_2
X_17586_ _17614_/A _17516_/Y _17597_/A _17585_/X VGND VGND VPWR VPWR _17586_/X sky130_fd_sc_hd__or4_4
XFILLER_223_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14798_ _14812_/C _14797_/X _14798_/C VGND VGND VPWR VPWR _14798_/X sky130_fd_sc_hd__or3_4
XFILLER_16_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22457__A _21587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16537_ _16536_/Y _16454_/A _16361_/X _16454_/A VGND VGND VPWR VPWR _16537_/X sky130_fd_sc_hd__a2bb2o_4
X_19325_ _19324_/Y _19322_/X _19279_/X _19322_/X VGND VGND VPWR VPWR _19325_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13749_ _25279_/Q VGND VGND VPWR VPWR _20157_/D sky130_fd_sc_hd__buf_2
XFILLER_177_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16468_ _16466_/Y _16461_/X _16467_/X _16461_/X VGND VGND VPWR VPWR _16468_/X sky130_fd_sc_hd__a2bb2o_4
X_19256_ _23801_/Q VGND VGND VPWR VPWR _22214_/B sky130_fd_sc_hd__inv_2
XFILLER_176_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15419_ _15087_/Y _15320_/D _15313_/A _15417_/B VGND VGND VPWR VPWR _15419_/X sky130_fd_sc_hd__a211o_4
X_18207_ _17972_/A _18207_/B VGND VGND VPWR VPWR _18207_/X sky130_fd_sc_hd__or2_4
XFILLER_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19187_ _19183_/Y _19186_/X _19144_/X _19186_/X VGND VGND VPWR VPWR _23826_/D sky130_fd_sc_hd__a2bb2o_4
X_16399_ _15091_/Y _16393_/X _16397_/X _16398_/X VGND VGND VPWR VPWR _24599_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_3_6_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18138_ _18032_/A _18138_/B VGND VGND VPWR VPWR _18138_/X sky130_fd_sc_hd__or2_4
XFILLER_8_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18069_ _18032_/A _19308_/A VGND VGND VPWR VPWR _18069_/X sky130_fd_sc_hd__or2_4
XANTENNA__17286__A _17284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15513__B1 HADDR[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20100_ _21898_/B _20096_/X _20099_/X _20096_/X VGND VGND VPWR VPWR _23503_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21080_ _22756_/B VGND VGND VPWR VPWR _21080_/X sky130_fd_sc_hd__buf_2
XFILLER_144_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20031_ _20031_/A VGND VGND VPWR VPWR _20031_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13827__B1 _13826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18645__A2_N _24138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24770_ _24765_/CLK _24770_/D HRESETn VGND VGND VPWR VPWR _12247_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19006__A _19006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21982_ _21983_/A _20318_/X _18350_/Y _23420_/Q VGND VGND VPWR VPWR _21982_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23721_ _23406_/CLK _23721_/D VGND VGND VPWR VPWR _23721_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20933_ _24059_/Q _20932_/B _20932_/Y VGND VGND VPWR VPWR _20933_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_199_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23652_ _24209_/CLK _23652_/D VGND VGND VPWR VPWR _13404_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ _16696_/Y _20846_/X _20855_/X _20863_/Y VGND VGND VPWR VPWR _20864_/X sky130_fd_sc_hd__o22a_4
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24795__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22603_ _22149_/X _22602_/X _22134_/A _25531_/Q _22554_/X VGND VGND VPWR VPWR _22603_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21271__A _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23583_ _23555_/CLK _23583_/D VGND VGND VPWR VPWR _23583_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12893__A _12813_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20325__B1 _19759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24724__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20795_ _20780_/X _20794_/Y _15572_/A _20784_/X VGND VGND VPWR VPWR _20795_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16365__A _16365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12802__B2 _24800_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25322_ _25158_/CLK _25322_/D HRESETn VGND VGND VPWR VPWR _13468_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_168_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22534_ _22431_/X VGND VGND VPWR VPWR _22534_/X sky130_fd_sc_hd__buf_2
XFILLER_167_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25253_ _24958_/CLK _13848_/X HRESETn VGND VGND VPWR VPWR _20476_/A sky130_fd_sc_hd__dfrtp_4
X_22465_ _21597_/X VGND VGND VPWR VPWR _22468_/A sky130_fd_sc_hd__buf_2
XANTENNA__22617__A2 _21031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24204_ _23456_/CLK _18348_/X HRESETn VGND VGND VPWR VPWR _13247_/A sky130_fd_sc_hd__dfrtp_4
X_21416_ _21178_/X _21400_/X _21415_/X VGND VGND VPWR VPWR _21416_/X sky130_fd_sc_hd__and3_4
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25184_ _23972_/CLK _14274_/X HRESETn VGND VGND VPWR VPWR _25184_/Q sky130_fd_sc_hd__dfrtp_4
X_22396_ _23690_/Q _22396_/B VGND VGND VPWR VPWR _22396_/X sky130_fd_sc_hd__or2_4
XFILLER_191_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24135_ _24148_/CLK _18801_/X HRESETn VGND VGND VPWR VPWR _24135_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15504__B1 HADDR[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21347_ _21347_/A _22181_/B VGND VGND VPWR VPWR _21347_/X sky130_fd_sc_hd__and2_4
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12080_ _25478_/Q VGND VGND VPWR VPWR _12080_/Y sky130_fd_sc_hd__inv_2
X_24066_ _24049_/CLK _24066_/D HRESETn VGND VGND VPWR VPWR _13655_/A sky130_fd_sc_hd__dfrtp_4
X_21278_ _13779_/X VGND VGND VPWR VPWR _21278_/X sky130_fd_sc_hd__buf_2
XFILLER_89_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23017_ _12240_/Y _23268_/A _23016_/X VGND VGND VPWR VPWR _23017_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_150_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25512__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20229_ _23455_/Q VGND VGND VPWR VPWR _20229_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21446__A _21019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17009__B1 _24717_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15770_ _19646_/A VGND VGND VPWR VPWR _15770_/X sky130_fd_sc_hd__buf_2
XFILLER_218_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21165__B _11700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12982_ _12982_/A VGND VGND VPWR VPWR _13068_/C sky130_fd_sc_hd__inv_2
X_24968_ _24073_/CLK _24968_/D HRESETn VGND VGND VPWR VPWR _13930_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_58_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14721_ _14720_/Y _14702_/X _14720_/A _14701_/A VGND VGND VPWR VPWR _14721_/X sky130_fd_sc_hd__o22a_4
XFILLER_217_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11933_ _11932_/X VGND VGND VPWR VPWR _11934_/B sky130_fd_sc_hd__inv_2
X_23919_ _23912_/CLK _23919_/D VGND VGND VPWR VPWR _18920_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_91_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24899_ _24900_/CLK _24899_/D HRESETn VGND VGND VPWR VPWR _15618_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18755__A _18760_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17440_ _17440_/A VGND VGND VPWR VPWR _17440_/X sky130_fd_sc_hd__buf_2
X_14652_ _19002_/B _19026_/C _19026_/D _19320_/A VGND VGND VPWR VPWR _14652_/X sky130_fd_sc_hd__and4_4
X_11864_ _11863_/Y _11864_/B VGND VGND VPWR VPWR _11864_/X sky130_fd_sc_hd__or2_4
XFILLER_205_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _18095_/A VGND VGND VPWR VPWR _18060_/A sky130_fd_sc_hd__buf_2
X_17371_ _17345_/A _17345_/B _17284_/X _17369_/B VGND VGND VPWR VPWR _17372_/A sky130_fd_sc_hd__a211o_4
XPHY_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _13563_/Y _14555_/X VGND VGND VPWR VPWR _14583_/Y sky130_fd_sc_hd__nand2_4
XFILLER_232_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24465__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ _11790_/Y _11778_/X _11793_/X _11794_/X VGND VGND VPWR VPWR _11795_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19182__B1 _19138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16322_ _24627_/Q VGND VGND VPWR VPWR _16322_/Y sky130_fd_sc_hd__inv_2
X_19110_ _19108_/Y _19109_/X _19063_/X _19109_/X VGND VGND VPWR VPWR _23853_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13534_ _13533_/Y _14547_/A _13533_/Y _14547_/A VGND VGND VPWR VPWR _13541_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19041_ _19039_/Y _19040_/X _18948_/X _19040_/X VGND VGND VPWR VPWR _19041_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16253_ _16251_/Y _16252_/X _16059_/X _16252_/X VGND VGND VPWR VPWR _16253_/X sky130_fd_sc_hd__a2bb2o_4
X_13465_ _13461_/Y _13464_/X _11761_/X _13464_/X VGND VGND VPWR VPWR _13465_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23266__C1 _23265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15204_ _15204_/A _15204_/B _15059_/X _15242_/B VGND VGND VPWR VPWR _15205_/C sky130_fd_sc_hd__or4_4
X_12416_ _12416_/A VGND VGND VPWR VPWR _12416_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16184_ _16183_/Y VGND VGND VPWR VPWR _16184_/X sky130_fd_sc_hd__buf_2
X_13396_ _13396_/A _23908_/Q VGND VGND VPWR VPWR _13397_/C sky130_fd_sc_hd__or2_4
XFILLER_127_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15135_ _15356_/A _24595_/Q _15356_/A _24595_/Q VGND VGND VPWR VPWR _15136_/D sky130_fd_sc_hd__a2bb2o_4
X_12347_ _12976_/C _24835_/Q _12976_/C _24835_/Q VGND VGND VPWR VPWR _12347_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15619__A _14403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15066_ _15066_/A _15065_/X VGND VGND VPWR VPWR _15067_/B sky130_fd_sc_hd__or2_4
X_19943_ _19943_/A VGND VGND VPWR VPWR _19943_/Y sky130_fd_sc_hd__inv_2
X_12278_ _12278_/A _12277_/X VGND VGND VPWR VPWR _12279_/B sky130_fd_sc_hd__or2_4
XFILLER_153_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14017_ _13986_/X _13987_/X _13995_/A VGND VGND VPWR VPWR _14017_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__25253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19874_ _19874_/A VGND VGND VPWR VPWR _19874_/X sky130_fd_sc_hd__buf_2
XFILLER_150_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18996__B1 _18951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18825_ pwm_S7 VGND VGND VPWR VPWR _18825_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23274__C _23266_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18756_ _18693_/C _18755_/X _18709_/X VGND VGND VPWR VPWR _18756_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24089__D _20961_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15968_ _15930_/Y VGND VGND VPWR VPWR _15968_/X sky130_fd_sc_hd__buf_2
XFILLER_208_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14482__B1 _14389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22544__B2 _21317_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17707_ _24213_/Q VGND VGND VPWR VPWR _17707_/X sky130_fd_sc_hd__buf_2
XFILLER_208_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14919_ _14909_/X _14919_/B _14915_/X _14919_/D VGND VGND VPWR VPWR _14935_/C sky130_fd_sc_hd__or4_4
X_15899_ _15701_/X _15887_/X _15764_/X _24788_/Q _15857_/A VGND VGND VPWR VPWR _15899_/X
+ sky130_fd_sc_hd__a32o_4
X_18687_ _24139_/Q VGND VGND VPWR VPWR _18778_/A sky130_fd_sc_hd__inv_2
X_17638_ _17569_/C _17638_/B VGND VGND VPWR VPWR _17648_/B sky130_fd_sc_hd__or2_4
XFILLER_17_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17569_ _17569_/A _17648_/A _17569_/C _17569_/D VGND VGND VPWR VPWR _17569_/X sky130_fd_sc_hd__or4_4
XANTENNA__22847__A2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19173__B1 _19057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19308_ _19308_/A VGND VGND VPWR VPWR _19308_/Y sky130_fd_sc_hd__inv_2
X_20580_ _23945_/Q _20580_/B VGND VGND VPWR VPWR _20580_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24135__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_124_0_HCLK clkbuf_7_62_0_HCLK/X VGND VGND VPWR VPWR _24866_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_187_0_HCLK clkbuf_7_93_0_HCLK/X VGND VGND VPWR VPWR _23932_/CLK sky130_fd_sc_hd__clkbuf_1
X_19239_ _22058_/B _19233_/X _16869_/X _19238_/X VGND VGND VPWR VPWR _19239_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15734__B1 _11721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20820__A1_N _20690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16913__A _16913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22250_ _21453_/X _22242_/X _22249_/X VGND VGND VPWR VPWR _22250_/X sky130_fd_sc_hd__and3_4
XFILLER_192_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21201_ _21209_/A _21201_/B VGND VGND VPWR VPWR _21202_/C sky130_fd_sc_hd__or2_4
X_22181_ _25250_/Q _22181_/B VGND VGND VPWR VPWR _22181_/X sky130_fd_sc_hd__and2_4
XFILLER_145_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21132_ _17438_/B VGND VGND VPWR VPWR _21132_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23024__A2 _22838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22650__A _22618_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21063_ _22136_/B VGND VGND VPWR VPWR _21109_/A sky130_fd_sc_hd__buf_2
XFILLER_235_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22232__B1 _21178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17744__A _17744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20014_ _22340_/B _20013_/X _19964_/X _20013_/X VGND VGND VPWR VPWR _23538_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18987__B1 _18985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11792__A _13797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24822_ _25428_/CLK _24822_/D HRESETn VGND VGND VPWR VPWR _24822_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24976__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16588__A1_N _16587_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14473__B1 _14392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25301__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16079__B _15670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24753_ _24753_/CLK _15973_/X HRESETn VGND VGND VPWR VPWR _22150_/A sky130_fd_sc_hd__dfrtp_4
X_21965_ _21968_/A _23686_/Q _25081_/Q _19589_/Y VGND VGND VPWR VPWR _21965_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24905__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23704_ _23706_/CLK _23704_/D VGND VGND VPWR VPWR _23704_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _20916_/A _20916_/B VGND VGND VPWR VPWR _20916_/X sky130_fd_sc_hd__and2_4
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24684_ _24704_/CLK _16158_/X HRESETn VGND VGND VPWR VPWR _21698_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_82_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21896_ _22069_/A VGND VGND VPWR VPWR _21896_/X sky130_fd_sc_hd__buf_2
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_20_0_HCLK clkbuf_7_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_20_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _23644_/CLK _19736_/X VGND VGND VPWR VPWR _13443_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _13644_/A VGND VGND VPWR VPWR _20847_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15973__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_83_0_HCLK clkbuf_7_83_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_83_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23566_ _23555_/CLK _19930_/X VGND VGND VPWR VPWR _19929_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20778_ _13108_/B _20771_/X _20777_/X VGND VGND VPWR VPWR _20778_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20313__A3 _13829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25305_ _25308_/CLK _13517_/X HRESETn VGND VGND VPWR VPWR SCLK_S2 sky130_fd_sc_hd__dfstp_4
XFILLER_167_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22517_ _22517_/A _22696_/B VGND VGND VPWR VPWR _22517_/Y sky130_fd_sc_hd__nor2_4
XFILLER_7_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23497_ _23497_/CLK _20119_/X VGND VGND VPWR VPWR _20118_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_127_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ _13389_/A _19100_/A VGND VGND VPWR VPWR _13251_/C sky130_fd_sc_hd__or2_4
X_25236_ _23976_/CLK _14068_/X HRESETn VGND VGND VPWR VPWR _25236_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22448_ _21319_/X VGND VGND VPWR VPWR _22876_/C sky130_fd_sc_hd__buf_2
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15740__A3 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12201_ _12201_/A VGND VGND VPWR VPWR _12201_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13181_ _13353_/A _13173_/X _13180_/X _11948_/A _11948_/B VGND VGND VPWR VPWR _13181_/X
+ sky130_fd_sc_hd__o32a_4
X_25167_ _25164_/CLK _25167_/D HRESETn VGND VGND VPWR VPWR _18372_/B sky130_fd_sc_hd__dfstp_4
X_22379_ _22379_/A _20031_/Y VGND VGND VPWR VPWR _22379_/X sky130_fd_sc_hd__or2_4
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12132_ _12097_/A _12131_/Y _12097_/A _12131_/Y VGND VGND VPWR VPWR _12132_/X sky130_fd_sc_hd__a2bb2o_4
X_24118_ _25100_/CLK _24118_/D HRESETn VGND VGND VPWR VPWR _20992_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25098_ _25098_/CLK _14565_/X HRESETn VGND VGND VPWR VPWR _25098_/Q sky130_fd_sc_hd__dfrtp_4
X_12063_ _12062_/Y _12060_/X _11765_/X _12060_/X VGND VGND VPWR VPWR _12063_/X sky130_fd_sc_hd__a2bb2o_4
X_16940_ _24280_/Q VGND VGND VPWR VPWR _16940_/Y sky130_fd_sc_hd__inv_2
X_24049_ _24049_/CLK _24049_/D HRESETn VGND VGND VPWR VPWR _20889_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18978__B1 _17415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21176__A _21176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16871_ _20102_/A VGND VGND VPWR VPWR _19820_/A sky130_fd_sc_hd__buf_2
XANTENNA__12798__A _25385_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22986__A1_N _17249_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18610_ _18610_/A VGND VGND VPWR VPWR _18789_/C sky130_fd_sc_hd__buf_2
XFILLER_219_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15822_ _12319_/Y _15820_/X _15752_/X _15820_/X VGND VGND VPWR VPWR _15822_/X sky130_fd_sc_hd__a2bb2o_4
X_19590_ _19576_/A VGND VGND VPWR VPWR _19590_/X sky130_fd_sc_hd__buf_2
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14464__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15753_ _12537_/Y _15750_/X _15752_/X _15750_/X VGND VGND VPWR VPWR _24864_/D sky130_fd_sc_hd__a2bb2o_4
X_18541_ _18523_/X _18541_/B _18540_/Y VGND VGND VPWR VPWR _24176_/D sky130_fd_sc_hd__and3_4
XANTENNA__21904__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12965_ _12967_/A _12959_/B _12965_/C VGND VGND VPWR VPWR _12965_/X sky130_fd_sc_hd__and3_4
XANTENNA__24646__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11916_ _11914_/Y _11907_/X _11915_/X _11907_/X VGND VGND VPWR VPWR _11916_/X sky130_fd_sc_hd__a2bb2o_4
X_14704_ _14704_/A VGND VGND VPWR VPWR _14704_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15684_ _15673_/X _15680_/A _15694_/A _15675_/Y _15683_/X VGND VGND VPWR VPWR _15684_/X
+ sky130_fd_sc_hd__a32o_4
X_18472_ _24161_/Q VGND VGND VPWR VPWR _18589_/A sky130_fd_sc_hd__inv_2
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12896_ _12836_/Y _12896_/B VGND VGND VPWR VPWR _12897_/C sky130_fd_sc_hd__or2_4
XANTENNA__14216__B1 _13826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14635_ _18090_/A VGND VGND VPWR VPWR _14636_/A sky130_fd_sc_hd__buf_2
X_17423_ _17420_/Y _17414_/X _17421_/X _17422_/X VGND VGND VPWR VPWR _24331_/D sky130_fd_sc_hd__a2bb2o_4
X_11847_ _11813_/X _11847_/B _11835_/X _11846_/X VGND VGND VPWR VPWR _11934_/C sky130_fd_sc_hd__or4_4
XFILLER_205_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13422__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14563_/A _14563_/B _14563_/C _14566_/D VGND VGND VPWR VPWR _14566_/X sky130_fd_sc_hd__and4_4
X_17354_ _17354_/A VGND VGND VPWR VPWR _17354_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11682_/Y VGND VGND VPWR VPWR _11778_/X sky130_fd_sc_hd__buf_2
XFILLER_158_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13517_ _20964_/B _13516_/X SCLK_S2 _20964_/B VGND VGND VPWR VPWR _13517_/X sky130_fd_sc_hd__a2bb2o_4
X_16305_ _24633_/Q VGND VGND VPWR VPWR _16305_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17285_ _17254_/X _17264_/X _17255_/A VGND VGND VPWR VPWR _17285_/X sky130_fd_sc_hd__o21a_4
XFILLER_147_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15716__B1 _15560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14497_ _14492_/B VGND VGND VPWR VPWR _14497_/Y sky130_fd_sc_hd__inv_2
X_16236_ _16236_/A VGND VGND VPWR VPWR _16236_/X sky130_fd_sc_hd__buf_2
X_19024_ _19024_/A VGND VGND VPWR VPWR _19024_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13448_ _13310_/X _13444_/X _13448_/C VGND VGND VPWR VPWR _13448_/X sky130_fd_sc_hd__or3_4
XANTENNA__23254__A2 _21031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20255__A _20243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16452__B _16540_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16167_ _16166_/X VGND VGND VPWR VPWR _16167_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13379_ _13312_/A _13379_/B VGND VGND VPWR VPWR _13380_/C sky130_fd_sc_hd__or2_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15118_ _15405_/A VGND VGND VPWR VPWR _15298_/A sky130_fd_sc_hd__inv_2
XFILLER_114_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16098_ _23157_/A VGND VGND VPWR VPWR _16098_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15049_ _15049_/A _15049_/B _15045_/X _15048_/X VGND VGND VPWR VPWR _15049_/X sky130_fd_sc_hd__or4_4
X_19926_ _19924_/Y _19920_/X _19606_/X _19925_/X VGND VGND VPWR VPWR _19926_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18969__B1 _18948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21086__A _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19857_ _19856_/Y VGND VGND VPWR VPWR _19857_/X sky130_fd_sc_hd__buf_2
X_18808_ _18788_/B _18812_/B VGND VGND VPWR VPWR _18808_/Y sky130_fd_sc_hd__nand2_4
XFILLER_205_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19788_ _23616_/Q VGND VGND VPWR VPWR _19788_/Y sky130_fd_sc_hd__inv_2
XFILLER_228_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15798__A3 _15719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18739_ _18739_/A _18738_/Y VGND VGND VPWR VPWR _18739_/X sky130_fd_sc_hd__or2_4
XFILLER_37_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24387__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16908__A _24265_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21750_ _21119_/X _21748_/Y _21596_/X _21749_/X VGND VGND VPWR VPWR _21750_/X sky130_fd_sc_hd__o22a_4
XFILLER_70_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24316__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18615__A1_N _16566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21740__A2 _15704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20701_ _20700_/Y _13112_/A _13113_/X VGND VGND VPWR VPWR _20701_/X sky130_fd_sc_hd__o21a_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21681_ _21487_/A _21681_/B VGND VGND VPWR VPWR _21682_/C sky130_fd_sc_hd__or2_4
XFILLER_211_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23420_ _23425_/CLK _20321_/X VGND VGND VPWR VPWR _23420_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12874__C _12588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20632_ _15462_/Y _20615_/X _20629_/X _20631_/X VGND VGND VPWR VPWR _20632_/X sky130_fd_sc_hd__a211o_4
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23351_ _11699_/A _15724_/A HWDATA[26] _25546_/Q _11681_/X VGND VGND VPWR VPWR _25546_/D
+ sky130_fd_sc_hd__a32o_4
X_20563_ _18875_/X _20563_/B _20553_/C VGND VGND VPWR VPWR _20563_/X sky130_fd_sc_hd__and3_4
XFILLER_50_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16643__A _16655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22302_ _25374_/Q _22299_/X _22301_/X VGND VGND VPWR VPWR _22302_/X sky130_fd_sc_hd__a21o_4
X_23282_ _21520_/X _23281_/X _21522_/X _15993_/A _23152_/X VGND VGND VPWR VPWR _23282_/X
+ sky130_fd_sc_hd__a32o_4
X_20494_ _20479_/A VGND VGND VPWR VPWR _20495_/C sky130_fd_sc_hd__buf_2
XANTENNA__12890__B _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15722__A3 _15721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23951__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25021_ _25021_/CLK _25021_/D HRESETn VGND VGND VPWR VPWR _25021_/Q sky130_fd_sc_hd__dfrtp_4
X_22233_ _21274_/X _22213_/X _22228_/X _22231_/Y _22232_/X VGND VGND VPWR VPWR _22233_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__22453__B1 _14911_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25104__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22164_ _16520_/A _21309_/X _21339_/X VGND VGND VPWR VPWR _22164_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16132__B1 _11739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22380__A _22380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21115_ _17239_/A _21111_/X _21114_/X VGND VGND VPWR VPWR _21115_/X sky130_fd_sc_hd__o21a_4
XFILLER_160_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22095_ _23091_/A _22095_/B _22095_/C VGND VGND VPWR VPWR _22095_/X sky130_fd_sc_hd__and3_4
X_21046_ _21041_/X _21045_/Y _12968_/A _21041_/X VGND VGND VPWR VPWR _21046_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_219_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14446__B1 _14403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24805_ _24804_/CLK _24805_/D HRESETn VGND VGND VPWR VPWR _24805_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_216_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22997_ _24568_/Q _22885_/X _22802_/X VGND VGND VPWR VPWR _22997_/X sky130_fd_sc_hd__o21a_4
XANTENNA__19385__B1 _19295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12750_ _12749_/Y _24785_/Q _12749_/Y _24785_/Q VGND VGND VPWR VPWR _12751_/D sky130_fd_sc_hd__a2bb2o_4
X_24736_ _24737_/CLK _16023_/X HRESETn VGND VGND VPWR VPWR _24736_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21948_ _21926_/A _21948_/B VGND VGND VPWR VPWR _21948_/X sky130_fd_sc_hd__or2_4
XFILLER_131_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16199__B1 _15567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24057__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _21327_/A VGND VGND VPWR VPWR _11701_/X sky130_fd_sc_hd__buf_2
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12681_/A _12681_/B VGND VGND VPWR VPWR _12681_/X sky130_fd_sc_hd__or2_4
X_24667_ _24667_/CLK _16213_/X HRESETn VGND VGND VPWR VPWR _22939_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_188_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21879_ _21019_/X VGND VGND VPWR VPWR _21879_/X sky130_fd_sc_hd__buf_2
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14419_/Y _14415_/X _14389_/X _14408_/A VGND VGND VPWR VPWR _14420_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _23458_/CLK _23618_/D VGND VGND VPWR VPWR _23618_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24598_ _24551_/CLK _16401_/X HRESETn VGND VGND VPWR VPWR _24598_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22108__A2_N _21721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _25159_/Q _14340_/X _25158_/Q _14345_/X VGND VGND VPWR VPWR _14351_/X sky130_fd_sc_hd__o22a_4
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23549_ _24317_/CLK _19982_/X VGND VGND VPWR VPWR _19979_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13434_/A _13302_/B _13302_/C VGND VGND VPWR VPWR _13302_/X sky130_fd_sc_hd__and3_4
XFILLER_183_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17070_ _17070_/A _17070_/B _17070_/C VGND VGND VPWR VPWR _24400_/D sky130_fd_sc_hd__and3_4
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _13508_/D _14281_/Y _14290_/A VGND VGND VPWR VPWR _25182_/D sky130_fd_sc_hd__o21a_4
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_170_0_HCLK clkbuf_7_85_0_HCLK/X VGND VGND VPWR VPWR _24088_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16371__B1 _15991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16021_ _16018_/Y _16019_/X _16020_/X _16019_/X VGND VGND VPWR VPWR _16021_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13233_ _13438_/A _13233_/B VGND VGND VPWR VPWR _13233_/X sky130_fd_sc_hd__or2_4
X_25219_ _25113_/CLK _25219_/D HRESETn VGND VGND VPWR VPWR _14105_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_27_0_HCLK clkbuf_8_26_0_HCLK/A VGND VGND VPWR VPWR _24297_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13164_ _13263_/A _13151_/X _13163_/X VGND VGND VPWR VPWR _13164_/X sky130_fd_sc_hd__or3_4
XFILLER_156_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22290__A _22290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12115_ _12115_/A _12125_/A VGND VGND VPWR VPWR _12129_/A sky130_fd_sc_hd__and2_4
XFILLER_123_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17871__B1 _16952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13095_ _12321_/Y _13095_/B VGND VGND VPWR VPWR _13097_/B sky130_fd_sc_hd__or2_4
X_17972_ _17972_/A _23761_/Q VGND VGND VPWR VPWR _17973_/C sky130_fd_sc_hd__or2_4
XANTENNA__24898__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19711_ _19360_/A VGND VGND VPWR VPWR _19711_/X sky130_fd_sc_hd__buf_2
X_12046_ _13462_/C _12058_/B _12160_/C _13457_/D VGND VGND VPWR VPWR _12047_/A sky130_fd_sc_hd__or4_4
X_16923_ _16923_/A VGND VGND VPWR VPWR _17752_/C sky130_fd_sc_hd__inv_2
XANTENNA__24827__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19642_ _19640_/Y _19641_/X _19540_/X _19641_/X VGND VGND VPWR VPWR _19642_/X sky130_fd_sc_hd__a2bb2o_4
X_16854_ _24413_/Q VGND VGND VPWR VPWR _16854_/X sky130_fd_sc_hd__buf_2
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15805_ _12354_/Y _15803_/X _11711_/X _15803_/X VGND VGND VPWR VPWR _24840_/D sky130_fd_sc_hd__a2bb2o_4
X_19573_ _22229_/B VGND VGND VPWR VPWR _19573_/X sky130_fd_sc_hd__buf_2
XFILLER_19_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24480__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13997_ _14028_/B _13978_/X _13979_/X _14019_/D VGND VGND VPWR VPWR _13997_/X sky130_fd_sc_hd__or4_4
X_16785_ _15005_/Y _16779_/X _16435_/X _16779_/X VGND VGND VPWR VPWR _16785_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_219_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18524_ _18560_/A _18479_/X VGND VGND VPWR VPWR _18524_/X sky130_fd_sc_hd__or2_4
XFILLER_65_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12948_ _12948_/A _12948_/B VGND VGND VPWR VPWR _12952_/B sky130_fd_sc_hd__or2_4
X_15736_ _15736_/A VGND VGND VPWR VPWR _15736_/X sky130_fd_sc_hd__buf_2
XFILLER_34_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18455_ _18774_/A VGND VGND VPWR VPWR _18580_/A sky130_fd_sc_hd__buf_2
X_12879_ _12879_/A _12879_/B VGND VGND VPWR VPWR _12880_/C sky130_fd_sc_hd__or2_4
X_15667_ _21323_/A VGND VGND VPWR VPWR _22530_/A sky130_fd_sc_hd__buf_2
XANTENNA__20930__B1 _20855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _17384_/X _17398_/X _21000_/B _24336_/Q _17401_/X VGND VGND VPWR VPWR _17406_/X
+ sky130_fd_sc_hd__a32o_4
X_14618_ _14614_/Y _14617_/Y _14613_/X _14616_/X VGND VGND VPWR VPWR _25082_/D sky130_fd_sc_hd__o22a_4
XFILLER_178_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15598_ _24907_/Q VGND VGND VPWR VPWR _15598_/Y sky130_fd_sc_hd__inv_2
X_18386_ _18373_/Y VGND VGND VPWR VPWR _18386_/X sky130_fd_sc_hd__buf_2
XFILLER_187_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14549_ _14549_/A _14549_/B VGND VGND VPWR VPWR _14550_/B sky130_fd_sc_hd__or2_4
X_17337_ _17245_/Y _17335_/A VGND VGND VPWR VPWR _17337_/X sky130_fd_sc_hd__or2_4
XANTENNA__17559__A _24714_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17268_ _17284_/A VGND VGND VPWR VPWR _17268_/X sky130_fd_sc_hd__buf_2
XANTENNA__16362__B1 _16361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19007_ _19000_/Y _19004_/X _19006_/X _19004_/X VGND VGND VPWR VPWR _23890_/D sky130_fd_sc_hd__a2bb2o_4
X_16219_ _22814_/A VGND VGND VPWR VPWR _16219_/Y sky130_fd_sc_hd__inv_2
X_17199_ _17169_/X _17178_/X _17188_/X _17198_/X VGND VGND VPWR VPWR _17228_/A sky130_fd_sc_hd__or4_4
XANTENNA__14912__B2 _14911_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16114__B1 _15946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14711__A _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19909_ _19909_/A VGND VGND VPWR VPWR _19909_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12687__C1 _12641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24568__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22920_ _22915_/X _22918_/X _22919_/X VGND VGND VPWR VPWR _22920_/X sky130_fd_sc_hd__or3_4
XANTENNA__15245__C _15261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22851_ _16120_/Y _22523_/B _15855_/B _11720_/Y _21051_/A VGND VGND VPWR VPWR _22851_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_244_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21802_ _21665_/A _19929_/Y VGND VGND VPWR VPWR _21803_/C sky130_fd_sc_hd__or2_4
XFILLER_37_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24150__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22782_ _12428_/C _22499_/X _24274_/Q _21056_/X VGND VGND VPWR VPWR _22782_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21174__B1 _16365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24521_ _24520_/CLK _24521_/D HRESETn VGND VGND VPWR VPWR _16605_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21733_ _21569_/X _21731_/X _21575_/X _21732_/X VGND VGND VPWR VPWR _21733_/X sky130_fd_sc_hd__o22a_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24452_ _24463_/CLK _24452_/D HRESETn VGND VGND VPWR VPWR _24452_/Q sky130_fd_sc_hd__dfrtp_4
X_21664_ _21473_/A _19952_/Y VGND VGND VPWR VPWR _21666_/B sky130_fd_sc_hd__or2_4
XFILLER_197_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25132__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23403_ _23675_/CLK _23403_/D VGND VGND VPWR VPWR _23403_/Q sky130_fd_sc_hd__dfxtp_4
X_20615_ _20615_/A VGND VGND VPWR VPWR _20615_/X sky130_fd_sc_hd__buf_2
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25356__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24383_ _24725_/CLK _17136_/X HRESETn VGND VGND VPWR VPWR _24383_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22674__B1 _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21595_ _21748_/A _21594_/X VGND VGND VPWR VPWR _21595_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__16373__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25195__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23334_ _24477_/Q _22661_/X _23178_/X VGND VGND VPWR VPWR _23334_/X sky130_fd_sc_hd__o21a_4
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20546_ _20546_/A VGND VGND VPWR VPWR _23937_/D sky130_fd_sc_hd__inv_2
XFILLER_192_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_243_0_HCLK clkbuf_8_243_0_HCLK/A VGND VGND VPWR VPWR _24080_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_193_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22426__B1 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23265_ _23091_/A _23265_/B _23264_/X VGND VGND VPWR VPWR _23265_/X sky130_fd_sc_hd__and3_4
X_20477_ _13873_/X _20515_/B _20477_/C VGND VGND VPWR VPWR _20477_/X sky130_fd_sc_hd__or3_4
XFILLER_192_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25004_ _25204_/CLK _25004_/D HRESETn VGND VGND VPWR VPWR _15288_/A sky130_fd_sc_hd__dfrtp_4
X_22216_ _22226_/A _22214_/X _22215_/X VGND VGND VPWR VPWR _22220_/B sky130_fd_sc_hd__and3_4
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16105__B1 _15939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23196_ _23160_/A _23186_/X _23196_/C _23195_/X VGND VGND VPWR VPWR _23196_/X sky130_fd_sc_hd__or4_4
XFILLER_105_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22147_ _15704_/A _22145_/X _22146_/X VGND VGND VPWR VPWR _22147_/X sky130_fd_sc_hd__and3_4
XFILLER_133_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15717__A _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24991__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22078_ _21622_/A VGND VGND VPWR VPWR _22378_/A sky130_fd_sc_hd__buf_2
XANTENNA__24920__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13920_ _13920_/A VGND VGND VPWR VPWR _13953_/A sky130_fd_sc_hd__inv_2
X_21029_ _22641_/B VGND VGND VPWR VPWR _21030_/A sky130_fd_sc_hd__buf_2
XANTENNA__24238__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13851_ _20476_/B VGND VGND VPWR VPWR _13851_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21454__A _17709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19358__B1 _19357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12802_ _12801_/X _24800_/Q _12801_/X _24800_/Q VGND VGND VPWR VPWR _12802_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_216_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13782_ _21379_/B VGND VGND VPWR VPWR _13783_/D sky130_fd_sc_hd__buf_2
X_16570_ _16569_/Y _16567_/X _16395_/X _16567_/X VGND VGND VPWR VPWR _24535_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12733_ _12732_/Y _24816_/Q _12732_/Y _24816_/Q VGND VGND VPWR VPWR _12733_/X sky130_fd_sc_hd__a2bb2o_4
X_15521_ _11674_/A VGND VGND VPWR VPWR _15640_/A sky130_fd_sc_hd__inv_2
X_24719_ _24737_/CLK _24719_/D HRESETn VGND VGND VPWR VPWR _24719_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15919__B1 _24781_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18763__A _24143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15452_ _13907_/B _15451_/X _15426_/X _13903_/A _15447_/X VGND VGND VPWR VPWR _24962_/D
+ sky130_fd_sc_hd__a32o_4
X_18240_ _18240_/A VGND VGND VPWR VPWR _18240_/X sky130_fd_sc_hd__buf_2
X_12664_ _12664_/A _12671_/A _12664_/C _12663_/X VGND VGND VPWR VPWR _12670_/B sky130_fd_sc_hd__or4_4
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14403_/A VGND VGND VPWR VPWR _14403_/X sky130_fd_sc_hd__buf_2
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_53_0_HCLK clkbuf_5_26_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_53_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15383_ _15296_/A _15296_/B _15409_/A _15382_/X VGND VGND VPWR VPWR _15383_/X sky130_fd_sc_hd__or4_4
X_18171_ _17987_/X _18171_/B VGND VGND VPWR VPWR _18171_/X sky130_fd_sc_hd__or2_4
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17379__A _17203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12595_ _12505_/Y _12644_/A VGND VGND VPWR VPWR _12595_/X sky130_fd_sc_hd__or2_4
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20517__B _20517_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ _14334_/A _14345_/A VGND VGND VPWR VPWR _14339_/B sky130_fd_sc_hd__or2_4
X_17122_ _17043_/B _17117_/B _17118_/Y _17053_/X VGND VGND VPWR VPWR _17123_/A sky130_fd_sc_hd__a211o_4
XFILLER_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25026__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17053_ _17381_/B VGND VGND VPWR VPWR _17053_/X sky130_fd_sc_hd__buf_2
XFILLER_128_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14265_ _14264_/Y _14259_/X _13798_/X _14247_/A VGND VGND VPWR VPWR _14265_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16004_ HWDATA[27] VGND VGND VPWR VPWR _16004_/X sky130_fd_sc_hd__buf_2
X_13216_ _13369_/A _13209_/X _13215_/X VGND VGND VPWR VPWR _13217_/C sky130_fd_sc_hd__or3_4
XANTENNA__21629__A _22225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14196_ _20489_/B VGND VGND VPWR VPWR _20517_/B sky130_fd_sc_hd__inv_2
XANTENNA__23090__B1 _22098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13147_ _13168_/A _13147_/B VGND VGND VPWR VPWR _13147_/X sky130_fd_sc_hd__or2_4
XFILLER_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13078_ _12981_/D _13074_/X VGND VGND VPWR VPWR _13078_/Y sky130_fd_sc_hd__nand2_4
X_17955_ _17940_/A _17955_/B VGND VGND VPWR VPWR _17955_/X sky130_fd_sc_hd__or2_4
XANTENNA__24661__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12029_ _12029_/A VGND VGND VPWR VPWR _12029_/Y sky130_fd_sc_hd__inv_2
X_16906_ _16906_/A VGND VGND VPWR VPWR _16906_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13147__A _13168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17886_ _17880_/A _17850_/X VGND VGND VPWR VPWR _17886_/Y sky130_fd_sc_hd__nand2_4
XFILLER_239_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19625_ _19716_/C _20220_/B _19273_/A _20220_/D VGND VGND VPWR VPWR _19626_/A sky130_fd_sc_hd__or4_4
XANTENNA__21364__A _23964_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16837_ _16841_/A VGND VGND VPWR VPWR _16837_/X sky130_fd_sc_hd__buf_2
XFILLER_93_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19349__B1 _19282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16458__A _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19556_ _22029_/B _19550_/X _11911_/X _19555_/X VGND VGND VPWR VPWR _23696_/D sky130_fd_sc_hd__a2bb2o_4
X_16768_ _15018_/Y _16766_/X _16420_/X _16766_/X VGND VGND VPWR VPWR _24456_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18507_ _18499_/B _18498_/X _18499_/A VGND VGND VPWR VPWR _18507_/X sky130_fd_sc_hd__o21a_4
X_15719_ HWDATA[26] VGND VGND VPWR VPWR _15719_/X sky130_fd_sc_hd__buf_2
XANTENNA__19769__A _19764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19487_ _19494_/A VGND VGND VPWR VPWR _19487_/X sky130_fd_sc_hd__buf_2
XFILLER_202_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16699_ _24486_/Q VGND VGND VPWR VPWR _16699_/Y sky130_fd_sc_hd__inv_2
X_18438_ _18438_/A _18438_/B _18438_/C _18437_/X VGND VGND VPWR VPWR _18438_/X sky130_fd_sc_hd__or4_4
XANTENNA__16583__B1 _16226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20708__A _20708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24119__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17289__A _17234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18369_ _18354_/A VGND VGND VPWR VPWR _18369_/Y sky130_fd_sc_hd__inv_2
X_20400_ _23387_/Q VGND VGND VPWR VPWR _20400_/Y sky130_fd_sc_hd__inv_2
X_21380_ _21278_/X _21376_/X _21378_/Y _21379_/X VGND VGND VPWR VPWR _21380_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16335__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14425__B _14425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20331_ _20331_/A VGND VGND VPWR VPWR _22251_/B sky130_fd_sc_hd__inv_2
XFILLER_134_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16886__B2 _14777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23050_ _21427_/A VGND VGND VPWR VPWR _23050_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_10_0_HCLK clkbuf_7_5_0_HCLK/X VGND VGND VPWR VPWR _23808_/CLK sky130_fd_sc_hd__clkbuf_1
X_20262_ _20261_/X VGND VGND VPWR VPWR _20262_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21539__A _21087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24560__D _16504_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24749__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22001_ _21960_/B VGND VGND VPWR VPWR _22001_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_73_0_HCLK clkbuf_7_36_0_HCLK/X VGND VGND VPWR VPWR _24744_/CLK sky130_fd_sc_hd__clkbuf_1
X_20193_ _21611_/B _20192_/X _20106_/X _20192_/X VGND VGND VPWR VPWR _20193_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14441__A _14096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19588__B1 _19587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23952_ _23951_/CLK _23952_/D HRESETn VGND VGND VPWR VPWR _23952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_243_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24331__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13872__A1 _23995_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22903_ _23043_/A _22903_/B VGND VGND VPWR VPWR _22913_/C sky130_fd_sc_hd__and2_4
XANTENNA__21274__A _21177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18260__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23883_ _23875_/CLK _23883_/D VGND VGND VPWR VPWR _19022_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_45_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16368__A _16368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22834_ _23129_/A _22830_/X _22831_/X _22833_/X VGND VGND VPWR VPWR _22835_/A sky130_fd_sc_hd__o22a_4
XFILLER_244_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22765_ _22764_/X VGND VGND VPWR VPWR _22766_/D sky130_fd_sc_hd__inv_2
XFILLER_197_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25537__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24504_ _24060_/CLK _16656_/X HRESETn VGND VGND VPWR VPWR _24504_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22817__B _22817_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19760__B1 _19759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21716_ _25105_/Q _22119_/B VGND VGND VPWR VPWR _21716_/Y sky130_fd_sc_hd__nand2_4
X_25484_ _23938_/CLK _12066_/X HRESETn VGND VGND VPWR VPWR _25484_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21721__B _21721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22696_ _22696_/A _22696_/B VGND VGND VPWR VPWR _22696_/Y sky130_fd_sc_hd__nor2_4
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24435_ _24462_/CLK _24435_/D HRESETn VGND VGND VPWR VPWR _24435_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_184_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21647_ _21643_/X _21646_/X _25273_/Q _18263_/X VGND VGND VPWR VPWR _21647_/X sky130_fd_sc_hd__o22a_4
XFILLER_200_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12380_ _12204_/Y _12264_/Y _12379_/X VGND VGND VPWR VPWR _12380_/X sky130_fd_sc_hd__or3_4
X_24366_ _24365_/CLK _24366_/D HRESETn VGND VGND VPWR VPWR _17292_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16326__B1 _16229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21578_ _21556_/Y _21564_/X _21567_/X _21577_/Y VGND VGND VPWR VPWR _21601_/B sky130_fd_sc_hd__a211o_4
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23317_ _22552_/X _23316_/X _22135_/C _24114_/Q _22555_/X VGND VGND VPWR VPWR _23317_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_126_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20529_ _20529_/A _20528_/X VGND VGND VPWR VPWR _20535_/B sky130_fd_sc_hd__or2_4
X_24297_ _24297_/CLK _17685_/X HRESETn VGND VGND VPWR VPWR _24297_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14050_ _13995_/A _14046_/X _14049_/X VGND VGND VPWR VPWR _14050_/Y sky130_fd_sc_hd__o21ai_4
X_23248_ _23248_/A _22890_/B VGND VGND VPWR VPWR _23251_/B sky130_fd_sc_hd__or2_4
XFILLER_134_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13001_ _13001_/A VGND VGND VPWR VPWR _13001_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23179_ _15046_/A _23002_/X _23178_/X VGND VGND VPWR VPWR _23179_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24419__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15166__B _15242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19579__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18758__A _18692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17740_ _16950_/X VGND VGND VPWR VPWR _17810_/A sky130_fd_sc_hd__buf_2
XFILLER_153_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14952_ _15065_/A _16810_/A _14951_/A _16810_/A VGND VGND VPWR VPWR _14952_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24072__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13903_ _13903_/A _13903_/B _13917_/B _13880_/X VGND VGND VPWR VPWR _14231_/A sky130_fd_sc_hd__or4_4
XFILLER_248_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17671_ _17519_/Y _17670_/X VGND VGND VPWR VPWR _17671_/X sky130_fd_sc_hd__or2_4
XFILLER_235_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17381__B _17381_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24001__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14883_ _14883_/A VGND VGND VPWR VPWR _14883_/Y sky130_fd_sc_hd__inv_2
X_19410_ _17956_/B VGND VGND VPWR VPWR _19410_/Y sky130_fd_sc_hd__inv_2
X_16622_ _16621_/X VGND VGND VPWR VPWR _16622_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13834_ _13552_/Y _13832_/X _13791_/X _13832_/X VGND VGND VPWR VPWR _13834_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19341_ _19341_/A _13596_/A _19163_/C VGND VGND VPWR VPWR _19342_/A sky130_fd_sc_hd__or3_4
XFILLER_216_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13765_ _13765_/A VGND VGND VPWR VPWR _14395_/A sky130_fd_sc_hd__buf_2
X_16553_ _16552_/Y _16548_/X _16467_/X _16548_/X VGND VGND VPWR VPWR _16553_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17010__A1_N _15993_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15504_ _15503_/Y _15499_/X HADDR[15] _15499_/X VGND VGND VPWR VPWR _15504_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12716_ _12716_/A _12716_/B VGND VGND VPWR VPWR _12721_/B sky130_fd_sc_hd__or2_4
X_19272_ _23794_/Q VGND VGND VPWR VPWR _19272_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13696_ _13679_/A _13694_/X _13695_/Y _13690_/X _11804_/A VGND VGND VPWR VPWR _25292_/D
+ sky130_fd_sc_hd__a32o_4
X_16484_ _16481_/Y _16482_/X _16483_/X _16482_/X VGND VGND VPWR VPWR _24568_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16565__B1 _16391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18223_ _18094_/A _18223_/B _18222_/X VGND VGND VPWR VPWR _18227_/B sky130_fd_sc_hd__and3_4
X_12647_ _12560_/A _12650_/B VGND VGND VPWR VPWR _12648_/C sky130_fd_sc_hd__or2_4
X_15435_ _13927_/B _15432_/X _15427_/X _13913_/X _15433_/X VGND VGND VPWR VPWR _15435_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15366_ _15366_/A _15370_/B VGND VGND VPWR VPWR _15366_/Y sky130_fd_sc_hd__nand2_4
X_18154_ _18014_/A _18154_/B VGND VGND VPWR VPWR _18155_/C sky130_fd_sc_hd__or2_4
X_12578_ _12578_/A VGND VGND VPWR VPWR _12578_/Y sky130_fd_sc_hd__inv_2
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17105_ _17105_/A _17099_/X _17104_/Y VGND VGND VPWR VPWR _24391_/D sky130_fd_sc_hd__and3_4
X_14317_ _25169_/Q _12151_/X _14316_/Y VGND VGND VPWR VPWR _25169_/D sky130_fd_sc_hd__o21a_4
X_15297_ _15417_/A VGND VGND VPWR VPWR _15409_/A sky130_fd_sc_hd__inv_2
X_18085_ _18085_/A _18083_/X _18085_/C VGND VGND VPWR VPWR _18085_/X sky130_fd_sc_hd__and3_4
XFILLER_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14248_ _14242_/Y _14247_/X _13824_/X _14247_/X VGND VGND VPWR VPWR _14248_/X sky130_fd_sc_hd__a2bb2o_4
X_17036_ _17036_/A VGND VGND VPWR VPWR _17125_/A sky130_fd_sc_hd__inv_2
XANTENNA__24842__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14179_ _16366_/A _14179_/B VGND VGND VPWR VPWR _14184_/A sky130_fd_sc_hd__or2_4
XFILLER_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21078__B _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18987_ _18983_/Y _18977_/X _18985_/X _18986_/X VGND VGND VPWR VPWR _23896_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17938_ _17942_/A _17938_/B _17938_/C VGND VGND VPWR VPWR _17938_/X sky130_fd_sc_hd__and3_4
XFILLER_100_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17869_ _16925_/Y _17853_/D VGND VGND VPWR VPWR _17873_/B sky130_fd_sc_hd__or2_4
XFILLER_66_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19608_ _19605_/Y _19599_/X _19606_/X _19607_/X VGND VGND VPWR VPWR _19608_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20880_ _13649_/X VGND VGND VPWR VPWR _20880_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21129__B1 _21127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19539_ _19526_/A VGND VGND VPWR VPWR _19539_/X sky130_fd_sc_hd__buf_2
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22550_ _24525_/Q _21098_/X _21738_/X _22549_/X VGND VGND VPWR VPWR _22550_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16556__B1 _16382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18860__A2_N _18613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21501_ _22393_/A VGND VGND VPWR VPWR _21501_/X sky130_fd_sc_hd__buf_2
XFILLER_195_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22481_ _22638_/B VGND VGND VPWR VPWR _22901_/B sky130_fd_sc_hd__buf_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24220_ _24233_/CLK _24220_/D HRESETn VGND VGND VPWR VPWR _13682_/A sky130_fd_sc_hd__dfrtp_4
X_21432_ _21431_/X VGND VGND VPWR VPWR _21525_/A sky130_fd_sc_hd__buf_2
XFILLER_148_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24151_ _24146_/CLK _24151_/D HRESETn VGND VGND VPWR VPWR _24151_/Q sky130_fd_sc_hd__dfrtp_4
X_21363_ _14179_/B _21343_/B VGND VGND VPWR VPWR _21556_/A sky130_fd_sc_hd__or2_4
XFILLER_190_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23102_ _23035_/X _23101_/X _22858_/X _24845_/Q _23037_/X VGND VGND VPWR VPWR _23102_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20314_ _21984_/D VGND VGND VPWR VPWR _21974_/A sky130_fd_sc_hd__inv_2
XFILLER_163_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24082_ _23926_/CLK _24082_/D HRESETn VGND VGND VPWR VPWR _20437_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__23054__B1 _17744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21294_ _21864_/B VGND VGND VPWR VPWR _21294_/X sky130_fd_sc_hd__buf_2
XFILLER_190_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24583__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23033_ _23028_/Y _23032_/Y _22854_/X VGND VGND VPWR VPWR _23033_/X sky130_fd_sc_hd__o21a_4
X_20245_ _20245_/A VGND VGND VPWR VPWR _22198_/B sky130_fd_sc_hd__inv_2
XANTENNA__24512__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21419__D _21418_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20176_ _21263_/B _20171_/X _20133_/X _20158_/Y VGND VGND VPWR VPWR _23475_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21716__B _22119_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24984_ _24985_/CLK _15398_/X HRESETn VGND VGND VPWR VPWR _15093_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_85_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23935_ _23932_/CLK _20987_/B HRESETn VGND VGND VPWR VPWR _23935_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__22580__A2 _21031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11880_ _11853_/X _11850_/Y _11869_/A _25515_/Q VGND VGND VPWR VPWR _11881_/A sky130_fd_sc_hd__a211o_4
X_23866_ _23610_/CLK _23866_/D VGND VGND VPWR VPWR _23866_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16795__B1 _15545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22817_ _16492_/A _22817_/B _22817_/C VGND VGND VPWR VPWR _22817_/X sky130_fd_sc_hd__and3_4
XANTENNA__25371__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23797_ _23806_/CLK _23797_/D VGND VGND VPWR VPWR _23797_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16826__A _24428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22332__A2 _21349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13550_ _22695_/A _25097_/Q _22695_/A _25097_/Q VGND VGND VPWR VPWR _13550_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22748_ _24763_/Q _22487_/X VGND VGND VPWR VPWR _22748_/X sky130_fd_sc_hd__or2_4
X_25536_ _25538_/CLK _25536_/D HRESETn VGND VGND VPWR VPWR _25536_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_197_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12501_ _12500_/Y _24886_/Q _12500_/Y _24886_/Q VGND VGND VPWR VPWR _12501_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_198_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13481_ _13480_/Y _13476_/X _13459_/X _13464_/A VGND VGND VPWR VPWR _25317_/D sky130_fd_sc_hd__a2bb2o_4
X_25467_ _25109_/CLK _12158_/X HRESETn VGND VGND VPWR VPWR SCLK_S3 sky130_fd_sc_hd__dfstp_4
X_22679_ _20744_/Y _22992_/A _20883_/Y _21597_/X VGND VGND VPWR VPWR _22679_/X sky130_fd_sc_hd__o22a_4
X_15220_ _15203_/X _15214_/X _15219_/Y VGND VGND VPWR VPWR _25026_/D sky130_fd_sc_hd__and3_4
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12432_ _12428_/B _12431_/X VGND VGND VPWR VPWR _12433_/B sky130_fd_sc_hd__or2_4
X_24418_ _24419_/CLK _24418_/D HRESETn VGND VGND VPWR VPWR _24418_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25398_ _25397_/CLK _25398_/D HRESETn VGND VGND VPWR VPWR _12818_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15151_ _15150_/Y _24610_/Q _15150_/Y _24610_/Q VGND VGND VPWR VPWR _15156_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12363_ _12990_/A _24850_/Q _12990_/A _24850_/Q VGND VGND VPWR VPWR _12363_/X sky130_fd_sc_hd__a2bb2o_4
X_24349_ _24667_/CLK _24349_/D HRESETn VGND VGND VPWR VPWR _24349_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14102_ _23956_/Q _14087_/X _14102_/C VGND VGND VPWR VPWR _14102_/X sky130_fd_sc_hd__or3_4
XFILLER_165_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15082_ _15082_/A VGND VGND VPWR VPWR _15082_/Y sky130_fd_sc_hd__inv_2
X_12294_ _25361_/Q VGND VGND VPWR VPWR _13005_/A sky130_fd_sc_hd__inv_2
XANTENNA__15522__B2 _15519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14033_ _14008_/A _14007_/D _13967_/Y _14007_/B VGND VGND VPWR VPWR _14033_/X sky130_fd_sc_hd__or4_4
X_18910_ _18910_/A _18910_/B _18326_/C VGND VGND VPWR VPWR _19047_/C sky130_fd_sc_hd__or3_4
XANTENNA__12336__B2 _24832_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19890_ _19890_/A VGND VGND VPWR VPWR _21676_/B sky130_fd_sc_hd__inv_2
XFILLER_107_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24253__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18841_ _16512_/A _24135_/Q _16512_/Y _18789_/A VGND VGND VPWR VPWR _18841_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18772_ _18691_/B _18767_/B _18735_/X _18768_/Y VGND VGND VPWR VPWR _18773_/A sky130_fd_sc_hd__a211o_4
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15984_ _15984_/A _14365_/B _14365_/C _15984_/D VGND VGND VPWR VPWR _15985_/B sky130_fd_sc_hd__or4_4
XFILLER_94_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17723_ _17723_/A VGND VGND VPWR VPWR _22257_/A sky130_fd_sc_hd__buf_2
X_14935_ _14935_/A _14905_/X _14935_/C _14935_/D VGND VGND VPWR VPWR _14935_/X sky130_fd_sc_hd__or4_4
XANTENNA__25459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17654_ _17653_/X VGND VGND VPWR VPWR _24305_/D sky130_fd_sc_hd__inv_2
XFILLER_180_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14866_ _14865_/X VGND VGND VPWR VPWR _14866_/X sky130_fd_sc_hd__buf_2
XFILLER_36_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16605_ _16605_/A VGND VGND VPWR VPWR _16605_/Y sky130_fd_sc_hd__inv_2
X_13817_ _13810_/A VGND VGND VPWR VPWR _13817_/X sky130_fd_sc_hd__buf_2
X_17585_ _17585_/A _17584_/X VGND VGND VPWR VPWR _17585_/X sky130_fd_sc_hd__or2_4
XFILLER_16_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14797_ _25051_/Q _14796_/X _25052_/Q VGND VGND VPWR VPWR _14797_/X sky130_fd_sc_hd__or3_4
XFILLER_189_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19324_ _23777_/Q VGND VGND VPWR VPWR _19324_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16536_ _24547_/Q VGND VGND VPWR VPWR _16536_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25041__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13748_ _13744_/X _13745_/X _13747_/Y VGND VGND VPWR VPWR _13748_/Y sky130_fd_sc_hd__a21oi_4
X_19255_ _19251_/Y _19254_/X _16860_/X _19254_/X VGND VGND VPWR VPWR _23802_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16467_ HWDATA[27] VGND VGND VPWR VPWR _16467_/X sky130_fd_sc_hd__buf_2
X_13679_ _13679_/A VGND VGND VPWR VPWR _13692_/B sky130_fd_sc_hd__inv_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18951__A _18951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18206_ _18027_/A _23747_/Q VGND VGND VPWR VPWR _18208_/B sky130_fd_sc_hd__or2_4
X_15418_ _15418_/A _15418_/B _15402_/X VGND VGND VPWR VPWR _15418_/X sky130_fd_sc_hd__and3_4
X_19186_ _19191_/A VGND VGND VPWR VPWR _19186_/X sky130_fd_sc_hd__buf_2
Xclkbuf_5_23_0_HCLK clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_46_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16398_ _16387_/A VGND VGND VPWR VPWR _16398_/X sky130_fd_sc_hd__buf_2
XFILLER_129_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18137_ _18030_/A _18137_/B _18137_/C VGND VGND VPWR VPWR _18141_/B sky130_fd_sc_hd__and3_4
X_15349_ _15349_/A VGND VGND VPWR VPWR _15349_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21834__B2 _21833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18068_ _18030_/A _18068_/B _18067_/X VGND VGND VPWR VPWR _18072_/B sky130_fd_sc_hd__and3_4
XFILLER_208_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12300__A2_N _24820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16710__B1 _16353_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13524__B1 _13459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17019_ _24403_/Q VGND VGND VPWR VPWR _17019_/Y sky130_fd_sc_hd__inv_2
X_20030_ _21201_/B _20025_/X _20008_/X _20012_/Y VGND VGND VPWR VPWR _20030_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18906__A1_N _17517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_147_0_HCLK clkbuf_7_73_0_HCLK/X VGND VGND VPWR VPWR _25492_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__23976__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21981_ _21978_/X _21979_/X _21980_/X VGND VGND VPWR VPWR _21981_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_227_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23720_ _23406_/CLK _23720_/D VGND VGND VPWR VPWR _23720_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20932_ _24059_/Q _20932_/B VGND VGND VPWR VPWR _20932_/Y sky130_fd_sc_hd__nor2_4
XFILLER_39_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25129__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23651_ _24209_/CLK _23651_/D VGND VGND VPWR VPWR _13436_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ _24043_/Q _20857_/X _20862_/X VGND VGND VPWR VPWR _20863_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_241_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22314__A2 _14182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22602_ _22602_/A _21101_/A VGND VGND VPWR VPWR _22602_/X sky130_fd_sc_hd__or2_4
XFILLER_230_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23582_ _23555_/CLK _19889_/X VGND VGND VPWR VPWR _19888_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16529__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20794_ _20793_/A _20793_/B _20793_/Y VGND VGND VPWR VPWR _20794_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25321_ _25158_/CLK _25321_/D HRESETn VGND VGND VPWR VPWR _25321_/Q sky130_fd_sc_hd__dfrtp_4
X_22533_ _21737_/X VGND VGND VPWR VPWR _22533_/X sky130_fd_sc_hd__buf_2
XFILLER_179_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25252_ _25230_/CLK _13854_/X HRESETn VGND VGND VPWR VPWR _20476_/B sky130_fd_sc_hd__dfrtp_4
X_22464_ _22463_/X VGND VGND VPWR VPWR _22472_/B sky130_fd_sc_hd__inv_2
XANTENNA__24764__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24203_ _23456_/CLK _18349_/Y HRESETn VGND VGND VPWR VPWR _13189_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_148_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21415_ _25064_/Q _21407_/X _21414_/X VGND VGND VPWR VPWR _21415_/X sky130_fd_sc_hd__or3_4
XFILLER_136_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25183_ _25308_/CLK _25183_/D HRESETn VGND VGND VPWR VPWR _13509_/A sky130_fd_sc_hd__dfrtp_4
X_22395_ _22395_/A VGND VGND VPWR VPWR _22395_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24134_ _24148_/CLK _18803_/Y HRESETn VGND VGND VPWR VPWR _24134_/Q sky130_fd_sc_hd__dfrtp_4
X_21346_ _21346_/A VGND VGND VPWR VPWR _22181_/B sky130_fd_sc_hd__buf_2
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23027__B1 _12356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24065_ _24060_/CLK _20959_/X HRESETn VGND VGND VPWR VPWR _24065_/Q sky130_fd_sc_hd__dfrtp_4
X_21277_ _19594_/A _20307_/X _23699_/Q _21215_/X VGND VGND VPWR VPWR _21277_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23016_ _12804_/Y _21879_/X _16940_/Y _22826_/X VGND VGND VPWR VPWR _23016_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20228_ _20226_/Y _20222_/X _19746_/X _20227_/X VGND VGND VPWR VPWR _20228_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_43_0_HCLK clkbuf_7_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_87_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15725__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20159_ _20158_/Y VGND VGND VPWR VPWR _20159_/X sky130_fd_sc_hd__buf_2
X_12981_ _13097_/A _12321_/Y _12981_/C _12981_/D VGND VGND VPWR VPWR _12981_/X sky130_fd_sc_hd__or4_4
XFILLER_92_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24967_ _24967_/CLK _15445_/X HRESETn VGND VGND VPWR VPWR _13932_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_217_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18757__A1 _18693_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19954__B1 _19617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14720_ _14720_/A VGND VGND VPWR VPWR _14720_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13245__A _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11932_ _11967_/A _11932_/B _11932_/C VGND VGND VPWR VPWR _11932_/X sky130_fd_sc_hd__and3_4
X_23918_ _23912_/CLK _18923_/X VGND VGND VPWR VPWR _13334_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_245_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16768__B1 _16420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20564__A1 _14428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24898_ _24900_/CLK _15624_/X HRESETn VGND VGND VPWR VPWR _24898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_72_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22558__A _22558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11863_ _11796_/B VGND VGND VPWR VPWR _11863_/Y sky130_fd_sc_hd__inv_2
X_14651_ _13615_/A VGND VGND VPWR VPWR _19320_/A sky130_fd_sc_hd__buf_2
X_23849_ _23831_/CLK _19123_/X VGND VGND VPWR VPWR _18012_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _18026_/A VGND VGND VPWR VPWR _18095_/A sky130_fd_sc_hd__buf_2
XPHY_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _17351_/A _17366_/B _17370_/C VGND VGND VPWR VPWR _17370_/X sky130_fd_sc_hd__and3_4
XPHY_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _11682_/Y VGND VGND VPWR VPWR _11794_/X sky130_fd_sc_hd__buf_2
X_14582_ _14557_/X _14575_/X _14581_/Y _14579_/X _13566_/A VGND VGND VPWR VPWR _25092_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16321_ _16317_/Y _16319_/X _16320_/X _16319_/X VGND VGND VPWR VPWR _24628_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ _25267_/Q VGND VGND VPWR VPWR _13533_/Y sky130_fd_sc_hd__inv_2
X_25519_ _25499_/CLK _11862_/X HRESETn VGND VGND VPWR VPWR _25519_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19040_ _19028_/A VGND VGND VPWR VPWR _19040_/X sky130_fd_sc_hd__buf_2
X_13464_ _13464_/A VGND VGND VPWR VPWR _13464_/X sky130_fd_sc_hd__buf_2
X_16252_ _16239_/A VGND VGND VPWR VPWR _16252_/X sky130_fd_sc_hd__buf_2
XANTENNA__23266__B1 _23261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22293__A _21748_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12415_ _12415_/A _12412_/B _12414_/X VGND VGND VPWR VPWR _12416_/A sky130_fd_sc_hd__or3_4
X_15203_ _15241_/A VGND VGND VPWR VPWR _15203_/X sky130_fd_sc_hd__buf_2
XFILLER_173_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13395_ _13285_/A _13395_/B VGND VGND VPWR VPWR _13395_/X sky130_fd_sc_hd__or2_4
X_16183_ _16368_/A _16540_/B VGND VGND VPWR VPWR _16183_/Y sky130_fd_sc_hd__nor2_4
XFILLER_154_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24434__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12346_ _25350_/Q VGND VGND VPWR VPWR _12976_/C sky130_fd_sc_hd__inv_2
X_15134_ _15369_/A VGND VGND VPWR VPWR _15356_/A sky130_fd_sc_hd__inv_2
X_15065_ _15065_/A _14995_/X _15055_/X _15064_/X VGND VGND VPWR VPWR _15065_/X sky130_fd_sc_hd__or4_4
X_19942_ _22346_/B _19941_/X _19600_/X _19941_/X VGND VGND VPWR VPWR _19942_/X sky130_fd_sc_hd__a2bb2o_4
X_12277_ _12232_/Y _12240_/Y _12265_/X _12402_/B VGND VGND VPWR VPWR _12277_/X sky130_fd_sc_hd__or4_4
XFILLER_99_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14016_ _13984_/B _14010_/X _14536_/B VGND VGND VPWR VPWR _14059_/A sky130_fd_sc_hd__a21o_4
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19873_ _23587_/Q VGND VGND VPWR VPWR _21200_/B sky130_fd_sc_hd__inv_2
XANTENNA__15259__B1 _15185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18824_ _18744_/A _18815_/B _18824_/C VGND VGND VPWR VPWR _18824_/X sky130_fd_sc_hd__and3_4
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22529__C1 _22528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18755_ _18760_/A _18755_/B _18692_/Y _18746_/X VGND VGND VPWR VPWR _18755_/X sky130_fd_sc_hd__or4_4
XANTENNA__25293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_0_0_HCLK clkbuf_5_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_15967_ _12209_/Y _15964_/X _15752_/X _15964_/X VGND VGND VPWR VPWR _15967_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14482__B2 _14468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22544__A2 _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17706_ _17706_/A VGND VGND VPWR VPWR _17706_/X sky130_fd_sc_hd__buf_2
XFILLER_208_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14918_ _25015_/Q _14917_/A _15059_/A _14917_/Y VGND VGND VPWR VPWR _14919_/D sky130_fd_sc_hd__o22a_4
XANTENNA__25222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18686_ _18686_/A _18686_/B _18682_/X _18686_/D VGND VGND VPWR VPWR _18745_/D sky130_fd_sc_hd__or4_4
XFILLER_64_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15898_ _15701_/X _15887_/X _15830_/X _24789_/Q _15857_/A VGND VGND VPWR VPWR _24789_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22468__A _22468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17637_ _17569_/D _17637_/B VGND VGND VPWR VPWR _17638_/B sky130_fd_sc_hd__or2_4
X_14849_ _14840_/X _14848_/Y _24958_/Q _14840_/X VGND VGND VPWR VPWR _14849_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23290__C _22140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17568_ _17568_/A VGND VGND VPWR VPWR _17569_/D sky130_fd_sc_hd__inv_2
XFILLER_51_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22847__A3 _16724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19307_ _19305_/Y _19300_/X _19282_/X _19306_/X VGND VGND VPWR VPWR _23784_/D sky130_fd_sc_hd__a2bb2o_4
X_16519_ _16517_/Y _16513_/X _16518_/X _16513_/X VGND VGND VPWR VPWR _24554_/D sky130_fd_sc_hd__a2bb2o_4
X_17499_ _24301_/Q VGND VGND VPWR VPWR _17499_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19238_ _19232_/Y VGND VGND VPWR VPWR _19238_/X sky130_fd_sc_hd__buf_2
XFILLER_176_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19169_ _19169_/A VGND VGND VPWR VPWR _19169_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24175__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21200_ _21205_/A _21200_/B VGND VGND VPWR VPWR _21202_/B sky130_fd_sc_hd__or2_4
XFILLER_191_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22180_ _22179_/X VGND VGND VPWR VPWR _22180_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24104__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21131_ _21117_/Y _21119_/X _21122_/X _21130_/X VGND VGND VPWR VPWR _21131_/X sky130_fd_sc_hd__a211o_4
XFILLER_160_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22232__A1 _13538_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21062_ _22525_/A VGND VGND VPWR VPWR _21062_/X sky130_fd_sc_hd__buf_2
XANTENNA__21547__A _21545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18436__B1 _22996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20013_ _20012_/Y VGND VGND VPWR VPWR _20013_/X sky130_fd_sc_hd__buf_2
XANTENNA__15545__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16998__B1 _24737_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24821_ _24804_/CLK _15834_/X HRESETn VGND VGND VPWR VPWR _24821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17760__A _24274_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21964_ _21964_/A _19592_/Y VGND VGND VPWR VPWR _21964_/X sky130_fd_sc_hd__and2_4
X_24752_ _24800_/CLK _24752_/D HRESETn VGND VGND VPWR VPWR _24752_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_227_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20915_ _24055_/Q VGND VGND VPWR VPWR _20916_/A sky130_fd_sc_hd__inv_2
X_23703_ _24208_/CLK _23703_/D VGND VGND VPWR VPWR _23703_/Q sky130_fd_sc_hd__dfxtp_4
X_24683_ _24704_/CLK _24683_/D HRESETn VGND VGND VPWR VPWR _21521_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21895_ _21911_/A _21892_/X _21894_/X VGND VGND VPWR VPWR _21895_/X sky130_fd_sc_hd__and3_4
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15280__A _15311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23634_ _25326_/CLK _19741_/X VGND VGND VPWR VPWR _23634_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ _20846_/A VGND VGND VPWR VPWR _20846_/X sky130_fd_sc_hd__buf_2
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24945__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23565_ _24297_/CLK _23565_/D VGND VGND VPWR VPWR _19931_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20777_ _20776_/Y _20777_/B VGND VGND VPWR VPWR _20777_/X sky130_fd_sc_hd__and2_4
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22516_ _13820_/Y _22051_/X VGND VGND VPWR VPWR _22516_/X sky130_fd_sc_hd__and2_4
X_25304_ _25492_/CLK _25304_/D HRESETn VGND VGND VPWR VPWR _25304_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23496_ _23490_/CLK _23496_/D VGND VGND VPWR VPWR _23496_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23002__A _23002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22447_ _17352_/B _22430_/X _25441_/Q _22769_/A VGND VGND VPWR VPWR _22447_/X sky130_fd_sc_hd__a2bb2o_4
X_25235_ _25230_/CLK _25235_/D HRESETn VGND VGND VPWR VPWR _13979_/C sky130_fd_sc_hd__dfrtp_4
X_12200_ _12189_/X _12193_/X _12196_/X _12199_/X VGND VGND VPWR VPWR _12215_/C sky130_fd_sc_hd__or4_4
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13180_ _13176_/X _13179_/X _13162_/X VGND VGND VPWR VPWR _13180_/X sky130_fd_sc_hd__o21a_4
X_25166_ _25164_/CLK _14325_/X HRESETn VGND VGND VPWR VPWR _25166_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22378_ _22378_/A _20240_/Y VGND VGND VPWR VPWR _22378_/X sky130_fd_sc_hd__or2_4
XFILLER_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22841__A _21579_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12131_ _12131_/A VGND VGND VPWR VPWR _12131_/Y sky130_fd_sc_hd__inv_2
X_24117_ _24325_/CLK _18898_/X HRESETn VGND VGND VPWR VPWR _20994_/A sky130_fd_sc_hd__dfrtp_4
X_21329_ _21582_/A VGND VGND VPWR VPWR _21338_/A sky130_fd_sc_hd__inv_2
XFILLER_191_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25097_ _24188_/CLK _14567_/X HRESETn VGND VGND VPWR VPWR _25097_/Q sky130_fd_sc_hd__dfrtp_4
X_12062_ _25485_/Q VGND VGND VPWR VPWR _12062_/Y sky130_fd_sc_hd__inv_2
X_24048_ _24487_/CLK _24048_/D HRESETn VGND VGND VPWR VPWR _24048_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16870_ _16868_/Y _16865_/X _16869_/X _16865_/X VGND VGND VPWR VPWR _24410_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15821_ _12293_/Y _15820_/X _13818_/X _15820_/X VGND VGND VPWR VPWR _24830_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16695__A1_N _16694_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_130_0_HCLK clkbuf_7_65_0_HCLK/X VGND VGND VPWR VPWR _23627_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_46_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18540_ _18467_/A _18540_/B VGND VGND VPWR VPWR _18540_/Y sky130_fd_sc_hd__nand2_4
X_15752_ HWDATA[9] VGND VGND VPWR VPWR _15752_/X sky130_fd_sc_hd__buf_2
X_12964_ _12833_/C _12958_/B VGND VGND VPWR VPWR _12965_/C sky130_fd_sc_hd__nand2_4
XFILLER_234_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_193_0_HCLK clkbuf_7_96_0_HCLK/X VGND VGND VPWR VPWR _24678_/CLK sky130_fd_sc_hd__clkbuf_1
X_14703_ _21787_/A _14697_/X _14702_/X VGND VGND VPWR VPWR _14703_/Y sky130_fd_sc_hd__a21oi_4
X_11915_ _19610_/A VGND VGND VPWR VPWR _11915_/X sky130_fd_sc_hd__buf_2
X_18471_ _18567_/A _18409_/Y _18577_/A _18471_/D VGND VGND VPWR VPWR _18478_/A sky130_fd_sc_hd__or4_4
X_15683_ _15676_/Y _15686_/A _15686_/B VGND VGND VPWR VPWR _15683_/X sky130_fd_sc_hd__or3_4
XFILLER_205_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12895_ _12895_/A _12894_/Y VGND VGND VPWR VPWR _12897_/B sky130_fd_sc_hd__or2_4
XFILLER_233_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17422_ _17429_/A VGND VGND VPWR VPWR _17422_/X sky130_fd_sc_hd__buf_2
XFILLER_221_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14634_ _18026_/A VGND VGND VPWR VPWR _18090_/A sky130_fd_sc_hd__inv_2
X_11846_ _11837_/X _11846_/B _11842_/X _11846_/D VGND VGND VPWR VPWR _11846_/X sky130_fd_sc_hd__or4_4
XFILLER_233_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24686__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17347_/C _17352_/X _17284_/X _17349_/B VGND VGND VPWR VPWR _17354_/A sky130_fd_sc_hd__a211o_4
XFILLER_14_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _25523_/Q VGND VGND VPWR VPWR _11777_/Y sky130_fd_sc_hd__inv_2
X_14565_ _14543_/Y _14546_/X _14563_/X _25098_/Q _14564_/Y VGND VGND VPWR VPWR _14565_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_198_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24615__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16304_ _16303_/Y _16298_/X _15942_/X _16298_/X VGND VGND VPWR VPWR _24634_/D sky130_fd_sc_hd__a2bb2o_4
X_13516_ _13503_/Y _13515_/Y SCLK_S2 _13514_/X VGND VGND VPWR VPWR _13516_/X sky130_fd_sc_hd__o22a_4
XFILLER_158_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23239__B1 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17284_ _17284_/A VGND VGND VPWR VPWR _17284_/X sky130_fd_sc_hd__buf_2
X_14496_ _14494_/X _14495_/Y _14490_/B VGND VGND VPWR VPWR _14496_/X sky130_fd_sc_hd__a21o_4
XANTENNA_clkbuf_4_1_0_HCLK_A clkbuf_3_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19023_ _19022_/Y _19018_/X _18998_/X _19011_/A VGND VGND VPWR VPWR _23883_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16235_ _24659_/Q VGND VGND VPWR VPWR _16235_/Y sky130_fd_sc_hd__inv_2
X_13447_ _13314_/X _13447_/B _13446_/X VGND VGND VPWR VPWR _13448_/C sky130_fd_sc_hd__and3_4
XFILLER_9_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14973__A2_N _16796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13378_ _13220_/X _19706_/A VGND VGND VPWR VPWR _13378_/X sky130_fd_sc_hd__or2_4
X_16166_ _14765_/A _14756_/A VGND VGND VPWR VPWR _16166_/X sky130_fd_sc_hd__or2_4
XANTENNA__18666__B1 _16610_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15117_ _24597_/Q VGND VGND VPWR VPWR _15117_/Y sky130_fd_sc_hd__inv_2
X_12329_ _24837_/Q VGND VGND VPWR VPWR _12329_/Y sky130_fd_sc_hd__inv_2
X_16097_ _16096_/Y _16092_/X _16004_/X _16092_/X VGND VGND VPWR VPWR _24708_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15048_ _25034_/Q _15046_/Y _25028_/Q _15047_/Y VGND VGND VPWR VPWR _15048_/X sky130_fd_sc_hd__a2bb2o_4
X_19925_ _19932_/A VGND VGND VPWR VPWR _19925_/X sky130_fd_sc_hd__buf_2
XFILLER_114_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20225__B1 _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19856_ _19856_/A VGND VGND VPWR VPWR _19856_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25403__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18807_ _18686_/A _18809_/B _18806_/Y VGND VGND VPWR VPWR _24133_/D sky130_fd_sc_hd__o21a_4
X_19787_ _19786_/Y _19784_/X _19743_/X _19784_/X VGND VGND VPWR VPWR _19787_/X sky130_fd_sc_hd__a2bb2o_4
X_16999_ _16035_/Y _24388_/Q _16035_/Y _24388_/Q VGND VGND VPWR VPWR _17000_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18738_ _18729_/B VGND VGND VPWR VPWR _18738_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22629__C _22628_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18669_ _18647_/X _18669_/B _18669_/C _18668_/X VGND VGND VPWR VPWR _18670_/B sky130_fd_sc_hd__or4_4
X_20700_ _13113_/A VGND VGND VPWR VPWR _20700_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21680_ _21654_/A _19469_/Y VGND VGND VPWR VPWR _21680_/X sky130_fd_sc_hd__or2_4
XFILLER_212_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22926__A _23062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20631_ _17388_/B _20630_/Y _20621_/C VGND VGND VPWR VPWR _20631_/X sky130_fd_sc_hd__and3_4
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24356__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23350_ _23350_/A _25170_/Q VGND VGND VPWR VPWR _23363_/A sky130_fd_sc_hd__and2_4
XFILLER_20_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20562_ _18875_/A _18874_/X VGND VGND VPWR VPWR _20563_/B sky130_fd_sc_hd__nand2_4
XFILLER_177_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22301_ _22300_/Y _22287_/X _13116_/A _21292_/X VGND VGND VPWR VPWR _22301_/X sky130_fd_sc_hd__a2bb2o_4
X_23281_ _24642_/Q _21528_/B VGND VGND VPWR VPWR _23281_/X sky130_fd_sc_hd__or2_4
XFILLER_192_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20493_ _20529_/A _20492_/X VGND VGND VPWR VPWR _24079_/D sky130_fd_sc_hd__or2_4
XFILLER_192_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25020_ _25021_/CLK _15240_/Y HRESETn VGND VGND VPWR VPWR _25020_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12890__C _12588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22232_ _13538_/Y _22735_/B _21178_/X VGND VGND VPWR VPWR _22232_/X sky130_fd_sc_hd__a21o_4
XANTENNA__20059__A3 _15830_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22453__A1 _15003_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22453__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22661__A _22145_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22163_ _22163_/A _22701_/B VGND VGND VPWR VPWR _22163_/X sky130_fd_sc_hd__or2_4
XANTENNA__23991__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21114_ _21859_/A VGND VGND VPWR VPWR _21114_/X sky130_fd_sc_hd__buf_2
X_22094_ _14940_/A _22417_/B _21730_/A _22093_/X VGND VGND VPWR VPWR _22095_/C sky130_fd_sc_hd__a211o_4
XANTENNA__17474__B _17448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20216__B1 _19711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15891__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21045_ _21045_/A VGND VGND VPWR VPWR _21045_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_12_0_HCLK_A clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24804_ _24804_/CLK _15876_/X HRESETn VGND VGND VPWR VPWR _22901_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_203_0_HCLK clkbuf_8_202_0_HCLK/A VGND VGND VPWR VPWR _24985_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_216_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22996_ _22996_/A _22800_/B VGND VGND VPWR VPWR _22996_/X sky130_fd_sc_hd__or2_4
XFILLER_234_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24735_ _24737_/CLK _16026_/X HRESETn VGND VGND VPWR VPWR _24735_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_9_0_HCLK clkbuf_7_4_0_HCLK/X VGND VGND VPWR VPWR _23494_/CLK sky130_fd_sc_hd__clkbuf_1
X_21947_ _17720_/A _21947_/B VGND VGND VPWR VPWR _21949_/B sky130_fd_sc_hd__or2_4
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11700_ _11700_/A VGND VGND VPWR VPWR _21327_/A sky130_fd_sc_hd__inv_2
XFILLER_242_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12680_/A VGND VGND VPWR VPWR _12686_/A sky130_fd_sc_hd__buf_2
XFILLER_15_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ _22298_/A _21872_/X _21099_/X _21877_/X VGND VGND VPWR VPWR _21882_/A sky130_fd_sc_hd__a211o_4
X_24666_ _24667_/CLK _16216_/X HRESETn VGND VGND VPWR VPWR _22927_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_187_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _16715_/Y _20825_/X _24035_/Q _20828_/X VGND VGND VPWR VPWR _20830_/A sky130_fd_sc_hd__o22a_4
X_23617_ _23458_/CLK _19787_/X VGND VGND VPWR VPWR _23617_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24097__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24597_ _24597_/CLK _24597_/D HRESETn VGND VGND VPWR VPWR _24597_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14350_ _14344_/X _14348_/X _25485_/Q _14349_/X VGND VGND VPWR VPWR _14350_/X sky130_fd_sc_hd__o22a_4
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23548_ _24317_/CLK _19985_/X VGND VGND VPWR VPWR _19983_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_156_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24026__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13301_ _13369_/A _13296_/X _13300_/X VGND VGND VPWR VPWR _13302_/C sky130_fd_sc_hd__or3_4
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14281_ _14281_/A VGND VGND VPWR VPWR _14281_/Y sky130_fd_sc_hd__inv_2
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23479_ _23487_/CLK _23479_/D VGND VGND VPWR VPWR _23479_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13232_ _13225_/A VGND VGND VPWR VPWR _13438_/A sky130_fd_sc_hd__buf_2
X_16020_ HWDATA[21] VGND VGND VPWR VPWR _16020_/X sky130_fd_sc_hd__buf_2
X_25218_ _25224_/CLK _25218_/D HRESETn VGND VGND VPWR VPWR _14090_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__18648__B1 _16587_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13163_ _13155_/X _13160_/X _13162_/X VGND VGND VPWR VPWR _13163_/X sky130_fd_sc_hd__o21a_4
XFILLER_164_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25149_ _25146_/CLK _25149_/D HRESETn VGND VGND VPWR VPWR _25149_/Q sky130_fd_sc_hd__dfrtp_4
X_12114_ _24103_/Q _12120_/A VGND VGND VPWR VPWR _12125_/A sky130_fd_sc_hd__and2_4
X_13094_ _13068_/C _13068_/D VGND VGND VPWR VPWR _13095_/B sky130_fd_sc_hd__or2_4
X_17971_ _14639_/A VGND VGND VPWR VPWR _17972_/A sky130_fd_sc_hd__buf_2
XFILLER_78_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20207__B1 _19746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19710_ _13410_/B VGND VGND VPWR VPWR _19710_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15882__B1 _24801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12045_ _17436_/C VGND VGND VPWR VPWR _13457_/D sky130_fd_sc_hd__buf_2
X_16922_ _24698_/Q _16921_/Y _16152_/Y _16925_/A VGND VGND VPWR VPWR _16929_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15185__A _15185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_13_0_HCLK clkbuf_5_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19641_ _19641_/A VGND VGND VPWR VPWR _19641_/X sky130_fd_sc_hd__buf_2
X_16853_ _16852_/Y _16793_/X _16716_/X _16793_/X VGND VGND VPWR VPWR _16853_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15804_ _12296_/Y _15803_/X _15581_/X _15803_/X VGND VGND VPWR VPWR _24841_/D sky130_fd_sc_hd__a2bb2o_4
X_19572_ _19572_/A VGND VGND VPWR VPWR _22229_/B sky130_fd_sc_hd__buf_2
X_16784_ _16781_/Y _16779_/X _16783_/X _16779_/X VGND VGND VPWR VPWR _16784_/X sky130_fd_sc_hd__a2bb2o_4
X_13996_ _13990_/A VGND VGND VPWR VPWR _14028_/B sky130_fd_sc_hd__buf_2
XANTENNA__24867__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18523_ _18580_/A VGND VGND VPWR VPWR _18523_/X sky130_fd_sc_hd__buf_2
XFILLER_206_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15735_ HWDATA[16] VGND VGND VPWR VPWR _15735_/X sky130_fd_sc_hd__buf_2
X_12947_ _12781_/Y _12947_/B VGND VGND VPWR VPWR _12948_/B sky130_fd_sc_hd__or2_4
XFILLER_61_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13433__A _13433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18454_ _18745_/C VGND VGND VPWR VPWR _18774_/A sky130_fd_sc_hd__buf_2
X_15666_ _15666_/A VGND VGND VPWR VPWR _21323_/A sky130_fd_sc_hd__buf_2
X_12878_ _12878_/A _12878_/B VGND VGND VPWR VPWR _12880_/B sky130_fd_sc_hd__or2_4
XFILLER_222_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20930__A1 _16659_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17384_/X _17398_/X _24336_/Q _21000_/A _17401_/X VGND VGND VPWR VPWR _24337_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21650__A _13726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14617_ _14616_/X VGND VGND VPWR VPWR _14617_/Y sky130_fd_sc_hd__inv_2
X_11829_ _11829_/A VGND VGND VPWR VPWR _11829_/Y sky130_fd_sc_hd__inv_2
X_18385_ _24193_/Q VGND VGND VPWR VPWR _18385_/Y sky130_fd_sc_hd__inv_2
X_15597_ _15595_/Y _15596_/X _11730_/X _15596_/X VGND VGND VPWR VPWR _15597_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17336_ _17336_/A _17335_/Y VGND VGND VPWR VPWR _17338_/B sky130_fd_sc_hd__or2_4
XFILLER_147_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14548_ _14548_/A VGND VGND VPWR VPWR _14548_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20694__B1 _20690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17267_ _17228_/X VGND VGND VPWR VPWR _17284_/A sky130_fd_sc_hd__inv_2
X_14479_ _18951_/A VGND VGND VPWR VPWR _14479_/X sky130_fd_sc_hd__buf_2
X_19006_ _19006_/A VGND VGND VPWR VPWR _19006_/X sky130_fd_sc_hd__buf_2
X_16218_ _16217_/Y _16215_/X _15951_/X _16215_/X VGND VGND VPWR VPWR _16218_/X sky130_fd_sc_hd__a2bb2o_4
X_17198_ _17190_/X _17192_/X _17198_/C _17198_/D VGND VGND VPWR VPWR _17198_/X sky130_fd_sc_hd__or4_4
XANTENNA__22481__A _22638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16149_ _22191_/A VGND VGND VPWR VPWR _16149_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15873__B1 _15581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22738__A2 _22429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19908_ _19907_/Y _19905_/X _19817_/X _19905_/X VGND VGND VPWR VPWR _23575_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19064__B1 _19063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19839_ _23600_/Q VGND VGND VPWR VPWR _19839_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22850_ _12780_/Y _21437_/X _22849_/X _12547_/Y _21085_/X VGND VGND VPWR VPWR _22850_/X
+ sky130_fd_sc_hd__o32a_4
X_21801_ _21661_/A _21801_/B VGND VGND VPWR VPWR _21803_/B sky130_fd_sc_hd__or2_4
XFILLER_225_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22781_ _22781_/A _22781_/B _22781_/C _22780_/X VGND VGND VPWR VPWR _22781_/X sky130_fd_sc_hd__or4_4
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24537__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21732_ _18383_/Y _12057_/X _12104_/Y _21570_/X VGND VGND VPWR VPWR _21732_/X sky130_fd_sc_hd__o22a_4
X_24520_ _24520_/CLK _24520_/D HRESETn VGND VGND VPWR VPWR _24520_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_33_0_HCLK clkbuf_7_16_0_HCLK/X VGND VGND VPWR VPWR _23490_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22656__A _21077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_96_0_HCLK clkbuf_7_48_0_HCLK/X VGND VGND VPWR VPWR _24365_/CLK sky130_fd_sc_hd__clkbuf_1
X_21663_ _21472_/A _21663_/B _21662_/X VGND VGND VPWR VPWR _21663_/X sky130_fd_sc_hd__and3_4
X_24451_ _24419_/CLK _24451_/D HRESETn VGND VGND VPWR VPWR _14986_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24190__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20614_ _17399_/X VGND VGND VPWR VPWR _20615_/A sky130_fd_sc_hd__inv_2
X_23402_ _23675_/CLK _23402_/D VGND VGND VPWR VPWR _23402_/Q sky130_fd_sc_hd__dfxtp_4
X_24382_ _24725_/CLK _17138_/X HRESETn VGND VGND VPWR VPWR _24382_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22674__A1 _16587_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21594_ _21597_/A _21591_/X _22290_/A _21593_/X VGND VGND VPWR VPWR _21594_/X sky130_fd_sc_hd__o22a_4
XFILLER_177_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23333_ _16363_/A _23301_/B VGND VGND VPWR VPWR _23333_/X sky130_fd_sc_hd__or2_4
X_20545_ _14158_/Y _20543_/X _20600_/A _20544_/X VGND VGND VPWR VPWR _20546_/A sky130_fd_sc_hd__a211o_4
XANTENNA__17177__A2_N _17239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14174__A _20503_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23264_ _24443_/Q _21542_/X _22098_/X _23263_/X VGND VGND VPWR VPWR _23264_/X sky130_fd_sc_hd__a211o_4
X_20476_ _20476_/A _20476_/B _25254_/Q VGND VGND VPWR VPWR _20477_/C sky130_fd_sc_hd__or3_4
XANTENNA__25396__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22215_ _22210_/A _22215_/B VGND VGND VPWR VPWR _22215_/X sky130_fd_sc_hd__or2_4
X_25003_ _24953_/CLK _15327_/X HRESETn VGND VGND VPWR VPWR _25003_/Q sky130_fd_sc_hd__dfrtp_4
X_23195_ _23108_/X _23192_/Y _23155_/X _23194_/X VGND VGND VPWR VPWR _23195_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25325__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22146_ _21297_/Y VGND VGND VPWR VPWR _22146_/X sky130_fd_sc_hd__buf_2
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15864__B1 _15560_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19055__B1 _18985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22077_ _22373_/A _22075_/X _22077_/C VGND VGND VPWR VPWR _22077_/X sky130_fd_sc_hd__and3_4
XANTENNA__12678__B1 _12627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15734__A1_N _12547_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21028_ _11701_/X VGND VGND VPWR VPWR _22641_/B sky130_fd_sc_hd__buf_2
XFILLER_247_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18661__A1_N _16564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13850_ _13849_/X VGND VGND VPWR VPWR _13850_/X sky130_fd_sc_hd__buf_2
XANTENNA__23372__D scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24960__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12801_ _12800_/Y VGND VGND VPWR VPWR _12801_/X sky130_fd_sc_hd__buf_2
X_13781_ _13780_/Y VGND VGND VPWR VPWR _21379_/B sky130_fd_sc_hd__buf_2
XANTENNA__24278__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22979_ _22979_/A VGND VGND VPWR VPWR _22979_/Y sky130_fd_sc_hd__inv_2
X_15520_ _15518_/Y _15519_/X HADDR[9] _15519_/X VGND VGND VPWR VPWR _24934_/D sky130_fd_sc_hd__a2bb2o_4
X_12732_ _25399_/Q VGND VGND VPWR VPWR _12732_/Y sky130_fd_sc_hd__inv_2
X_24718_ _24737_/CLK _24718_/D HRESETn VGND VGND VPWR VPWR _24718_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_204_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24207__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16041__B1 _11739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15451_ _15451_/A VGND VGND VPWR VPWR _15451_/X sky130_fd_sc_hd__buf_2
X_12663_ _12564_/Y _12675_/A VGND VGND VPWR VPWR _12663_/X sky130_fd_sc_hd__or2_4
X_24649_ _24650_/CLK _24649_/D HRESETn VGND VGND VPWR VPWR _24649_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16564__A _16564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ HWDATA[6] VGND VGND VPWR VPWR _14403_/A sky130_fd_sc_hd__buf_2
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _18032_/A _18170_/B VGND VGND VPWR VPWR _18170_/X sky130_fd_sc_hd__or2_4
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_4_0_HCLK clkbuf_5_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _15087_/Y _15285_/Y VGND VGND VPWR VPWR _15382_/X sky130_fd_sc_hd__or2_4
XFILLER_230_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _25429_/Q VGND VGND VPWR VPWR _12594_/Y sky130_fd_sc_hd__inv_2
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ _17142_/A _17119_/X _17121_/C VGND VGND VPWR VPWR _24386_/D sky130_fd_sc_hd__and3_4
XFILLER_51_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14333_ _14337_/A VGND VGND VPWR VPWR _14345_/A sky130_fd_sc_hd__buf_2
XANTENNA__20517__C _20496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17052_ _17087_/A VGND VGND VPWR VPWR _17381_/B sky130_fd_sc_hd__inv_2
XFILLER_171_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14264_ _14264_/A VGND VGND VPWR VPWR _14264_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16003_ _24743_/Q VGND VGND VPWR VPWR _16003_/Y sky130_fd_sc_hd__inv_2
X_13215_ _13300_/A _13212_/X _13214_/X VGND VGND VPWR VPWR _13215_/X sky130_fd_sc_hd__and3_4
XANTENNA__15908__A _15908_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25066__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14195_ _20517_/A _14188_/X _13829_/X _14190_/X VGND VGND VPWR VPWR _14195_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_152_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13146_ _13170_/A _23794_/Q VGND VGND VPWR VPWR _13148_/B sky130_fd_sc_hd__or2_4
X_13077_ _12981_/C _13079_/B _13076_/Y VGND VGND VPWR VPWR _25346_/D sky130_fd_sc_hd__o21a_4
X_17954_ _17950_/X _17953_/X _18020_/A VGND VGND VPWR VPWR _17954_/X sky130_fd_sc_hd__o21a_4
XFILLER_151_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12332__A _24821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12028_ _12026_/Y _12027_/X _12029_/A _12027_/X VGND VGND VPWR VPWR _12028_/X sky130_fd_sc_hd__a2bb2o_4
X_16905_ _16144_/A _24266_/Q _16144_/Y _16904_/Y VGND VGND VPWR VPWR _16905_/X sky130_fd_sc_hd__o22a_4
XFILLER_239_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17885_ _17866_/A _17885_/B _17884_/Y VGND VGND VPWR VPWR _24260_/D sky130_fd_sc_hd__and3_4
XANTENNA__15870__A3 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15643__A _13797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16836_ _14895_/Y _16834_/X _15965_/A _16834_/X VGND VGND VPWR VPWR _24424_/D sky130_fd_sc_hd__a2bb2o_4
X_19624_ _13147_/B VGND VGND VPWR VPWR _19624_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16280__B1 _15991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19555_ _19549_/Y VGND VGND VPWR VPWR _19555_/X sky130_fd_sc_hd__buf_2
X_16767_ _16765_/Y _16766_/X _15748_/X _16766_/X VGND VGND VPWR VPWR _24457_/D sky130_fd_sc_hd__a2bb2o_4
X_13979_ _25237_/Q _25236_/Q _13979_/C _25234_/Q VGND VGND VPWR VPWR _13979_/X sky130_fd_sc_hd__or4_4
XANTENNA__24630__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18506_ _18497_/A _18506_/B _18506_/C VGND VGND VPWR VPWR _18506_/X sky130_fd_sc_hd__and3_4
X_15718_ _12515_/Y _15714_/X _15564_/X _15717_/X VGND VGND VPWR VPWR _15718_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19486_ _23720_/Q VGND VGND VPWR VPWR _22010_/B sky130_fd_sc_hd__inv_2
X_16698_ _16696_/Y _16692_/X _16601_/X _16697_/X VGND VGND VPWR VPWR _16698_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18437_ _16225_/Y _24173_/Q _16225_/Y _24173_/Q VGND VGND VPWR VPWR _18437_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15649_ _15648_/X VGND VGND VPWR VPWR _15649_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16474__A _24571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18368_ _18356_/X _18354_/Y _18367_/X _21979_/A _18357_/Y VGND VGND VPWR VPWR _24200_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17319_ _17179_/Y _17319_/B VGND VGND VPWR VPWR _17320_/C sky130_fd_sc_hd__nand2_4
X_18299_ _17731_/X _18298_/X _17731_/X _18298_/X VGND VGND VPWR VPWR _24215_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20330_ _22343_/B _20329_/X _19600_/A _20329_/X VGND VGND VPWR VPWR _23417_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22408__A1 _24265_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13522__A1_N SSn_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23100__A _23077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14897__B2 _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20261_ _21006_/B _20261_/B VGND VGND VPWR VPWR _20261_/X sky130_fd_sc_hd__or2_4
XFILLER_116_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15818__A _11706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22000_ _21642_/A VGND VGND VPWR VPWR _22735_/B sky130_fd_sc_hd__buf_2
XFILLER_89_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20192_ _20180_/A VGND VGND VPWR VPWR _20192_/X sky130_fd_sc_hd__buf_2
XFILLER_115_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24340__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12242__A _25437_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24789__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13321__A1 _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23951_ _23951_/CLK scl_i_S4 HRESETn VGND VGND VPWR VPWR _23952_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_229_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17752__B _16917_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24718__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22902_ _21424_/X _22901_/X _21427_/X _12521_/A _21428_/X VGND VGND VPWR VPWR _22903_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15553__A _15553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23882_ _23774_/CLK _23882_/D VGND VGND VPWR VPWR _19024_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_229_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16368__B _16792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16271__B1 _24645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22833_ _16675_/Y _22794_/A _15591_/Y _22832_/X VGND VGND VPWR VPWR _22833_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24371__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22764_ _22747_/Y _22752_/Y _22760_/Y _21445_/X _22763_/X VGND VGND VPWR VPWR _22764_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_198_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24300__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22386__A _22386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16023__B1 _15946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24503_ _25021_/CLK _24503_/D HRESETn VGND VGND VPWR VPWR _24503_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21290__A _21290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21715_ _21715_/A _14246_/A VGND VGND VPWR VPWR _21719_/A sky130_fd_sc_hd__or2_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22817__C _22817_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19760__B2 _19740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22695_ _22695_/A _22619_/B VGND VGND VPWR VPWR _22695_/X sky130_fd_sc_hd__and2_4
X_25483_ _25158_/CLK _25483_/D HRESETn VGND VGND VPWR VPWR _25483_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21646_ _23685_/Q _21959_/B _19538_/A _22397_/B VGND VGND VPWR VPWR _21646_/X sky130_fd_sc_hd__o22a_4
X_24434_ _24462_/CLK _16815_/X HRESETn VGND VGND VPWR VPWR _14964_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_12_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22647__A1 _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12731__A1_N _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21577_ _21576_/X VGND VGND VPWR VPWR _21577_/Y sky130_fd_sc_hd__inv_2
X_24365_ _24365_/CLK _24365_/D HRESETn VGND VGND VPWR VPWR _23078_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25506__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20528_ _15451_/A _20514_/C _20526_/Y _20527_/X VGND VGND VPWR VPWR _20528_/X sky130_fd_sc_hd__a211o_4
X_23316_ _23316_/A _23156_/X VGND VGND VPWR VPWR _23316_/X sky130_fd_sc_hd__or2_4
X_24296_ _24297_/CLK _24296_/D HRESETn VGND VGND VPWR VPWR _17530_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15728__A _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20459_ _14530_/A _20458_/Y VGND VGND VPWR VPWR _20459_/Y sky130_fd_sc_hd__nor2_4
X_23247_ _23228_/X _23231_/X _23235_/Y _23246_/X VGND VGND VPWR VPWR HRDATA[28] sky130_fd_sc_hd__a211o_4
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14632__A _14630_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13000_ _13000_/A _12285_/Y _13059_/A _13000_/D VGND VGND VPWR VPWR _13001_/A sky130_fd_sc_hd__or4_4
XANTENNA__15043__A1_N _15249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23178_ _23178_/A VGND VGND VPWR VPWR _23178_/X sky130_fd_sc_hd__buf_2
XFILLER_133_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22129_ _21537_/X VGND VGND VPWR VPWR _22129_/X sky130_fd_sc_hd__buf_2
XANTENNA__13248__A _13285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14951_ _14951_/A VGND VGND VPWR VPWR _15065_/A sky130_fd_sc_hd__buf_2
XFILLER_248_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16559__A _24539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24459__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13902_ _13902_/A VGND VGND VPWR VPWR _14232_/B sky130_fd_sc_hd__inv_2
XFILLER_236_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17670_ _17670_/A _17670_/B VGND VGND VPWR VPWR _17670_/X sky130_fd_sc_hd__or2_4
XFILLER_236_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14882_ _15249_/A _24425_/Q _15249_/A _24425_/Q VGND VGND VPWR VPWR _14882_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16262__B1 _15976_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16621_ _14756_/A _16171_/X _13577_/B VGND VGND VPWR VPWR _16621_/X sky130_fd_sc_hd__o21a_4
X_13833_ _13559_/Y _13828_/X _13788_/X _13832_/X VGND VGND VPWR VPWR _13833_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13076__B1 _13019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22335__B1 _22322_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18774__A _18774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19340_ _17948_/B VGND VGND VPWR VPWR _19340_/Y sky130_fd_sc_hd__inv_2
X_16552_ _24542_/Q VGND VGND VPWR VPWR _16552_/Y sky130_fd_sc_hd__inv_2
XFILLER_244_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13764_ _13763_/X VGND VGND VPWR VPWR _13772_/C sky130_fd_sc_hd__buf_2
XFILLER_16_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24041__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15503_ _24940_/Q VGND VGND VPWR VPWR _15503_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12715_ _12714_/X VGND VGND VPWR VPWR _12715_/Y sky130_fd_sc_hd__inv_2
X_19271_ _21249_/B _19266_/X _19091_/X _19253_/Y VGND VGND VPWR VPWR _19271_/X sky130_fd_sc_hd__a2bb2o_4
X_16483_ HWDATA[21] VGND VGND VPWR VPWR _16483_/X sky130_fd_sc_hd__buf_2
X_13695_ _13678_/A _13678_/B VGND VGND VPWR VPWR _13695_/Y sky130_fd_sc_hd__nand2_4
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18222_ _18222_/A _23835_/Q VGND VGND VPWR VPWR _18222_/X sky130_fd_sc_hd__or2_4
XFILLER_188_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15434_ _13913_/X _15432_/X _15427_/X _24974_/Q _15433_/X VGND VGND VPWR VPWR _15434_/X
+ sky130_fd_sc_hd__a32o_4
X_12646_ _12638_/X VGND VGND VPWR VPWR _12650_/B sky130_fd_sc_hd__inv_2
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ _18053_/A _23773_/Q VGND VGND VPWR VPWR _18155_/B sky130_fd_sc_hd__or2_4
XFILLER_157_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15365_ _15352_/A _15361_/X _15364_/Y VGND VGND VPWR VPWR _24993_/D sky130_fd_sc_hd__and3_4
XFILLER_8_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12577_ _12568_/X _12577_/B _12573_/X _12577_/D VGND VGND VPWR VPWR _12577_/X sky130_fd_sc_hd__or4_4
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17104_ _16984_/Y _17103_/X VGND VGND VPWR VPWR _17104_/Y sky130_fd_sc_hd__nand2_4
X_14316_ _14315_/X VGND VGND VPWR VPWR _14316_/Y sky130_fd_sc_hd__inv_2
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18084_ _18222_/A _23879_/Q VGND VGND VPWR VPWR _18085_/C sky130_fd_sc_hd__or2_4
X_15296_ _15296_/A _15296_/B _15068_/Y _15390_/A VGND VGND VPWR VPWR _15299_/B sky130_fd_sc_hd__or4_4
XFILLER_8_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17035_ _17035_/A _16971_/Y _16975_/Y _16957_/Y VGND VGND VPWR VPWR _17042_/A sky130_fd_sc_hd__or4_4
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14247_ _14247_/A VGND VGND VPWR VPWR _14247_/X sky130_fd_sc_hd__buf_2
XFILLER_7_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15638__A _14366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14882__A1_N _15249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14542__A HREADY VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18014__A _18014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14178_ _15984_/A _14178_/B _14365_/C _14365_/D VGND VGND VPWR VPWR _14179_/B sky130_fd_sc_hd__or4_4
XANTENNA__15828__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16893__A2_N _24274_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13158__A _13157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13129_ _13129_/A VGND VGND VPWR VPWR _13129_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19019__B1 _18948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18986_ _18986_/A VGND VGND VPWR VPWR _18986_/X sky130_fd_sc_hd__buf_2
XANTENNA__24882__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14897__A1_N _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17937_ _17949_/A _17937_/B VGND VGND VPWR VPWR _17938_/C sky130_fd_sc_hd__or2_4
XANTENNA__24811__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17868_ _17867_/X VGND VGND VPWR VPWR _17868_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24129__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16253__B1 _16059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19607_ _19598_/Y VGND VGND VPWR VPWR _19607_/X sky130_fd_sc_hd__buf_2
X_16819_ _14936_/Y _16816_/X HWDATA[17] _16816_/X VGND VGND VPWR VPWR _24431_/D sky130_fd_sc_hd__a2bb2o_4
X_17799_ _24283_/Q _17798_/Y VGND VGND VPWR VPWR _17801_/B sky130_fd_sc_hd__or2_4
XFILLER_19_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19538_ _19538_/A VGND VGND VPWR VPWR _19538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12814__B1 _12813_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21822__B _21649_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16005__B1 _16004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19469_ _19469_/A VGND VGND VPWR VPWR _19469_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21500_ _21274_/X VGND VGND VPWR VPWR _22393_/A sky130_fd_sc_hd__buf_2
XFILLER_195_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13621__A _13579_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22480_ _22769_/A _22479_/X VGND VGND VPWR VPWR _22480_/X sky130_fd_sc_hd__and2_4
XFILLER_195_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21431_ _22189_/A VGND VGND VPWR VPWR _21431_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_107_0_HCLK clkbuf_7_53_0_HCLK/X VGND VGND VPWR VPWR _24662_/CLK sky130_fd_sc_hd__clkbuf_1
X_24150_ _24146_/CLK _24150_/D HRESETn VGND VGND VPWR VPWR _24150_/Q sky130_fd_sc_hd__dfrtp_4
X_21362_ _21361_/X VGND VGND VPWR VPWR _21362_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21852__A2 _12086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20313_ _20306_/X _19573_/X _13829_/A _22003_/A _20310_/X VGND VGND VPWR VPWR _23423_/D
+ sky130_fd_sc_hd__a32o_4
X_23101_ _23101_/A _22897_/X VGND VGND VPWR VPWR _23101_/X sky130_fd_sc_hd__or2_4
X_24081_ _24074_/CLK _24081_/D HRESETn VGND VGND VPWR VPWR _20524_/B sky130_fd_sc_hd__dfrtp_4
X_21293_ _21519_/A VGND VGND VPWR VPWR _21864_/B sky130_fd_sc_hd__buf_2
X_23032_ _23031_/X VGND VGND VPWR VPWR _23032_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17269__C1 _17268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20244_ _20240_/Y _20243_/X _16854_/X _20243_/X VGND VGND VPWR VPWR _23450_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_150_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15819__B1 _24831_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20175_ _23475_/Q VGND VGND VPWR VPWR _21263_/B sky130_fd_sc_hd__inv_2
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24983_ _24985_/CLK _24983_/D HRESETn VGND VGND VPWR VPWR _24983_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24552__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22565__B1 _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23934_ _23951_/CLK _20985_/X HRESETn VGND VGND VPWR VPWR _20986_/A sky130_fd_sc_hd__dfstp_4
XFILLER_85_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23865_ _24413_/CLK _19077_/X VGND VGND VPWR VPWR _19076_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22816_ _22816_/A VGND VGND VPWR VPWR _22817_/C sky130_fd_sc_hd__buf_2
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23796_ _23859_/CLK _19269_/X VGND VGND VPWR VPWR _23796_/Q sky130_fd_sc_hd__dfxtp_4
X_25535_ _25533_/CLK _11731_/X HRESETn VGND VGND VPWR VPWR _25535_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22747_ _22632_/A _22747_/B VGND VGND VPWR VPWR _22747_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12281__B2 _24831_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12500_ _12613_/A VGND VGND VPWR VPWR _12500_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13480_ _13480_/A VGND VGND VPWR VPWR _13480_/Y sky130_fd_sc_hd__inv_2
X_25466_ _25466_/CLK _25466_/D HRESETn VGND VGND VPWR VPWR _12159_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_200_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_66_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_66_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22678_ _16272_/X _22678_/B VGND VGND VPWR VPWR _22678_/Y sky130_fd_sc_hd__nor2_4
XFILLER_232_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12431_ _12428_/C _12428_/D VGND VGND VPWR VPWR _12431_/X sky130_fd_sc_hd__or2_4
X_24417_ _24574_/CLK _16848_/X HRESETn VGND VGND VPWR VPWR _16847_/A sky130_fd_sc_hd__dfrtp_4
X_21629_ _22225_/A VGND VGND VPWR VPWR _21771_/A sky130_fd_sc_hd__buf_2
XANTENNA__25340__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25397_ _25397_/CLK _12861_/X HRESETn VGND VGND VPWR VPWR _25397_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15150_ _15150_/A VGND VGND VPWR VPWR _15150_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12362_ _25365_/Q VGND VGND VPWR VPWR _12990_/A sky130_fd_sc_hd__inv_2
X_24348_ _24346_/CLK _17365_/X HRESETn VGND VGND VPWR VPWR _24348_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14101_ _25223_/Q VGND VGND VPWR VPWR _14108_/A sky130_fd_sc_hd__inv_2
X_12293_ _24830_/Q VGND VGND VPWR VPWR _12293_/Y sky130_fd_sc_hd__inv_2
X_15081_ _24590_/Q VGND VGND VPWR VPWR _15081_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24279_ _24278_/CLK _24279_/D HRESETn VGND VGND VPWR VPWR _24279_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14032_ _14032_/A VGND VGND VPWR VPWR _14032_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18769__A _18769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18840_ _18836_/X _18840_/B _18838_/X _18839_/X VGND VGND VPWR VPWR _18840_/X sky130_fd_sc_hd__or4_4
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18771_ _18752_/A _18769_/X _18771_/C VGND VGND VPWR VPWR _18771_/X sky130_fd_sc_hd__and3_4
X_15983_ _23138_/A VGND VGND VPWR VPWR _15983_/X sky130_fd_sc_hd__buf_2
XANTENNA__24293__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22186__A1_N _20510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22556__B1 _12511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17722_ _24214_/Q VGND VGND VPWR VPWR _17723_/A sky130_fd_sc_hd__inv_2
XFILLER_236_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15193__A _15165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14934_ _14923_/X _14934_/B _14930_/X _14934_/D VGND VGND VPWR VPWR _14935_/D sky130_fd_sc_hd__or4_4
XFILLER_36_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24222__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17653_ _17569_/D _17637_/B _17604_/X _17651_/B VGND VGND VPWR VPWR _17653_/X sky130_fd_sc_hd__a211o_4
X_14865_ _14859_/C _23994_/Q VGND VGND VPWR VPWR _14865_/X sky130_fd_sc_hd__or2_4
XFILLER_63_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16604_ _16603_/Y _16598_/X _16518_/X _16598_/X VGND VGND VPWR VPWR _16604_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13816_ _13531_/Y _13813_/X _11748_/X _13813_/X VGND VGND VPWR VPWR _13816_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15921__A _15670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17584_ _17563_/Y _17545_/Y _17584_/C _17583_/X VGND VGND VPWR VPWR _17584_/X sky130_fd_sc_hd__or4_4
XFILLER_217_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25499__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14796_ _14796_/A _14796_/B _14811_/A VGND VGND VPWR VPWR _14796_/X sky130_fd_sc_hd__or3_4
X_19323_ _19319_/Y _19322_/X _19301_/X _19322_/X VGND VGND VPWR VPWR _23778_/D sky130_fd_sc_hd__a2bb2o_4
X_16535_ _16534_/Y _16454_/A _16358_/X _16454_/A VGND VGND VPWR VPWR _16535_/X sky130_fd_sc_hd__a2bb2o_4
X_13747_ _13746_/X VGND VGND VPWR VPWR _13747_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15640__B _15640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17735__B1 _17731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19254_ _19253_/Y VGND VGND VPWR VPWR _19254_/X sky130_fd_sc_hd__buf_2
X_16466_ _24574_/Q VGND VGND VPWR VPWR _16466_/Y sky130_fd_sc_hd__inv_2
X_13678_ _13678_/A _13678_/B VGND VGND VPWR VPWR _13679_/A sky130_fd_sc_hd__or2_4
X_18205_ _18044_/A _18205_/B _18204_/X VGND VGND VPWR VPWR _18205_/X sky130_fd_sc_hd__or3_4
XANTENNA__22124__A1_N _20517_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15417_ _15417_/A _15417_/B VGND VGND VPWR VPWR _15418_/B sky130_fd_sc_hd__or2_4
XFILLER_31_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12629_ _12628_/X VGND VGND VPWR VPWR _25429_/D sky130_fd_sc_hd__inv_2
X_19185_ _19184_/X VGND VGND VPWR VPWR _19191_/A sky130_fd_sc_hd__buf_2
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25081__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16397_ HWDATA[19] VGND VGND VPWR VPWR _16397_/X sky130_fd_sc_hd__buf_2
XFILLER_129_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14191__A1_N _20496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18136_ _18104_/A _18136_/B VGND VGND VPWR VPWR _18137_/C sky130_fd_sc_hd__or2_4
X_15348_ _15293_/B _15347_/X VGND VGND VPWR VPWR _15349_/A sky130_fd_sc_hd__or2_4
XANTENNA__25010__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21834__A2 _21832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18067_ _18104_/A _23759_/Q VGND VGND VPWR VPWR _18067_/X sky130_fd_sc_hd__or2_4
X_15279_ _15241_/A _15273_/B _15278_/Y VGND VGND VPWR VPWR _15279_/X sky130_fd_sc_hd__and3_4
XFILLER_171_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17018_ _17087_/A VGND VGND VPWR VPWR _17070_/A sky130_fd_sc_hd__buf_2
XFILLER_132_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19660__B1 _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18969_ _18968_/Y _18966_/X _18948_/X _18966_/X VGND VGND VPWR VPWR _18969_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_239_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21980_ _21983_/A _23421_/Q _18350_/A _20320_/Y VGND VGND VPWR VPWR _21980_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21833__A _21325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20931_ _20931_/A VGND VGND VPWR VPWR _20931_/Y sky130_fd_sc_hd__inv_2
XFILLER_215_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20862_ _20862_/A _20862_/B _20862_/C VGND VGND VPWR VPWR _20862_/X sky130_fd_sc_hd__and3_4
X_23650_ _25326_/CLK _23650_/D VGND VGND VPWR VPWR _13152_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23945__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22601_ _21077_/A _22598_/X _21114_/X _22600_/X VGND VGND VPWR VPWR _22601_/Y sky130_fd_sc_hd__a22oi_4
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20793_ _20793_/A _20793_/B VGND VGND VPWR VPWR _20793_/Y sky130_fd_sc_hd__nor2_4
X_23581_ _24297_/CLK _19892_/X VGND VGND VPWR VPWR _19890_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13460__B1 _13459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25320_ _25158_/CLK _25320_/D HRESETn VGND VGND VPWR VPWR _25320_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22532_ _24590_/Q _22532_/B VGND VGND VPWR VPWR _22539_/B sky130_fd_sc_hd__or2_4
X_25251_ _25230_/CLK _13857_/X HRESETn VGND VGND VPWR VPWR _20673_/A sky130_fd_sc_hd__dfrtp_4
X_22463_ _22696_/B _22461_/X _13800_/X _22462_/X VGND VGND VPWR VPWR _22463_/X sky130_fd_sc_hd__o22a_4
XFILLER_183_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24202_ _25081_/CLK _18364_/X HRESETn VGND VGND VPWR VPWR _18361_/A sky130_fd_sc_hd__dfrtp_4
X_21414_ _21410_/X _21413_/X _14672_/A VGND VGND VPWR VPWR _21414_/X sky130_fd_sc_hd__o21a_4
X_22394_ _22394_/A _22394_/B _22335_/X _22393_/Y VGND VGND VPWR VPWR _22394_/X sky130_fd_sc_hd__or4_4
X_25182_ _25479_/CLK _25182_/D HRESETn VGND VGND VPWR VPWR _13508_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_148_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14960__B1 _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21345_ _21720_/A VGND VGND VPWR VPWR _21345_/Y sky130_fd_sc_hd__inv_2
X_24133_ _24133_/CLK _24133_/D HRESETn VGND VGND VPWR VPWR _24133_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12499__A2_N _24866_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23027__B2 _22846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14182__A _14182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21276_ _13804_/Y VGND VGND VPWR VPWR _22582_/A sky130_fd_sc_hd__buf_2
X_24064_ _24060_/CLK _20955_/X HRESETn VGND VGND VPWR VPWR _20953_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24733__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_HCLK clkbuf_3_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_20227_ _20227_/A VGND VGND VPWR VPWR _20227_/X sky130_fd_sc_hd__buf_2
X_23015_ _22946_/A _23015_/B _23014_/X VGND VGND VPWR VPWR _23015_/X sky130_fd_sc_hd__and3_4
XFILLER_150_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16465__B1 _16464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17662__C1 _17593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20158_ _20158_/A VGND VGND VPWR VPWR _20158_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12980_ _12980_/A VGND VGND VPWR VPWR _12981_/D sky130_fd_sc_hd__inv_2
X_20089_ _24413_/Q VGND VGND VPWR VPWR _20089_/X sky130_fd_sc_hd__buf_2
X_24966_ _24967_/CLK _15446_/X HRESETn VGND VGND VPWR VPWR _13888_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11931_ _11931_/A VGND VGND VPWR VPWR _11934_/A sky130_fd_sc_hd__inv_2
X_23917_ _25308_/CLK _18926_/X VGND VGND VPWR VPWR _23917_/Q sky130_fd_sc_hd__dfxtp_4
X_24897_ _24037_/CLK _24897_/D HRESETn VGND VGND VPWR VPWR _15625_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22558__B _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15741__A HWDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14650_ _14650_/A VGND VGND VPWR VPWR _19026_/C sky130_fd_sc_hd__buf_2
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18755__C _18692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11862_ _11801_/Y _11864_/B _25519_/Q _11861_/Y VGND VGND VPWR VPWR _11862_/X sky130_fd_sc_hd__o22a_4
X_23848_ _23831_/CLK _19127_/X VGND VGND VPWR VPWR _18053_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_45_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _17943_/A _19116_/B _17943_/A _19116_/B VGND VGND VPWR VPWR _14787_/A sky130_fd_sc_hd__a2bb2o_4
XPHY_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _14557_/A _14557_/B VGND VGND VPWR VPWR _14581_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__18474__D _18400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25521__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _13459_/A VGND VGND VPWR VPWR _11793_/X sky130_fd_sc_hd__buf_2
X_23779_ _24252_/CLK _19318_/X VGND VGND VPWR VPWR _18202_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16320_ HWDATA[16] VGND VGND VPWR VPWR _16320_/X sky130_fd_sc_hd__buf_2
XANTENNA__13261__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ _13530_/Y _25088_/Q _13531_/Y _25094_/Q VGND VGND VPWR VPWR _13541_/A sky130_fd_sc_hd__a2bb2o_4
X_25518_ _25499_/CLK _25518_/D HRESETn VGND VGND VPWR VPWR _11796_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_198_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16251_ _22163_/A VGND VGND VPWR VPWR _16251_/Y sky130_fd_sc_hd__inv_2
X_13463_ _13462_/X VGND VGND VPWR VPWR _13464_/A sky130_fd_sc_hd__inv_2
X_25449_ _24765_/CLK _25449_/D HRESETn VGND VGND VPWR VPWR _12175_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_158_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15202_ _15201_/X VGND VGND VPWR VPWR _25030_/D sky130_fd_sc_hd__inv_2
X_12414_ _12402_/B _12378_/X _12240_/Y VGND VGND VPWR VPWR _12414_/X sky130_fd_sc_hd__o21a_4
X_16182_ _16182_/A VGND VGND VPWR VPWR _16540_/B sky130_fd_sc_hd__buf_2
X_13394_ _13394_/A _13394_/B _13394_/C VGND VGND VPWR VPWR _13402_/B sky130_fd_sc_hd__or3_4
XFILLER_182_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_153_0_HCLK clkbuf_7_76_0_HCLK/X VGND VGND VPWR VPWR _25466_/CLK sky130_fd_sc_hd__clkbuf_1
X_15133_ _15361_/A _24597_/Q _24997_/Q _15084_/Y VGND VGND VPWR VPWR _15136_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12345_ _13046_/A _24837_/Q _25356_/Q _12296_/Y VGND VGND VPWR VPWR _12348_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23018__B2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15064_ _15059_/X _15063_/X VGND VGND VPWR VPWR _15064_/X sky130_fd_sc_hd__or2_4
X_19941_ _19946_/A VGND VGND VPWR VPWR _19941_/X sky130_fd_sc_hd__buf_2
X_12276_ _12271_/X _12275_/X VGND VGND VPWR VPWR _12402_/B sky130_fd_sc_hd__or2_4
XFILLER_107_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20822__A _20822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24474__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12714__C1 _12641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14015_ _14014_/X VGND VGND VPWR VPWR _14536_/B sky130_fd_sc_hd__inv_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19872_ _19871_/Y _19869_/X _19620_/X _19869_/X VGND VGND VPWR VPWR _19872_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19642__B1 _19540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24403__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18823_ _18616_/X _18823_/B VGND VGND VPWR VPWR _18824_/C sky130_fd_sc_hd__or2_4
XFILLER_96_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22529__B1 _22508_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15966_ _12178_/Y _15964_/X _15965_/X _15964_/X VGND VGND VPWR VPWR _15966_/X sky130_fd_sc_hd__a2bb2o_4
X_18754_ _18753_/X VGND VGND VPWR VPWR _24146_/D sky130_fd_sc_hd__inv_2
XFILLER_236_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16208__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14917_ _14917_/A VGND VGND VPWR VPWR _14917_/Y sky130_fd_sc_hd__inv_2
X_17705_ _17704_/X VGND VGND VPWR VPWR _17706_/A sky130_fd_sc_hd__inv_2
XANTENNA__17850__B _17555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15897_ _12784_/Y _15896_/X _15623_/X _15896_/X VGND VGND VPWR VPWR _15897_/X sky130_fd_sc_hd__a2bb2o_4
X_18685_ _18633_/A _18783_/A _18610_/A _18786_/A VGND VGND VPWR VPWR _18686_/D sky130_fd_sc_hd__or4_4
XFILLER_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14848_ _14848_/A VGND VGND VPWR VPWR _14848_/Y sky130_fd_sc_hd__inv_2
X_17636_ _17636_/A VGND VGND VPWR VPWR _17636_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17567_ _24306_/Q VGND VGND VPWR VPWR _17569_/C sky130_fd_sc_hd__inv_2
XFILLER_63_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14779_ _14769_/B _14777_/X _14778_/Y VGND VGND VPWR VPWR _14779_/X sky130_fd_sc_hd__o21a_4
XFILLER_210_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13171__A _13168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16518_ _14400_/A VGND VGND VPWR VPWR _16518_/X sky130_fd_sc_hd__buf_2
X_19306_ _19299_/Y VGND VGND VPWR VPWR _19306_/X sky130_fd_sc_hd__buf_2
X_17498_ _11725_/Y _24307_/Q _11725_/Y _24307_/Q VGND VGND VPWR VPWR _17506_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16449_ _16441_/X _16448_/X _16361_/X _16448_/X VGND VGND VPWR VPWR _24579_/D sky130_fd_sc_hd__a2bb2o_4
X_19237_ _23808_/Q VGND VGND VPWR VPWR _22058_/B sky130_fd_sc_hd__inv_2
XANTENNA__23257__A1 _12204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16931__B2 _17744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19168_ _19167_/Y _19165_/X _19122_/X _19165_/X VGND VGND VPWR VPWR _23833_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18119_ _18222_/A _19037_/A VGND VGND VPWR VPWR _18120_/C sky130_fd_sc_hd__or2_4
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19099_ _19098_/Y _19096_/X _18981_/X _19096_/X VGND VGND VPWR VPWR _23857_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21130_ _22466_/A _21130_/B _21129_/X VGND VGND VPWR VPWR _21130_/X sky130_fd_sc_hd__and3_4
XANTENNA__16695__B1 _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22768__B1 _24836_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21061_ _21098_/A VGND VGND VPWR VPWR _21061_/X sky130_fd_sc_hd__buf_2
XFILLER_160_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18827__A2_N _18769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24144__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20012_ _20012_/A VGND VGND VPWR VPWR _20012_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24820_ _24819_/CLK _15835_/X HRESETn VGND VGND VPWR VPWR _24820_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_246_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24751_ _25375_/CLK _24751_/D HRESETn VGND VGND VPWR VPWR _24751_/Q sky130_fd_sc_hd__dfrtp_4
X_21963_ _14606_/A _19594_/Y _21964_/A _19592_/Y VGND VGND VPWR VPWR _21963_/X sky130_fd_sc_hd__o22a_4
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23702_ _24208_/CLK _19537_/X VGND VGND VPWR VPWR _23702_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15561__A _15553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20914_ _20914_/A VGND VGND VPWR VPWR _24054_/D sky130_fd_sc_hd__inv_2
XFILLER_242_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24682_ _24681_/CLK _16162_/X HRESETn VGND VGND VPWR VPWR _21435_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21894_ _22386_/A _21894_/B VGND VGND VPWR VPWR _21894_/X sky130_fd_sc_hd__or2_4
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23633_ _23458_/CLK _19744_/X VGND VGND VPWR VPWR _23633_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20844_/X VGND VGND VPWR VPWR _20845_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13081__A _13085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23564_ _24297_/CLK _23564_/D VGND VGND VPWR VPWR _19934_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20776_ _13108_/B VGND VGND VPWR VPWR _20776_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25303_ _25492_/CLK _25303_/D HRESETn VGND VGND VPWR VPWR _13523_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22515_ _22515_/A VGND VGND VPWR VPWR _22515_/X sky130_fd_sc_hd__buf_2
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23495_ _23487_/CLK _23495_/D VGND VGND VPWR VPWR _20123_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24985__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25234_ _23976_/CLK _14071_/X HRESETn VGND VGND VPWR VPWR _25234_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22446_ _21439_/X VGND VGND VPWR VPWR _22769_/A sky130_fd_sc_hd__buf_2
XFILLER_109_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11724__A1_N _11720_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24914__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25165_ _25164_/CLK _25165_/D HRESETn VGND VGND VPWR VPWR _25165_/Q sky130_fd_sc_hd__dfrtp_4
X_22377_ _22373_/X _22376_/X _14666_/X VGND VGND VPWR VPWR _22377_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__19872__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_226_0_HCLK clkbuf_8_227_0_HCLK/A VGND VGND VPWR VPWR _25249_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_151_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12130_ _12115_/A _12125_/A _12129_/Y VGND VGND VPWR VPWR _12131_/A sky130_fd_sc_hd__o21a_4
X_24116_ _24209_/CLK _18899_/Y HRESETn VGND VGND VPWR VPWR _11929_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16686__B1 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21328_ _21327_/X VGND VGND VPWR VPWR _21582_/A sky130_fd_sc_hd__buf_2
X_25096_ _24188_/CLK _25096_/D HRESETn VGND VGND VPWR VPWR _13555_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_190_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12361__A2_N _24823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22759__B1 _21832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12061_ _12049_/Y _12060_/X _11761_/X _12060_/X VGND VGND VPWR VPWR _25486_/D sky130_fd_sc_hd__a2bb2o_4
X_21259_ _22056_/A _21259_/B VGND VGND VPWR VPWR _21259_/X sky130_fd_sc_hd__or2_4
X_24047_ _24427_/CLK _20882_/X HRESETn VGND VGND VPWR VPWR _24047_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23375__D _20822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15820_ _15820_/A VGND VGND VPWR VPWR _15820_/X sky130_fd_sc_hd__buf_2
XFILLER_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15751_ _12511_/Y _15750_/X _13818_/X _15750_/X VGND VGND VPWR VPWR _24865_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21473__A _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12963_ _12952_/A _12963_/B _12962_/Y VGND VGND VPWR VPWR _25370_/D sky130_fd_sc_hd__and3_4
X_24949_ _25285_/CLK _24949_/D HRESETn VGND VGND VPWR VPWR _14664_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_38_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14702_ _14701_/Y VGND VGND VPWR VPWR _14702_/X sky130_fd_sc_hd__buf_2
XFILLER_234_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11914_ _19613_/A VGND VGND VPWR VPWR _11914_/Y sky130_fd_sc_hd__inv_2
X_18470_ _18470_/A VGND VGND VPWR VPWR _18479_/B sky130_fd_sc_hd__inv_2
X_15682_ _24784_/Q _15679_/Y _15681_/X _13579_/B VGND VGND VPWR VPWR _15686_/B sky130_fd_sc_hd__a211o_4
X_12894_ _12896_/B VGND VGND VPWR VPWR _12894_/Y sky130_fd_sc_hd__inv_2
X_17421_ _14407_/A VGND VGND VPWR VPWR _17421_/X sky130_fd_sc_hd__buf_2
X_14633_ _13596_/B _14632_/Y _18009_/A _14632_/Y VGND VGND VPWR VPWR _14633_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_233_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11845_ _11843_/A _11844_/A _13686_/A _11844_/Y VGND VGND VPWR VPWR _11846_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12227__B2 _24762_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17352_ _17358_/A _17352_/B _17352_/C VGND VGND VPWR VPWR _17352_/X sky130_fd_sc_hd__or3_4
XPHY_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14563_/X _14544_/X _25276_/Q VGND VGND VPWR VPWR _14564_/Y sky130_fd_sc_hd__o21ai_4
XPHY_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _11772_/Y _11766_/X _11775_/X _11766_/X VGND VGND VPWR VPWR _11776_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16303_/A VGND VGND VPWR VPWR _16303_/Y sky130_fd_sc_hd__inv_2
X_13515_ _13514_/X VGND VGND VPWR VPWR _13515_/Y sky130_fd_sc_hd__inv_2
X_17283_ _17230_/X _17281_/X _17282_/X VGND VGND VPWR VPWR _24368_/D sky130_fd_sc_hd__and3_4
X_14495_ _23957_/Q VGND VGND VPWR VPWR _14495_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_36_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19022_ _19022_/A VGND VGND VPWR VPWR _19022_/Y sky130_fd_sc_hd__inv_2
X_16234_ _16232_/Y _16230_/X _16233_/X _16230_/X VGND VGND VPWR VPWR _16234_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17531__A1_N _25521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13446_ _13227_/X _13446_/B VGND VGND VPWR VPWR _13446_/X sky130_fd_sc_hd__or2_4
XFILLER_167_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24655__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16165_ _14775_/Y _16165_/B VGND VGND VPWR VPWR _16173_/A sky130_fd_sc_hd__and2_4
X_13377_ _13345_/A _13373_/X _13376_/X VGND VGND VPWR VPWR _13377_/X sky130_fd_sc_hd__or3_4
XFILLER_186_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15116_ _15116_/A _15116_/B _15102_/X _15115_/X VGND VGND VPWR VPWR _15116_/X sky130_fd_sc_hd__or4_4
X_12328_ _12289_/X _12328_/B _12328_/C _12328_/D VGND VGND VPWR VPWR _12370_/A sky130_fd_sc_hd__or4_4
X_16096_ _23193_/A VGND VGND VPWR VPWR _16096_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15047_ _15047_/A VGND VGND VPWR VPWR _15047_/Y sky130_fd_sc_hd__inv_2
X_19924_ _19924_/A VGND VGND VPWR VPWR _19924_/Y sky130_fd_sc_hd__inv_2
X_12259_ _12253_/X _12255_/X _12259_/C _12259_/D VGND VGND VPWR VPWR _12259_/X sky130_fd_sc_hd__or4_4
XFILLER_69_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19855_ _19939_/A _18279_/X _19455_/X VGND VGND VPWR VPWR _19856_/A sky130_fd_sc_hd__or3_4
X_18806_ _18686_/A _18809_/B _18709_/X VGND VGND VPWR VPWR _18806_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_95_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19786_ _23617_/Q VGND VGND VPWR VPWR _19786_/Y sky130_fd_sc_hd__inv_2
X_16998_ _16029_/Y _24390_/Q _24737_/Q _17032_/A VGND VGND VPWR VPWR _17000_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18737_ _18736_/X VGND VGND VPWR VPWR _24150_/D sky130_fd_sc_hd__inv_2
X_15949_ _15931_/X VGND VGND VPWR VPWR _15949_/X sky130_fd_sc_hd__buf_2
XFILLER_243_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18668_ _18663_/X _18668_/B _18668_/C _18668_/D VGND VGND VPWR VPWR _18668_/X sky130_fd_sc_hd__or4_4
XFILLER_236_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17619_ _17511_/Y _17615_/X VGND VGND VPWR VPWR _17619_/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12218__B2 _22150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_118_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_237_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_18599_ _24137_/Q VGND VGND VPWR VPWR _18791_/A sky130_fd_sc_hd__buf_2
XANTENNA__18692__A _24142_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20630_ _20630_/A _17386_/X VGND VGND VPWR VPWR _20630_/Y sky130_fd_sc_hd__nand2_4
X_20561_ _20560_/X VGND VGND VPWR VPWR _23940_/D sky130_fd_sc_hd__inv_2
X_22300_ _24041_/Q VGND VGND VPWR VPWR _22300_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20492_ _20517_/A _15432_/A _20490_/X _15432_/A _20491_/X VGND VGND VPWR VPWR _20492_/X
+ sky130_fd_sc_hd__a32o_4
X_23280_ _23280_/A _23280_/B VGND VGND VPWR VPWR _23287_/C sky130_fd_sc_hd__and2_4
XANTENNA__24396__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22231_ _22231_/A VGND VGND VPWR VPWR _22231_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22453__A2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24325__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22162_ _23176_/A _22162_/B _22161_/X VGND VGND VPWR VPWR _22195_/A sky130_fd_sc_hd__and3_4
XFILLER_117_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21113_ _22429_/A VGND VGND VPWR VPWR _21859_/A sky130_fd_sc_hd__inv_2
XFILLER_160_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22093_ _14986_/A _22420_/B _21339_/X VGND VGND VPWR VPWR _22093_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_8_56_0_HCLK clkbuf_7_28_0_HCLK/X VGND VGND VPWR VPWR _23398_/CLK sky130_fd_sc_hd__clkbuf_1
X_21044_ _12592_/A _15649_/Y _21042_/X _21043_/X VGND VGND VPWR VPWR _21045_/A sky130_fd_sc_hd__a211o_4
XFILLER_87_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17771__A _23320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24956__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24803_ _24874_/CLK _15877_/X HRESETn VGND VGND VPWR VPWR _22861_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16840__B1 _16518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21293__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23960__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22995_ _22995_/A VGND VGND VPWR VPWR _23209_/A sky130_fd_sc_hd__buf_2
XFILLER_216_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24734_ _24737_/CLK _16028_/X HRESETn VGND VGND VPWR VPWR _24734_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_243_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21946_ _21942_/X _21945_/X _17725_/A VGND VGND VPWR VPWR _21946_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24665_ _24667_/CLK _16218_/X HRESETn VGND VGND VPWR VPWR _22883_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21877_ _22435_/A _21875_/X _21439_/X _21876_/X VGND VGND VPWR VPWR _21877_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22126__D1 _22125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _23458_/CLK _23616_/D VGND VGND VPWR VPWR _23616_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ _20919_/A VGND VGND VPWR VPWR _20828_/X sky130_fd_sc_hd__buf_2
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24596_ _24594_/CLK _24596_/D HRESETn VGND VGND VPWR VPWR _16404_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23547_ _23534_/CLK _19987_/X VGND VGND VPWR VPWR _19986_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20759_ _13107_/C VGND VGND VPWR VPWR _20759_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14635__A _18090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13300_/A _13297_/X _13299_/X VGND VGND VPWR VPWR _13300_/X sky130_fd_sc_hd__and3_4
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ _14280_/A _14285_/A _14283_/A _14283_/B VGND VGND VPWR VPWR _14281_/A sky130_fd_sc_hd__or4_4
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23478_ _23487_/CLK _23478_/D VGND VGND VPWR VPWR _23478_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13231_ _13397_/A VGND VGND VPWR VPWR _13231_/X sky130_fd_sc_hd__buf_2
X_25217_ _25224_/CLK _14144_/X HRESETn VGND VGND VPWR VPWR _14089_/C sky130_fd_sc_hd__dfrtp_4
X_22429_ _22429_/A VGND VGND VPWR VPWR _22429_/X sky130_fd_sc_hd__buf_2
XANTENNA__24066__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13162_ _13394_/A VGND VGND VPWR VPWR _13162_/X sky130_fd_sc_hd__buf_2
X_25148_ _24326_/CLK _14387_/X HRESETn VGND VGND VPWR VPWR _25148_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12113_ _24101_/Q _24102_/Q VGND VGND VPWR VPWR _12120_/A sky130_fd_sc_hd__and2_4
XANTENNA__15466__A _14380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13093_ _13092_/X VGND VGND VPWR VPWR _25339_/D sky130_fd_sc_hd__inv_2
X_17970_ _18027_/A _23769_/Q VGND VGND VPWR VPWR _17973_/B sky130_fd_sc_hd__or2_4
X_25079_ _25081_/CLK _25079_/D HRESETn VGND VGND VPWR VPWR _14606_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14370__A _14096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12044_ _12043_/Y VGND VGND VPWR VPWR _17436_/C sky130_fd_sc_hd__buf_2
X_16921_ _16921_/A VGND VGND VPWR VPWR _16921_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19640_ _13375_/B VGND VGND VPWR VPWR _19640_/Y sky130_fd_sc_hd__inv_2
X_16852_ _16852_/A VGND VGND VPWR VPWR _16852_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15803_ _15792_/X VGND VGND VPWR VPWR _15803_/X sky130_fd_sc_hd__buf_2
X_16783_ _18965_/A VGND VGND VPWR VPWR _16783_/X sky130_fd_sc_hd__buf_2
X_19571_ _19570_/X VGND VGND VPWR VPWR _19572_/A sky130_fd_sc_hd__inv_2
X_13995_ _13995_/A _13995_/B _25234_/Q _13995_/D VGND VGND VPWR VPWR _13995_/X sky130_fd_sc_hd__and4_4
XFILLER_46_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15734_ _12547_/Y _15731_/X _11721_/X _15731_/X VGND VGND VPWR VPWR _15734_/X sky130_fd_sc_hd__a2bb2o_4
X_18522_ _18522_/A VGND VGND VPWR VPWR _18522_/Y sky130_fd_sc_hd__inv_2
X_12946_ _12945_/X VGND VGND VPWR VPWR _25376_/D sky130_fd_sc_hd__inv_2
XFILLER_46_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15665_ _21587_/A VGND VGND VPWR VPWR _15665_/X sky130_fd_sc_hd__buf_2
X_18453_ _18425_/X _18453_/B VGND VGND VPWR VPWR _18745_/C sky130_fd_sc_hd__or2_4
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12877_ _12879_/B VGND VGND VPWR VPWR _12878_/B sky130_fd_sc_hd__inv_2
XANTENNA__15937__A2 _15928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20930__A2 _20846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _21968_/A _14610_/A _14615_/A _13623_/X VGND VGND VPWR VPWR _14616_/X sky130_fd_sc_hd__o22a_4
X_17404_ _17384_/X _17398_/X _23992_/Q _21002_/B _17401_/X VGND VGND VPWR VPWR _24338_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _11826_/A _24236_/Q _11826_/Y _22541_/A VGND VGND VPWR VPWR _11835_/B sky130_fd_sc_hd__o22a_4
X_18384_ _18383_/Y _18379_/X _24193_/Q _18379_/X VGND VGND VPWR VPWR _18384_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21650__B _21649_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15596_ _15576_/A VGND VGND VPWR VPWR _15596_/X sky130_fd_sc_hd__buf_2
XFILLER_187_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12253__A2_N _24751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24836__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17335_ _17335_/A VGND VGND VPWR VPWR _17335_/Y sky130_fd_sc_hd__inv_2
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14547_/A VGND VGND VPWR VPWR _14563_/A sky130_fd_sc_hd__buf_2
XFILLER_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11759_ _25527_/Q VGND VGND VPWR VPWR _11759_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17266_ _17191_/Y _17231_/X _17265_/X VGND VGND VPWR VPWR _17266_/X sky130_fd_sc_hd__or3_4
XANTENNA__21891__B1 _22205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14478_ HWDATA[1] VGND VGND VPWR VPWR _18951_/A sky130_fd_sc_hd__buf_2
XFILLER_147_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16217_ _22883_/A VGND VGND VPWR VPWR _16217_/Y sky130_fd_sc_hd__inv_2
X_19005_ HWDATA[7] VGND VGND VPWR VPWR _19006_/A sky130_fd_sc_hd__buf_2
X_13429_ _13397_/A _13427_/X _13429_/C VGND VGND VPWR VPWR _13429_/X sky130_fd_sc_hd__and3_4
X_17197_ _24614_/Q _24343_/Q _16355_/Y _17242_/B VGND VGND VPWR VPWR _17198_/D sky130_fd_sc_hd__o22a_4
XFILLER_174_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16148_ _16147_/Y _16142_/X _16055_/X _16142_/X VGND VGND VPWR VPWR _24688_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16079_ _16077_/A _15670_/X VGND VGND VPWR VPWR _16079_/X sky130_fd_sc_hd__or2_4
XFILLER_103_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19907_ _23575_/Q VGND VGND VPWR VPWR _19907_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19838_ _22209_/B _19835_/X _19810_/X _19835_/X VGND VGND VPWR VPWR _23601_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19769_ _19764_/A VGND VGND VPWR VPWR _19769_/X sky130_fd_sc_hd__buf_2
X_21800_ _21472_/A _21800_/B _21799_/X VGND VGND VPWR VPWR _21800_/X sky130_fd_sc_hd__and3_4
X_22780_ _22774_/X _22777_/Y _22493_/X _22779_/X VGND VGND VPWR VPWR _22780_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16000__A _24744_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21174__A2 _15662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21731_ _13496_/Y _21570_/X _12024_/Y _21571_/X VGND VGND VPWR VPWR _21731_/X sky130_fd_sc_hd__o22a_4
XFILLER_224_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24450_ _24463_/CLK _24450_/D HRESETn VGND VGND VPWR VPWR _15022_/A sky130_fd_sc_hd__dfrtp_4
X_21662_ _21662_/A _21662_/B VGND VGND VPWR VPWR _21662_/X sky130_fd_sc_hd__or2_4
XFILLER_240_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24577__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23401_ _25272_/CLK _20371_/X VGND VGND VPWR VPWR _23401_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20613_ _13956_/A _20613_/B _15424_/C VGND VGND VPWR VPWR _23966_/D sky130_fd_sc_hd__and3_4
X_24381_ _24725_/CLK _24381_/D HRESETn VGND VGND VPWR VPWR _24381_/Q sky130_fd_sc_hd__dfrtp_4
X_21593_ _21593_/A _11704_/A VGND VGND VPWR VPWR _21593_/X sky130_fd_sc_hd__and2_4
XFILLER_177_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14455__A _14455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22674__A2 _22821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24506__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23332_ _22708_/A _23329_/X _23331_/X VGND VGND VPWR VPWR _23337_/C sky130_fd_sc_hd__and3_4
X_20544_ _20544_/A _18888_/A VGND VGND VPWR VPWR _20544_/X sky130_fd_sc_hd__and2_4
XANTENNA__17550__B2 _24113_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23263_ _24475_/Q _23263_/B _23263_/C VGND VGND VPWR VPWR _23263_/X sky130_fd_sc_hd__and3_4
XANTENNA__22426__A2 _22419_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20475_ _20502_/B VGND VGND VPWR VPWR _20515_/B sky130_fd_sc_hd__buf_2
X_25002_ _24953_/CLK _25002_/D HRESETn VGND VGND VPWR VPWR _15082_/A sky130_fd_sc_hd__dfrtp_4
X_22214_ _22209_/A _22214_/B VGND VGND VPWR VPWR _22214_/X sky130_fd_sc_hd__or2_4
X_23194_ _22552_/X _23193_/X _23050_/X _24110_/Q _22555_/X VGND VGND VPWR VPWR _23194_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20192__A _20180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22145_ _24617_/Q _22145_/B VGND VGND VPWR VPWR _22145_/X sky130_fd_sc_hd__or2_4
XFILLER_121_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22076_ _22387_/A _20038_/Y VGND VGND VPWR VPWR _22077_/C sky130_fd_sc_hd__or2_4
XFILLER_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25365__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21027_ _21027_/A _22423_/A VGND VGND VPWR VPWR _21027_/X sky130_fd_sc_hd__or2_4
XFILLER_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12800_ _12800_/A VGND VGND VPWR VPWR _12800_/Y sky130_fd_sc_hd__inv_2
X_13780_ _13779_/X VGND VGND VPWR VPWR _13780_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22978_ _22486_/X _22977_/X _22489_/X _24737_/Q _22865_/X VGND VGND VPWR VPWR _22979_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_216_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12731_ _12830_/A _24796_/Q _12830_/A _24796_/Q VGND VGND VPWR VPWR _12731_/X sky130_fd_sc_hd__a2bb2o_4
X_24717_ _24639_/CLK _16072_/X HRESETn VGND VGND VPWR VPWR _24717_/Q sky130_fd_sc_hd__dfrtp_4
X_21929_ _22343_/A _20336_/Y VGND VGND VPWR VPWR _21933_/B sky130_fd_sc_hd__or2_4
XFILLER_203_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15450_ _13903_/A _15444_/X _15441_/X _13935_/B _15447_/X VGND VGND VPWR VPWR _24963_/D
+ sky130_fd_sc_hd__a32o_4
X_12662_ _12555_/Y _12662_/B VGND VGND VPWR VPWR _12675_/A sky130_fd_sc_hd__or2_4
X_24648_ _24592_/CLK _16264_/X HRESETn VGND VGND VPWR VPWR _21335_/A sky130_fd_sc_hd__dfrtp_4
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_101_0_HCLK clkbuf_6_50_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_202_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14394_/Y _14398_/X _14400_/X _14398_/X VGND VGND VPWR VPWR _25145_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23311__B1 _24886_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21546__A2_N _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14987__A2_N _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15380_/X VGND VGND VPWR VPWR _24988_/D sky130_fd_sc_hd__inv_2
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12592_/Y VGND VGND VPWR VPWR _12681_/A sky130_fd_sc_hd__buf_2
X_24579_ _24678_/CLK _24579_/D HRESETn VGND VGND VPWR VPWR _24579_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24247__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ _17120_/A _17120_/B VGND VGND VPWR VPWR _17121_/C sky130_fd_sc_hd__or2_4
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _14329_/C _14332_/B VGND VGND VPWR VPWR _14337_/A sky130_fd_sc_hd__or2_4
XFILLER_128_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_5_21_0_HCLK_A clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17051_ _17070_/A _17051_/B _17051_/C VGND VGND VPWR VPWR _24404_/D sky130_fd_sc_hd__and3_4
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _14261_/Y _14259_/X _14262_/X _14259_/X VGND VGND VPWR VPWR _14263_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_167_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16002_ _16000_/Y _15998_/X _16001_/X _15998_/X VGND VGND VPWR VPWR _16002_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13214_ _13260_/A _13214_/B VGND VGND VPWR VPWR _13214_/X sky130_fd_sc_hd__or2_4
XFILLER_136_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14194_ _25207_/Q VGND VGND VPWR VPWR _20517_/A sky130_fd_sc_hd__inv_2
XANTENNA__23090__A2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13145_ _13397_/A VGND VGND VPWR VPWR _13172_/A sky130_fd_sc_hd__buf_2
XFILLER_124_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13076_ _12981_/C _13079_/B _13019_/X VGND VGND VPWR VPWR _13076_/Y sky130_fd_sc_hd__a21oi_4
X_17953_ _17942_/A _17951_/X _17952_/X VGND VGND VPWR VPWR _17953_/X sky130_fd_sc_hd__and3_4
XFILLER_239_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12027_ _12014_/Y VGND VGND VPWR VPWR _12027_/X sky130_fd_sc_hd__buf_2
X_16904_ _24266_/Q VGND VGND VPWR VPWR _16904_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25035__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17884_ _16917_/Y _17880_/X VGND VGND VPWR VPWR _17884_/Y sky130_fd_sc_hd__nand2_4
X_19623_ _21193_/B _19616_/X _19475_/X _19598_/Y VGND VGND VPWR VPWR _19623_/X sky130_fd_sc_hd__a2bb2o_4
X_16835_ _16833_/Y _16834_/X _15748_/X _16834_/X VGND VGND VPWR VPWR _24425_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13444__A _13254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19554_ _23696_/Q VGND VGND VPWR VPWR _22029_/B sky130_fd_sc_hd__inv_2
X_13978_ _13978_/A VGND VGND VPWR VPWR _13978_/X sky130_fd_sc_hd__buf_2
X_16766_ _16766_/A VGND VGND VPWR VPWR _16766_/X sky130_fd_sc_hd__buf_2
XFILLER_202_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18505_ _18505_/A _18493_/B VGND VGND VPWR VPWR _18506_/C sky130_fd_sc_hd__or2_4
XFILLER_222_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12929_ _12833_/X _12958_/B VGND VGND VPWR VPWR _12929_/X sky130_fd_sc_hd__or2_4
X_15717_ _15713_/X VGND VGND VPWR VPWR _15717_/X sky130_fd_sc_hd__buf_2
XFILLER_206_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16697_ _16692_/A VGND VGND VPWR VPWR _16697_/X sky130_fd_sc_hd__buf_2
X_19485_ _22258_/B _19482_/X _11906_/X _19482_/X VGND VGND VPWR VPWR _23721_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18436_ _16219_/Y _24175_/Q _22996_/A _18468_/A VGND VGND VPWR VPWR _18438_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15648_ _21138_/A _17436_/C _16446_/D _12160_/C VGND VGND VPWR VPWR _15648_/X sky130_fd_sc_hd__or4_4
XFILLER_210_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24670__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15579_ _15578_/Y _15576_/X _11695_/X _15576_/X VGND VGND VPWR VPWR _15579_/X sky130_fd_sc_hd__a2bb2o_4
X_18367_ _18354_/A _18353_/X VGND VGND VPWR VPWR _18367_/X sky130_fd_sc_hd__or2_4
XFILLER_187_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17318_ _17200_/Y _17318_/B VGND VGND VPWR VPWR _17319_/B sky130_fd_sc_hd__or2_4
X_18298_ _18292_/X _18298_/B VGND VGND VPWR VPWR _18298_/X sky130_fd_sc_hd__or2_4
XANTENNA__14346__A1 MSO_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17249_ _17329_/A _17248_/Y _17249_/C _17249_/D VGND VGND VPWR VPWR _17249_/X sky130_fd_sc_hd__or4_4
XFILLER_135_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14346__B2 _14340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22408__A2 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20260_ _21266_/B _20255_/X _20133_/X _20243_/A VGND VGND VPWR VPWR _20260_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20191_ _20191_/A VGND VGND VPWR VPWR _21611_/B sky130_fd_sc_hd__inv_2
XANTENNA__16638__A3 _15702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15809__A1_N _12329_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23950_ _25211_/CLK _20600_/Y HRESETn VGND VGND VPWR VPWR _23950_/Q sky130_fd_sc_hd__dfrtp_4
X_22901_ _22901_/A _22901_/B VGND VGND VPWR VPWR _22901_/X sky130_fd_sc_hd__or2_4
XFILLER_243_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23881_ _23844_/CLK _19031_/X VGND VGND VPWR VPWR _18002_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13609__B1 _18060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22832_ _21592_/A VGND VGND VPWR VPWR _22832_/X sky130_fd_sc_hd__buf_2
XFILLER_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22667__A _22667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24758__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22763_ _12801_/X _22761_/X _22762_/X VGND VGND VPWR VPWR _22763_/X sky130_fd_sc_hd__o21a_4
X_24502_ _25021_/CLK _24502_/D HRESETn VGND VGND VPWR VPWR _24502_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21714_ _21289_/X _21700_/X _21703_/X _21710_/X _21713_/X VGND VGND VPWR VPWR _21714_/X
+ sky130_fd_sc_hd__o41a_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25482_ _25158_/CLK _25482_/D HRESETn VGND VGND VPWR VPWR _25482_/Q sky130_fd_sc_hd__dfrtp_4
X_22694_ _22694_/A VGND VGND VPWR VPWR _22726_/A sky130_fd_sc_hd__inv_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24433_ _24462_/CLK _16817_/X HRESETn VGND VGND VPWR VPWR _14922_/A sky130_fd_sc_hd__dfrtp_4
X_21645_ _21960_/B VGND VGND VPWR VPWR _22397_/B sky130_fd_sc_hd__buf_2
XANTENNA__13801__B _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22647__A2 _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24364_ _24634_/CLK _24364_/D HRESETn VGND VGND VPWR VPWR _17298_/A sky130_fd_sc_hd__dfrtp_4
X_21576_ _21569_/X _21572_/X _21573_/X _21575_/X VGND VGND VPWR VPWR _21576_/X sky130_fd_sc_hd__o22a_4
X_23315_ _23315_/A VGND VGND VPWR VPWR _23315_/Y sky130_fd_sc_hd__inv_2
X_20527_ _20480_/X _20495_/X _20504_/A _20519_/A VGND VGND VPWR VPWR _20527_/X sky130_fd_sc_hd__or4_4
XFILLER_126_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15534__B1 HADDR[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24295_ _24305_/CLK _24295_/D HRESETn VGND VGND VPWR VPWR _24295_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23246_ _23182_/A _23237_/Y _23246_/C _23246_/D VGND VGND VPWR VPWR _23246_/X sky130_fd_sc_hd__or4_4
X_20458_ _20430_/A _20456_/X _20464_/C _20457_/X VGND VGND VPWR VPWR _20458_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25546__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23177_ _24606_/Q _23177_/B VGND VGND VPWR VPWR _23181_/B sky130_fd_sc_hd__or2_4
X_20389_ _20389_/A VGND VGND VPWR VPWR _20389_/X sky130_fd_sc_hd__buf_2
XFILLER_97_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22128_ _21319_/X VGND VGND VPWR VPWR _22140_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_26_0_HCLK clkbuf_7_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_26_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14950_ _25031_/Q VGND VGND VPWR VPWR _14951_/A sky130_fd_sc_hd__inv_2
X_22059_ _21896_/X _22059_/B _22058_/X VGND VGND VPWR VPWR _22059_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_89_0_HCLK clkbuf_7_89_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_89_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13901_ _13907_/A _13887_/Y _13897_/X _13907_/C _13900_/X VGND VGND VPWR VPWR _13901_/X
+ sky130_fd_sc_hd__a32o_4
X_14881_ _14880_/Y VGND VGND VPWR VPWR _15249_/A sky130_fd_sc_hd__buf_2
XFILLER_48_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13264__A _13289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13832_ _13832_/A VGND VGND VPWR VPWR _13832_/X sky130_fd_sc_hd__buf_2
X_16620_ _16619_/Y _16541_/X _16361_/X _16541_/X VGND VGND VPWR VPWR _16620_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16586__A1_N _16584_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22577__A _22539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22335__A1 _21345_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24499__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16551_ _16550_/Y _16548_/X _16464_/X _16548_/X VGND VGND VPWR VPWR _16551_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21481__A _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13763_ _13807_/C VGND VGND VPWR VPWR _13763_/X sky130_fd_sc_hd__buf_2
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24428__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17211__B1 _24633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12714_ _12569_/Y _12690_/X _12711_/Y _12641_/X VGND VGND VPWR VPWR _12714_/X sky130_fd_sc_hd__a211o_4
X_15502_ _15501_/Y _15499_/X HADDR[16] _15499_/X VGND VGND VPWR VPWR _24941_/D sky130_fd_sc_hd__a2bb2o_4
X_16482_ _16470_/A VGND VGND VPWR VPWR _16482_/X sky130_fd_sc_hd__buf_2
X_19270_ _23795_/Q VGND VGND VPWR VPWR _21249_/B sky130_fd_sc_hd__inv_2
X_13694_ _13666_/Y VGND VGND VPWR VPWR _13694_/X sky130_fd_sc_hd__buf_2
XFILLER_16_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15433_ _15436_/B VGND VGND VPWR VPWR _15433_/X sky130_fd_sc_hd__buf_2
X_18221_ _18125_/A _23843_/Q VGND VGND VPWR VPWR _18223_/B sky130_fd_sc_hd__or2_4
XANTENNA__22099__B1 _21339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12645_ _12648_/A _12645_/B _12645_/C VGND VGND VPWR VPWR _25425_/D sky130_fd_sc_hd__and3_4
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24081__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ _15361_/A _15367_/B VGND VGND VPWR VPWR _15364_/Y sky130_fd_sc_hd__nand2_4
X_18152_ _18085_/A _18152_/B _18151_/X VGND VGND VPWR VPWR _18156_/B sky130_fd_sc_hd__and3_4
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12576_ _12567_/A _12574_/Y _12655_/A _24875_/Q VGND VGND VPWR VPWR _12577_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20825__A _20846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17514__A1 _25527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24010__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14315_ _25169_/Q _12151_/X _14314_/X VGND VGND VPWR VPWR _14315_/X sky130_fd_sc_hd__a21o_4
X_17103_ _17103_/A _17103_/B VGND VGND VPWR VPWR _17103_/X sky130_fd_sc_hd__or2_4
XFILLER_8_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18083_ _18118_/A _18083_/B VGND VGND VPWR VPWR _18083_/X sky130_fd_sc_hd__or2_4
XANTENNA__15525__B1 HADDR[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15295_ _15295_/A VGND VGND VPWR VPWR _15390_/A sky130_fd_sc_hd__inv_2
XFILLER_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17034_ _17034_/A VGND VGND VPWR VPWR _17043_/B sky130_fd_sc_hd__inv_2
X_14246_ _14246_/A _14212_/B VGND VGND VPWR VPWR _14247_/A sky130_fd_sc_hd__nor2_4
XFILLER_183_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15638__B _22829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14542__B HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22271__B1 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14177_ _14177_/A _14177_/B VGND VGND VPWR VPWR _14365_/D sky130_fd_sc_hd__or2_4
XANTENNA__25216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13128_ _13128_/A _20688_/B VGND VGND VPWR VPWR _13128_/X sky130_fd_sc_hd__and2_4
X_18985_ _18985_/A VGND VGND VPWR VPWR _18985_/X sky130_fd_sc_hd__buf_2
XFILLER_112_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13059_ _13059_/A _12984_/X VGND VGND VPWR VPWR _13059_/X sky130_fd_sc_hd__or2_4
X_17936_ _17940_/A _23778_/Q VGND VGND VPWR VPWR _17938_/B sky130_fd_sc_hd__or2_4
XFILLER_112_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17867_ _17849_/X _17862_/B _17793_/A _17864_/B VGND VGND VPWR VPWR _17867_/X sky130_fd_sc_hd__a211o_4
XFILLER_213_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17176__A2_N _17249_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19606_ _19606_/A VGND VGND VPWR VPWR _19606_/X sky130_fd_sc_hd__buf_2
X_16818_ _14908_/Y _16816_/X HWDATA[18] _16816_/X VGND VGND VPWR VPWR _24432_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17798_ _17800_/B VGND VGND VPWR VPWR _17798_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24851__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19537_ _19536_/Y _19531_/X _19377_/X _19531_/X VGND VGND VPWR VPWR _19537_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16749_ _16730_/A VGND VGND VPWR VPWR _16749_/X sky130_fd_sc_hd__buf_2
XANTENNA__20337__B1 _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16485__A _16485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24169__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19468_ _21813_/B _19463_/X _11920_/X _19463_/X VGND VGND VPWR VPWR _23726_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18419_ _16244_/A _24167_/Q _16244_/Y _18567_/A VGND VGND VPWR VPWR _18424_/B sky130_fd_sc_hd__o22a_4
XFILLER_194_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19399_ _19398_/Y _19396_/X _19351_/X _19396_/X VGND VGND VPWR VPWR _19399_/X sky130_fd_sc_hd__a2bb2o_4
X_21430_ _22298_/A _21430_/B VGND VGND VPWR VPWR _21430_/Y sky130_fd_sc_hd__nand2_4
XFILLER_147_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21837__B1 _15465_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21361_ _13483_/A _17436_/B _21357_/X _21568_/A _21360_/X VGND VGND VPWR VPWR _21361_/X
+ sky130_fd_sc_hd__o32a_4
X_23100_ _23077_/X _23081_/X _23092_/X _23099_/X VGND VGND VPWR VPWR HRDATA[24] sky130_fd_sc_hd__or4_4
X_20312_ _20306_/X _19573_/X _13826_/A _22266_/A _20310_/X VGND VGND VPWR VPWR _20312_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24080_ _24080_/CLK _20501_/X HRESETn VGND VGND VPWR VPWR _20479_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_162_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21292_ _21598_/A VGND VGND VPWR VPWR _21292_/X sky130_fd_sc_hd__buf_2
X_23031_ _22761_/X _23029_/X _22691_/X _23030_/X VGND VGND VPWR VPWR _23031_/X sky130_fd_sc_hd__o22a_4
X_20243_ _20243_/A VGND VGND VPWR VPWR _20243_/X sky130_fd_sc_hd__buf_2
XFILLER_115_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15819__B2 _15786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20174_ _21405_/B _20171_/X _20109_/X _20171_/X VGND VGND VPWR VPWR _23476_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15564__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24982_ _24980_/CLK _15403_/X HRESETn VGND VGND VPWR VPWR _15153_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24939__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23933_ _23951_/CLK _20983_/X HRESETn VGND VGND VPWR VPWR _20987_/B sky130_fd_sc_hd__dfstp_4
XFILLER_123_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17441__B1 _17440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23864_ _23610_/CLK _23864_/D VGND VGND VPWR VPWR _23864_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14255__B1 _13785_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24592__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22815_ _22132_/B VGND VGND VPWR VPWR _22817_/B sky130_fd_sc_hd__buf_2
XFILLER_44_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23795_ _23859_/CLK _19271_/X VGND VGND VPWR VPWR _23795_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16395__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24521__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25534_ _25533_/CLK _11736_/X HRESETn VGND VGND VPWR VPWR _25534_/Q sky130_fd_sc_hd__dfrtp_4
X_22746_ _21109_/A _22745_/X _22296_/X _24870_/Q _21098_/A VGND VGND VPWR VPWR _22747_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25465_ _25466_/CLK _25465_/D HRESETn VGND VGND VPWR VPWR _12163_/A sky130_fd_sc_hd__dfrtp_4
X_22677_ _16232_/Y _22454_/X _16413_/Y _22450_/X VGND VGND VPWR VPWR _22678_/B sky130_fd_sc_hd__o22a_4
X_12430_ _12201_/Y _12428_/X _12429_/Y VGND VGND VPWR VPWR _12430_/X sky130_fd_sc_hd__o21a_4
X_24416_ _24477_/CLK _16850_/X HRESETn VGND VGND VPWR VPWR _14932_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21628_ _22381_/A _19846_/Y VGND VGND VPWR VPWR _21631_/B sky130_fd_sc_hd__or2_4
X_25396_ _25397_/CLK _25396_/D HRESETn VGND VGND VPWR VPWR _12828_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12361_ _12360_/Y _24823_/Q _12982_/A _12332_/Y VGND VGND VPWR VPWR _12368_/A sky130_fd_sc_hd__a2bb2o_4
X_24347_ _24667_/CLK _24347_/D HRESETn VGND VGND VPWR VPWR _24347_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15739__A HWDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15507__B1 HADDR[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21559_ _21559_/A VGND VGND VPWR VPWR _21559_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14100_ _14115_/A VGND VGND VPWR VPWR _14100_/X sky130_fd_sc_hd__buf_2
XFILLER_138_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15080_ _15366_/A _16404_/A _15078_/Y _16404_/A VGND VGND VPWR VPWR _15089_/A sky130_fd_sc_hd__a2bb2o_4
X_12292_ _12291_/X _24836_/Q _12291_/A _24836_/Q VGND VGND VPWR VPWR _12301_/A sky130_fd_sc_hd__a2bb2o_4
X_24278_ _24278_/CLK _17820_/Y HRESETn VGND VGND VPWR VPWR _24278_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25380__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14031_ _25242_/Q _13995_/B _25234_/Q _13994_/A VGND VGND VPWR VPWR _14032_/A sky130_fd_sc_hd__or4_4
X_23229_ _12264_/Y _21532_/X _24286_/Q _22493_/X VGND VGND VPWR VPWR _23229_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13259__A _13334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18770_ _18689_/Y _18770_/B VGND VGND VPWR VPWR _18771_/C sky130_fd_sc_hd__or2_4
X_15982_ _21745_/B VGND VGND VPWR VPWR _23138_/A sky130_fd_sc_hd__buf_2
XANTENNA__22556__A1 _22552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22556__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17721_ _18280_/C _21473_/A _18280_/C _21473_/A VGND VGND VPWR VPWR _17736_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14933_ _25010_/Q _14932_/A _15273_/A _14932_/Y VGND VGND VPWR VPWR _14934_/D sky130_fd_sc_hd__o22a_4
XANTENNA__24609__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17432__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17652_ _17647_/A _17648_/B _17652_/C VGND VGND VPWR VPWR _17652_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_113_0_HCLK clkbuf_7_56_0_HCLK/X VGND VGND VPWR VPWR _24795_/CLK sky130_fd_sc_hd__clkbuf_1
X_14864_ _14859_/A VGND VGND VPWR VPWR _14864_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16603_ _24522_/Q VGND VGND VPWR VPWR _16603_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_176_0_HCLK clkbuf_7_88_0_HCLK/X VGND VGND VPWR VPWR _25158_/CLK sky130_fd_sc_hd__clkbuf_1
X_13815_ _13533_/Y _13813_/X _11743_/X _13813_/X VGND VGND VPWR VPWR _13815_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14795_ _25047_/Q _14795_/B _14810_/A VGND VGND VPWR VPWR _14796_/B sky130_fd_sc_hd__or3_4
X_17583_ _17571_/X _17628_/B VGND VGND VPWR VPWR _17583_/X sky130_fd_sc_hd__or2_4
XANTENNA__15994__B1 _15554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14818__A _14817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24262__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19322_ _19327_/A VGND VGND VPWR VPWR _19322_/X sky130_fd_sc_hd__buf_2
XFILLER_189_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13746_ _13739_/Y _13745_/X VGND VGND VPWR VPWR _13746_/X sky130_fd_sc_hd__or2_4
X_16534_ _16534_/A VGND VGND VPWR VPWR _16534_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15640__C _15640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19253_ _19253_/A VGND VGND VPWR VPWR _19253_/Y sky130_fd_sc_hd__inv_2
X_13677_ _11826_/Y _13677_/B VGND VGND VPWR VPWR _13678_/B sky130_fd_sc_hd__or2_4
X_16465_ _16463_/Y _16461_/X _16464_/X _16461_/X VGND VGND VPWR VPWR _16465_/X sky130_fd_sc_hd__a2bb2o_4
X_18204_ _17984_/X _18202_/X _18203_/X VGND VGND VPWR VPWR _18204_/X sky130_fd_sc_hd__and3_4
X_12628_ _12594_/Y _12626_/X _12627_/X _12623_/B VGND VGND VPWR VPWR _12628_/X sky130_fd_sc_hd__a211o_4
X_15416_ _15382_/X VGND VGND VPWR VPWR _15417_/B sky130_fd_sc_hd__inv_2
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16396_ _15142_/Y _16393_/X _16395_/X _16393_/X VGND VGND VPWR VPWR _16396_/X sky130_fd_sc_hd__a2bb2o_4
X_19184_ _19002_/B _19026_/C _19026_/D _19341_/A VGND VGND VPWR VPWR _19184_/X sky130_fd_sc_hd__and4_4
XFILLER_176_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12162__A1_N SSn_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15347_ _15347_/A _15347_/B VGND VGND VPWR VPWR _15347_/X sky130_fd_sc_hd__or2_4
X_18135_ _18103_/A _18135_/B VGND VGND VPWR VPWR _18137_/B sky130_fd_sc_hd__or2_4
XANTENNA__15649__A _15648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12559_ _12558_/Y _24868_/Q _12558_/Y _24868_/Q VGND VGND VPWR VPWR _12566_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_156_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15278_ _15272_/A _15243_/B VGND VGND VPWR VPWR _15278_/Y sky130_fd_sc_hd__nand2_4
X_18066_ _18103_/A _19350_/A VGND VGND VPWR VPWR _18068_/B sky130_fd_sc_hd__or2_4
XFILLER_171_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14229_ _25194_/Q VGND VGND VPWR VPWR _14229_/Y sky130_fd_sc_hd__inv_2
X_17017_ _17333_/A VGND VGND VPWR VPWR _17087_/A sky130_fd_sc_hd__buf_2
XFILLER_171_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17864__A _16915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25050__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18999__B1 _18998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18968_ _23901_/Q VGND VGND VPWR VPWR _18968_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17919_ _17918_/Y _15905_/X _17917_/B VGND VGND VPWR VPWR _17919_/X sky130_fd_sc_hd__a21o_4
XFILLER_224_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18899_ _11948_/A _11938_/B _11935_/X VGND VGND VPWR VPWR _18899_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_239_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_72_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_72_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17423__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20930_ _16659_/Y _20846_/A _20855_/X _20929_/X VGND VGND VPWR VPWR _20931_/A sky130_fd_sc_hd__o22a_4
XFILLER_94_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20861_ _24043_/Q VGND VGND VPWR VPWR _20862_/C sky130_fd_sc_hd__inv_2
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23972__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22600_ _22279_/A _22599_/X _21312_/X _24727_/Q _21708_/X VGND VGND VPWR VPWR _22600_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12799__B1 _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23580_ _24297_/CLK _23580_/D VGND VGND VPWR VPWR _19893_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20792_ _20791_/X VGND VGND VPWR VPWR _20792_/Y sky130_fd_sc_hd__inv_2
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18923__B1 _16783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22531_ _23301_/B VGND VGND VPWR VPWR _22532_/B sky130_fd_sc_hd__buf_2
XANTENNA__18427__A2_N _18467_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25250_ _25230_/CLK _13859_/X HRESETn VGND VGND VPWR VPWR _25250_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23985__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22462_ _12092_/Y _12058_/B _12000_/Y _13456_/X VGND VGND VPWR VPWR _22462_/X sky130_fd_sc_hd__o22a_4
X_24201_ _24257_/CLK _24201_/D HRESETn VGND VGND VPWR VPWR _18350_/A sky130_fd_sc_hd__dfrtp_4
X_21413_ _14681_/A _21411_/X _21412_/X VGND VGND VPWR VPWR _21413_/X sky130_fd_sc_hd__and3_4
X_25181_ _25171_/CLK _14287_/X HRESETn VGND VGND VPWR VPWR _25181_/Q sky130_fd_sc_hd__dfrtp_4
X_22393_ _22393_/A _22392_/Y VGND VGND VPWR VPWR _22393_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14463__A _14468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24132_ _24133_/CLK _24132_/D HRESETn VGND VGND VPWR VPWR _24132_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21344_ _21343_/X VGND VGND VPWR VPWR _21720_/A sky130_fd_sc_hd__buf_2
XFILLER_108_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16162__B1 _15901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23027__A2 _22718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13079__A _13085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24063_ _24060_/CLK _20951_/X HRESETn VGND VGND VPWR VPWR _20953_/B sky130_fd_sc_hd__dfrtp_4
X_21275_ _21258_/X _21273_/X _21274_/X VGND VGND VPWR VPWR _21275_/X sky130_fd_sc_hd__a21o_4
XFILLER_190_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23014_ _24738_/Q _21061_/X _21062_/X _23013_/X VGND VGND VPWR VPWR _23014_/X sky130_fd_sc_hd__a211o_4
X_20226_ _20226_/A VGND VGND VPWR VPWR _20226_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13807__A _13807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20157_ _13753_/X _13737_/X _20157_/C _20157_/D VGND VGND VPWR VPWR _20158_/A sky130_fd_sc_hd__or4_4
XANTENNA__14476__B1 _14384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24773__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24965_ _24967_/CLK _24965_/D HRESETn VGND VGND VPWR VPWR _13898_/B sky130_fd_sc_hd__dfrtp_4
X_20088_ _20088_/A VGND VGND VPWR VPWR _20088_/X sky130_fd_sc_hd__buf_2
XFILLER_134_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24702__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25138__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11930_ _17443_/A VGND VGND VPWR VPWR _11948_/B sky130_fd_sc_hd__inv_2
X_23916_ _23916_/CLK _18928_/X VGND VGND VPWR VPWR _18927_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24896_ _24678_/CLK _24896_/D HRESETn VGND VGND VPWR VPWR _24896_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14228__B1 _13521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19926__A1_N _19924_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11861_ _11860_/Y _11864_/B VGND VGND VPWR VPWR _11861_/Y sky130_fd_sc_hd__nor2_4
X_23847_ _23846_/CLK _19129_/X VGND VGND VPWR VPWR _19128_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_249_0_HCLK clkbuf_7_124_0_HCLK/X VGND VGND VPWR VPWR _24146_/CLK sky130_fd_sc_hd__clkbuf_1
X_13600_ _13600_/A VGND VGND VPWR VPWR _19116_/B sky130_fd_sc_hd__buf_2
XPHY_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14561_/B _14575_/X _14578_/X _14579_/X _25093_/Q VGND VGND VPWR VPWR _25093_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _13797_/A VGND VGND VPWR VPWR _13459_/A sky130_fd_sc_hd__buf_2
X_23778_ _23774_/CLK _23778_/D VGND VGND VPWR VPWR _23778_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13451__B2 _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18914__B1 _17415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13531_ _25266_/Q VGND VGND VPWR VPWR _13531_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22729_ _24595_/Q _22729_/B VGND VGND VPWR VPWR _22733_/B sky130_fd_sc_hd__or2_4
X_25517_ _25499_/CLK _11870_/X HRESETn VGND VGND VPWR VPWR _11796_/B sky130_fd_sc_hd__dfrtp_4
XPHY_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18390__A1 _24109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16250_ _16249_/Y _16245_/X _16055_/X _16245_/X VGND VGND VPWR VPWR _16250_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13462_ _12058_/C _12057_/X _13462_/C _13456_/X VGND VGND VPWR VPWR _13462_/X sky130_fd_sc_hd__or4_4
X_25448_ _25453_/CLK _12444_/X HRESETn VGND VGND VPWR VPWR _12236_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23266__A2 _23257_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15201_ _14982_/A _15201_/B _15200_/X VGND VGND VPWR VPWR _15201_/X sky130_fd_sc_hd__or3_4
XFILLER_139_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12413_ _12413_/A _12413_/B _12412_/X VGND VGND VPWR VPWR _25456_/D sky130_fd_sc_hd__and3_4
X_16181_ _16181_/A _16180_/X VGND VGND VPWR VPWR _16182_/A sky130_fd_sc_hd__or2_4
XANTENNA__15469__A _14392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13393_ _13393_/A _13393_/B _13392_/X VGND VGND VPWR VPWR _13394_/C sky130_fd_sc_hd__and3_4
X_25379_ _25373_/CLK _25379_/D HRESETn VGND VGND VPWR VPWR _12934_/A sky130_fd_sc_hd__dfrtp_4
X_15132_ _15132_/A VGND VGND VPWR VPWR _15361_/A sky130_fd_sc_hd__inv_2
X_12344_ _12344_/A VGND VGND VPWR VPWR _13046_/A sky130_fd_sc_hd__inv_2
XFILLER_154_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16153__B1 _16062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23018__A2 _21303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15063_ _15063_/A _14942_/Y _15063_/C _15062_/X VGND VGND VPWR VPWR _15063_/X sky130_fd_sc_hd__or4_4
X_19940_ _19939_/X VGND VGND VPWR VPWR _19946_/A sky130_fd_sc_hd__inv_2
X_12275_ _12275_/A _12275_/B _12275_/C _12274_/X VGND VGND VPWR VPWR _12275_/X sky130_fd_sc_hd__or4_4
XFILLER_126_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15900__B1 _15472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14014_ _14001_/A _14011_/Y _14034_/C _14014_/D VGND VGND VPWR VPWR _14014_/X sky130_fd_sc_hd__or4_4
XFILLER_175_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19871_ _19871_/A VGND VGND VPWR VPWR _19871_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18822_ _18744_/A _18815_/X _18822_/C VGND VGND VPWR VPWR _24127_/D sky130_fd_sc_hd__and3_4
X_18753_ _18658_/Y _18748_/B _18735_/X _18749_/Y VGND VGND VPWR VPWR _18753_/X sky130_fd_sc_hd__a211o_4
X_15965_ _15965_/A VGND VGND VPWR VPWR _15965_/X sky130_fd_sc_hd__buf_2
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24443__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17704_ _11797_/Y _25515_/Q _17704_/C _11851_/X VGND VGND VPWR VPWR _17704_/X sky130_fd_sc_hd__or4_4
Xclkbuf_6_59_0_HCLK clkbuf_6_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14916_ _25015_/Q VGND VGND VPWR VPWR _15059_/A sky130_fd_sc_hd__inv_2
X_18684_ _18683_/Y _18819_/A _18815_/A VGND VGND VPWR VPWR _18786_/A sky130_fd_sc_hd__or3_4
XFILLER_64_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14219__B1 _13829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15896_ _15889_/A VGND VGND VPWR VPWR _15896_/X sky130_fd_sc_hd__buf_2
XFILLER_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17635_ _17543_/Y _17629_/X _17604_/X _17631_/Y VGND VGND VPWR VPWR _17636_/A sky130_fd_sc_hd__a211o_4
X_14847_ _14810_/A _14810_/B _14810_/A _14810_/B VGND VGND VPWR VPWR _14848_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15967__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17566_ _24307_/Q VGND VGND VPWR VPWR _17648_/A sky130_fd_sc_hd__inv_2
XFILLER_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14778_ _14771_/X VGND VGND VPWR VPWR _14778_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12559__A2_N _24868_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18905__B1 _24113_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19305_ _18032_/B VGND VGND VPWR VPWR _19305_/Y sky130_fd_sc_hd__inv_2
X_16517_ _16517_/A VGND VGND VPWR VPWR _16517_/Y sky130_fd_sc_hd__inv_2
X_13729_ _14761_/B VGND VGND VPWR VPWR _13729_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17497_ _17490_/X _17497_/B _17497_/C _17497_/D VGND VGND VPWR VPWR _17497_/X sky130_fd_sc_hd__or4_4
XFILLER_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19236_ _22222_/B _19233_/X _16864_/X _19233_/X VGND VGND VPWR VPWR _19236_/X sky130_fd_sc_hd__a2bb2o_4
X_16448_ _16721_/A _16721_/B _22629_/A _21327_/B VGND VGND VPWR VPWR _16448_/X sky130_fd_sc_hd__and4_4
XANTENNA__16392__B1 _16391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19167_ _23833_/Q VGND VGND VPWR VPWR _19167_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16379_ _15085_/Y _16376_/X _16004_/X _16376_/X VGND VGND VPWR VPWR _24607_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11700__A _11700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19330__B1 _19194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18118_ _18118_/A _18118_/B VGND VGND VPWR VPWR _18118_/X sky130_fd_sc_hd__or2_4
X_19098_ _23857_/Q VGND VGND VPWR VPWR _19098_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22931__C _22930_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18049_ _18193_/A _18983_/A VGND VGND VPWR VPWR _18050_/C sky130_fd_sc_hd__or2_4
XFILLER_160_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21060_ _22807_/A VGND VGND VPWR VPWR _21098_/A sky130_fd_sc_hd__buf_2
XANTENNA__22005__A _22004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21547__C _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20011_ _19455_/A _18288_/X _18285_/A _19960_/X VGND VGND VPWR VPWR _20012_/A sky130_fd_sc_hd__or4_4
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16340__A1_N _16339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14458__B1 _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16003__A _24743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24184__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19397__B1 _19395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17729__A1_N _17725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24750_ _24753_/CLK _24750_/D HRESETn VGND VGND VPWR VPWR _21534_/A sky130_fd_sc_hd__dfrtp_4
X_21962_ _21962_/A _21962_/B VGND VGND VPWR VPWR _21962_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24113__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15407__C1 _15334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23701_ _24208_/CLK _19541_/X VGND VGND VPWR VPWR _19538_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_215_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20913_ _16670_/Y _20846_/A _20855_/X _20912_/Y VGND VGND VPWR VPWR _20914_/A sky130_fd_sc_hd__o22a_4
XFILLER_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24681_ _24681_/CLK _16164_/X HRESETn VGND VGND VPWR VPWR _21064_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_55_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21893_ _21884_/A VGND VGND VPWR VPWR _22386_/A sky130_fd_sc_hd__buf_2
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23632_ _23458_/CLK _23632_/D VGND VGND VPWR VPWR _19745_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ _16706_/Y _20825_/X _20834_/X _20843_/Y VGND VGND VPWR VPWR _20844_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_2_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_16_0_HCLK clkbuf_7_8_0_HCLK/X VGND VGND VPWR VPWR _23437_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23563_ _23555_/CLK _23563_/D VGND VGND VPWR VPWR _19936_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20775_ _20774_/X VGND VGND VPWR VPWR _20775_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25319__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25302_ _23735_/CLK _25302_/D HRESETn VGND VGND VPWR VPWR _15908_/A sky130_fd_sc_hd__dfstp_4
Xclkbuf_8_79_0_HCLK clkbuf_8_79_0_HCLK/A VGND VGND VPWR VPWR _24696_/CLK sky130_fd_sc_hd__clkbuf_1
X_22514_ _22514_/A VGND VGND VPWR VPWR _22528_/B sky130_fd_sc_hd__inv_2
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23494_ _23494_/CLK _23494_/D VGND VGND VPWR VPWR _20125_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16383__B1 _16382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25233_ _23976_/CLK _25233_/D HRESETn VGND VGND VPWR VPWR _25233_/Q sky130_fd_sc_hd__dfrtp_4
X_22445_ _17849_/X _22437_/A _12755_/A _22444_/X VGND VGND VPWR VPWR _22445_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14933__B2 _14932_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25164_ _25164_/CLK _25164_/D HRESETn VGND VGND VPWR VPWR _14326_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22376_ _22383_/A _22376_/B _22376_/C VGND VGND VPWR VPWR _22376_/X sky130_fd_sc_hd__and3_4
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24115_ _24208_/CLK _24115_/D HRESETn VGND VGND VPWR VPWR _17443_/A sky130_fd_sc_hd__dfrtp_4
X_21327_ _21327_/A _21327_/B VGND VGND VPWR VPWR _21327_/X sky130_fd_sc_hd__or2_4
X_25095_ _24188_/CLK _25095_/D HRESETn VGND VGND VPWR VPWR _14547_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_191_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22759__A1 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12060_ _12060_/A VGND VGND VPWR VPWR _12060_/X sky130_fd_sc_hd__buf_2
X_24046_ _24427_/CLK _20879_/X HRESETn VGND VGND VPWR VPWR _24046_/Q sky130_fd_sc_hd__dfrtp_4
X_21258_ _22213_/A _21248_/X _21257_/X VGND VGND VPWR VPWR _21258_/X sky130_fd_sc_hd__or3_4
XFILLER_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20209_ _20208_/Y _20206_/X _19702_/X _20206_/X VGND VGND VPWR VPWR _23463_/D sky130_fd_sc_hd__a2bb2o_4
X_21189_ _21189_/A VGND VGND VPWR VPWR _21209_/A sky130_fd_sc_hd__buf_2
XANTENNA__14449__B1 _14407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15752__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12962_ _12775_/Y _12959_/B VGND VGND VPWR VPWR _12962_/Y sky130_fd_sc_hd__nand2_4
X_15750_ _15759_/A VGND VGND VPWR VPWR _15750_/X sky130_fd_sc_hd__buf_2
XFILLER_218_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24948_ _24947_/CLK _15488_/X HRESETn VGND VGND VPWR VPWR _14177_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_161_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11913_ _19977_/A VGND VGND VPWR VPWR _19613_/A sky130_fd_sc_hd__buf_2
X_14701_ _14701_/A VGND VGND VPWR VPWR _14701_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12893_ _12813_/Y _12892_/X VGND VGND VPWR VPWR _12896_/B sky130_fd_sc_hd__or2_4
X_15681_ _15681_/A VGND VGND VPWR VPWR _15681_/X sky130_fd_sc_hd__buf_2
X_24879_ _24874_/CLK _24879_/D HRESETn VGND VGND VPWR VPWR _24879_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17420_ _24331_/Q VGND VGND VPWR VPWR _17420_/Y sky130_fd_sc_hd__inv_2
X_11844_ _11844_/A VGND VGND VPWR VPWR _11844_/Y sky130_fd_sc_hd__inv_2
X_14632_ _14630_/C VGND VGND VPWR VPWR _14632_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14563_/A _14563_/B _14563_/C _25097_/Q VGND VGND VPWR VPWR _14563_/X sky130_fd_sc_hd__and4_4
X_17351_ _17351_/A _17351_/B _17350_/X VGND VGND VPWR VPWR _24352_/D sky130_fd_sc_hd__and3_4
XPHY_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _14380_/A VGND VGND VPWR VPWR _11775_/X sky130_fd_sc_hd__buf_2
XFILLER_198_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16300_/Y _16298_/X _16301_/X _16298_/X VGND VGND VPWR VPWR _24635_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _25308_/Q _13512_/Y _13513_/X _13509_/X VGND VGND VPWR VPWR _13514_/X sky130_fd_sc_hd__a211o_4
X_14494_ _14490_/C VGND VGND VPWR VPWR _14494_/X sky130_fd_sc_hd__buf_2
X_17282_ _17175_/Y _17280_/A VGND VGND VPWR VPWR _17282_/X sky130_fd_sc_hd__or2_4
XFILLER_41_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16374__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19021_ _19020_/Y _19018_/X _18951_/X _19018_/X VGND VGND VPWR VPWR _23884_/D sky130_fd_sc_hd__a2bb2o_4
X_13445_ _13445_/A _19758_/A VGND VGND VPWR VPWR _13447_/B sky130_fd_sc_hd__or2_4
X_16233_ _16233_/A VGND VGND VPWR VPWR _16233_/X sky130_fd_sc_hd__buf_2
XANTENNA__15199__A _15165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22447__B1 _25441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12616__A _12680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22998__A1 _16566_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13376_ _13268_/X _13376_/B _13375_/X VGND VGND VPWR VPWR _13376_/X sky130_fd_sc_hd__and3_4
X_16164_ _16163_/Y _16086_/A _15475_/X _16086_/A VGND VGND VPWR VPWR _16164_/X sky130_fd_sc_hd__a2bb2o_4
X_12327_ _12317_/X _12327_/B _12327_/C _12327_/D VGND VGND VPWR VPWR _12328_/D sky130_fd_sc_hd__or4_4
X_15115_ _15105_/X _15108_/X _15111_/X _15115_/D VGND VGND VPWR VPWR _15115_/X sky130_fd_sc_hd__or4_4
X_16095_ _16094_/Y _16092_/X _16001_/X _16092_/X VGND VGND VPWR VPWR _24709_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24695__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15046_ _15046_/A VGND VGND VPWR VPWR _15046_/Y sky130_fd_sc_hd__inv_2
X_19923_ _19922_/Y _19920_/X _19603_/X _19920_/X VGND VGND VPWR VPWR _19923_/X sky130_fd_sc_hd__a2bb2o_4
X_12258_ _12257_/Y _22276_/A _12252_/X _24751_/Q VGND VGND VPWR VPWR _12259_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24624__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19854_ _19854_/A VGND VGND VPWR VPWR _22339_/B sky130_fd_sc_hd__inv_2
X_12189_ _12187_/A _22857_/A _12187_/Y _12188_/Y VGND VGND VPWR VPWR _12189_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18805_ _18788_/B _18812_/B VGND VGND VPWR VPWR _18809_/B sky130_fd_sc_hd__or2_4
XANTENNA__21664__A _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19785_ _19782_/Y _19784_/X _18250_/X _19784_/X VGND VGND VPWR VPWR _23618_/D sky130_fd_sc_hd__a2bb2o_4
X_16997_ _16014_/Y _17024_/A _16014_/Y _17024_/A VGND VGND VPWR VPWR _17000_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15662__A _15662_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18736_ _18730_/A _18730_/B _18735_/X _18732_/B VGND VGND VPWR VPWR _18736_/X sky130_fd_sc_hd__a211o_4
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15948_ HWDATA[19] VGND VGND VPWR VPWR _15948_/X sky130_fd_sc_hd__buf_2
XFILLER_209_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18667_ _16605_/Y _24132_/Q _16613_/Y _18683_/A VGND VGND VPWR VPWR _18668_/D sky130_fd_sc_hd__a2bb2o_4
X_15879_ _15700_/X VGND VGND VPWR VPWR _15879_/X sky130_fd_sc_hd__buf_2
XANTENNA__13182__A _11950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17618_ _17564_/Y _17616_/X _17617_/Y VGND VGND VPWR VPWR _17618_/X sky130_fd_sc_hd__o21a_4
X_18598_ _18598_/A VGND VGND VPWR VPWR _24158_/D sky130_fd_sc_hd__inv_2
XANTENNA__25483__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14612__B1 _14611_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_232_0_HCLK clkbuf_7_116_0_HCLK/X VGND VGND VPWR VPWR _25230_/CLK sky130_fd_sc_hd__clkbuf_1
X_17549_ _17549_/A VGND VGND VPWR VPWR _17587_/A sky130_fd_sc_hd__inv_2
XFILLER_211_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20560_ _14430_/Y _20543_/X _20557_/X _20559_/X VGND VGND VPWR VPWR _20560_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16722__A2_N _16721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19219_ _19218_/Y _19216_/X _19194_/X _19216_/X VGND VGND VPWR VPWR _19219_/X sky130_fd_sc_hd__a2bb2o_4
X_20491_ _23966_/Q _20479_/B _20477_/C VGND VGND VPWR VPWR _20491_/X sky130_fd_sc_hd__and3_4
XFILLER_164_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22230_ _19528_/A _22001_/Y _22051_/X _22229_/X VGND VGND VPWR VPWR _22231_/A sky130_fd_sc_hd__a211o_4
XFILLER_164_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16117__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22453__A3 _16724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22161_ _14885_/A _22807_/A _23001_/A _22160_/X VGND VGND VPWR VPWR _22161_/X sky130_fd_sc_hd__a211o_4
XFILLER_161_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21112_ _15985_/B VGND VGND VPWR VPWR _22429_/A sky130_fd_sc_hd__buf_2
X_22092_ _11704_/A VGND VGND VPWR VPWR _22417_/B sky130_fd_sc_hd__buf_2
XANTENNA__24365__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17617__B1 _17593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21043_ _24819_/Q _21089_/B VGND VGND VPWR VPWR _21043_/X sky130_fd_sc_hd__and2_4
XFILLER_114_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24802_ _24804_/CLK _15878_/X HRESETn VGND VGND VPWR VPWR _24802_/Q sky130_fd_sc_hd__dfrtp_4
X_22994_ _23062_/A _22993_/X VGND VGND VPWR VPWR _22994_/Y sky130_fd_sc_hd__nor2_4
XFILLER_86_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_42_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_85_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21945_ _21462_/A _21945_/B _21944_/X VGND VGND VPWR VPWR _21945_/X sky130_fd_sc_hd__and3_4
X_24733_ _24737_/CLK _16030_/X HRESETn VGND VGND VPWR VPWR _24733_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19790__B1 _19746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24664_ _24667_/CLK _24664_/D HRESETn VGND VGND VPWR VPWR _22814_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_231_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _24752_/Q _22136_/B _22816_/A _24824_/Q _23138_/A VGND VGND VPWR VPWR _21876_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_215_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23615_ _23627_/CLK _23615_/D VGND VGND VPWR VPWR _19791_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _20827_/A VGND VGND VPWR VPWR _20919_/A sky130_fd_sc_hd__buf_2
XFILLER_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24595_ _24594_/CLK _24595_/D HRESETn VGND VGND VPWR VPWR _24595_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23546_ _23415_/CLK _19992_/X VGND VGND VPWR VPWR _19988_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20758_ _20753_/X _20756_/Y _24908_/Q _20757_/X VGND VGND VPWR VPWR _24018_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16356__B1 _15976_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23013__B _22817_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23477_ _25510_/CLK _23477_/D VGND VGND VPWR VPWR _23477_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20689_ _20716_/A VGND VGND VPWR VPWR _20780_/A sky130_fd_sc_hd__buf_2
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13345_/A _13224_/X _13230_/C VGND VGND VPWR VPWR _13230_/X sky130_fd_sc_hd__or3_4
X_25216_ _25224_/CLK _25216_/D HRESETn VGND VGND VPWR VPWR _14103_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__12917__B1 _12862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22428_ _21099_/X VGND VGND VPWR VPWR _22781_/A sky130_fd_sc_hd__buf_2
XANTENNA__13185__A3 _13184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13161_ _13187_/A VGND VGND VPWR VPWR _13394_/A sky130_fd_sc_hd__buf_2
X_25147_ _25146_/CLK _25147_/D HRESETn VGND VGND VPWR VPWR _14388_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_170_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22359_ _21936_/A _22359_/B VGND VGND VPWR VPWR _22359_/X sky130_fd_sc_hd__or2_4
XFILLER_124_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12112_ _12111_/Y _12107_/X _11793_/X _12107_/X VGND VGND VPWR VPWR _25469_/D sky130_fd_sc_hd__a2bb2o_4
X_13092_ _13069_/A _13069_/B _13090_/B _13019_/X VGND VGND VPWR VPWR _13092_/X sky130_fd_sc_hd__a211o_4
X_25078_ _23889_/CLK _25078_/D HRESETn VGND VGND VPWR VPWR _25078_/Q sky130_fd_sc_hd__dfrtp_4
X_12043_ _12043_/A VGND VGND VPWR VPWR _12043_/Y sky130_fd_sc_hd__inv_2
X_16920_ _16892_/X _16920_/B _16910_/X _16920_/D VGND VGND VPWR VPWR _16950_/A sky130_fd_sc_hd__or4_4
X_24029_ _24060_/CLK _20804_/X HRESETn VGND VGND VPWR VPWR _13106_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_49_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24035__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_124_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_124_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16851_ _14939_/Y _16793_/X _16787_/X _16793_/X VGND VGND VPWR VPWR _24415_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15802_ _12356_/Y _15796_/X _11695_/X _15796_/X VGND VGND VPWR VPWR _24842_/D sky130_fd_sc_hd__a2bb2o_4
X_19570_ _19570_/A _21159_/A VGND VGND VPWR VPWR _19570_/X sky130_fd_sc_hd__or2_4
XFILLER_19_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16782_ HWDATA[3] VGND VGND VPWR VPWR _18965_/A sky130_fd_sc_hd__buf_2
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13994_ _13994_/A VGND VGND VPWR VPWR _13995_/D sky130_fd_sc_hd__inv_2
XFILLER_218_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18521_ _18823_/B _18521_/B _18520_/X VGND VGND VPWR VPWR _18522_/A sky130_fd_sc_hd__or3_4
X_15733_ _12543_/Y _15731_/X _11718_/X _15731_/X VGND VGND VPWR VPWR _15733_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_246_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12945_ _12756_/X _12931_/X _12872_/A _12941_/Y VGND VGND VPWR VPWR _12945_/X sky130_fd_sc_hd__a211o_4
XFILLER_234_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18452_ _18452_/A _18438_/X _18446_/X _18452_/D VGND VGND VPWR VPWR _18453_/B sky130_fd_sc_hd__or4_4
X_15664_ _15663_/X VGND VGND VPWR VPWR _21587_/A sky130_fd_sc_hd__buf_2
XFILLER_234_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16595__B1 _16420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ _12759_/Y _12885_/B VGND VGND VPWR VPWR _12879_/B sky130_fd_sc_hd__or2_4
XPHY_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15937__A3 _15719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17384_/X _17398_/X _21002_/B _24339_/Q _17401_/X VGND VGND VPWR VPWR _17403_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _14615_/A VGND VGND VPWR VPWR _21968_/A sky130_fd_sc_hd__inv_2
X_11827_ _24236_/Q VGND VGND VPWR VPWR _22541_/A sky130_fd_sc_hd__inv_2
X_18383_ _24194_/Q VGND VGND VPWR VPWR _18383_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22668__B1 _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _24908_/Q VGND VGND VPWR VPWR _15595_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11959__A1 _18900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11959__B2 _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17246_/Y _17333_/X VGND VGND VPWR VPWR _17335_/A sky130_fd_sc_hd__or2_4
XFILLER_81_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11755_/Y _11756_/X _11757_/X _11756_/X VGND VGND VPWR VPWR _25528_/D sky130_fd_sc_hd__a2bb2o_4
X_14546_ _14566_/D VGND VGND VPWR VPWR _14546_/X sky130_fd_sc_hd__buf_2
XFILLER_60_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16347__B1 _16062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21340__B1 _21339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_62_0_HCLK clkbuf_8_63_0_HCLK/A VGND VGND VPWR VPWR _25089_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17265_ _17265_/A _17264_/X VGND VGND VPWR VPWR _17265_/X sky130_fd_sc_hd__or2_4
X_11689_ _11687_/Y _11684_/X _11688_/X _11684_/X VGND VGND VPWR VPWR _25544_/D sky130_fd_sc_hd__a2bb2o_4
X_14477_ _14477_/A VGND VGND VPWR VPWR _14477_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19004_ _19011_/A VGND VGND VPWR VPWR _19004_/X sky130_fd_sc_hd__buf_2
XANTENNA__24876__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16216_ _16214_/Y _16210_/X _15948_/X _16215_/X VGND VGND VPWR VPWR _16216_/X sky130_fd_sc_hd__a2bb2o_4
X_13428_ _13396_/A _18953_/A VGND VGND VPWR VPWR _13429_/C sky130_fd_sc_hd__or2_4
XFILLER_162_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23093__B1 _12309_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17196_ _24343_/Q VGND VGND VPWR VPWR _17242_/B sky130_fd_sc_hd__inv_2
XANTENNA__24805__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21729__A2_N _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13359_ _13391_/A _23813_/Q VGND VGND VPWR VPWR _13361_/B sky130_fd_sc_hd__or2_4
X_16147_ _22405_/A VGND VGND VPWR VPWR _16147_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16078_ _11699_/X _15651_/A _15920_/X _24714_/Q _16077_/X VGND VGND VPWR VPWR _24714_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__13177__A _13157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15029_ _15065_/A _24469_/Q _15065_/A _24469_/Q VGND VGND VPWR VPWR _15029_/X sky130_fd_sc_hd__a2bb2o_4
X_19906_ _22084_/B _19900_/X _19813_/X _19905_/X VGND VGND VPWR VPWR _19906_/X sky130_fd_sc_hd__a2bb2o_4
X_19837_ _19837_/A VGND VGND VPWR VPWR _22209_/B sky130_fd_sc_hd__inv_2
XFILLER_229_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19768_ _19768_/A VGND VGND VPWR VPWR _19768_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18719_ _18774_/A _18697_/X VGND VGND VPWR VPWR _18719_/X sky130_fd_sc_hd__or2_4
Xclkbuf_5_29_0_HCLK clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19699_ _19694_/A VGND VGND VPWR VPWR _19699_/X sky130_fd_sc_hd__buf_2
XFILLER_232_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21730_ _21730_/A _21730_/B VGND VGND VPWR VPWR _21730_/X sky130_fd_sc_hd__and2_4
XFILLER_213_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16586__B1 _16229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21661_ _21661_/A _20340_/Y VGND VGND VPWR VPWR _21663_/B sky130_fd_sc_hd__or2_4
XANTENNA__22659__B1 _24868_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23400_ _25272_/CLK _20373_/X VGND VGND VPWR VPWR _23400_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_212_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20612_ _15451_/X VGND VGND VPWR VPWR _20613_/B sky130_fd_sc_hd__buf_2
X_24380_ _24725_/CLK _24380_/D HRESETn VGND VGND VPWR VPWR _24380_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16338__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21592_ _21592_/A VGND VGND VPWR VPWR _22290_/A sky130_fd_sc_hd__buf_2
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20134__B2 _20116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22953__A _24600_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23331_ _24546_/Q _23171_/X _22839_/X _23330_/X VGND VGND VPWR VPWR _23331_/X sky130_fd_sc_hd__a211o_4
XFILLER_177_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20543_ _20543_/A VGND VGND VPWR VPWR _20543_/X sky130_fd_sc_hd__buf_2
XFILLER_124_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23262_ _15104_/A _23088_/B VGND VGND VPWR VPWR _23265_/B sky130_fd_sc_hd__or2_4
XFILLER_193_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20474_ _23966_/Q VGND VGND VPWR VPWR _20502_/B sky130_fd_sc_hd__inv_2
X_25001_ _24953_/CLK _15336_/X HRESETn VGND VGND VPWR VPWR _15075_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24546__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22213_ _22213_/A _22213_/B _22213_/C VGND VGND VPWR VPWR _22213_/X sky130_fd_sc_hd__and3_4
XANTENNA__15567__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23193_ _23193_/A _23156_/X VGND VGND VPWR VPWR _23193_/X sky130_fd_sc_hd__or2_4
XFILLER_118_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22144_ _21533_/A VGND VGND VPWR VPWR _22145_/B sky130_fd_sc_hd__buf_2
X_22075_ _22367_/A _22075_/B VGND VGND VPWR VPWR _22075_/X sky130_fd_sc_hd__or2_4
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21026_ _22466_/A VGND VGND VPWR VPWR _22423_/A sky130_fd_sc_hd__buf_2
XFILLER_102_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14824__B1 _14215_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22977_ _24633_/Q _22904_/X VGND VGND VPWR VPWR _22977_/X sky130_fd_sc_hd__or2_4
XANTENNA__25334__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12730_ _12934_/A VGND VGND VPWR VPWR _12830_/A sky130_fd_sc_hd__inv_2
X_24716_ _24639_/CLK _16074_/X HRESETn VGND VGND VPWR VPWR _24716_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_216_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19502__A _19501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21928_ _21922_/X _21927_/X _17725_/A VGND VGND VPWR VPWR _21928_/X sky130_fd_sc_hd__o21a_4
XFILLER_43_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16577__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12661_ _12661_/A VGND VGND VPWR VPWR _25421_/D sky130_fd_sc_hd__inv_2
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21859_ _21859_/A _21859_/B _21859_/C VGND VGND VPWR VPWR _21859_/X sky130_fd_sc_hd__and3_4
X_24647_ _24592_/CLK _16266_/X HRESETn VGND VGND VPWR VPWR _16265_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_188_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22114__A2 _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _14400_/A VGND VGND VPWR VPWR _14400_/X sky130_fd_sc_hd__buf_2
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23311__B2 _21871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12063__B1 _11765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12592_/A VGND VGND VPWR VPWR _12592_/Y sky130_fd_sc_hd__inv_2
X_15380_ _15123_/Y _15375_/B _15376_/Y _15334_/X VGND VGND VPWR VPWR _15380_/X sky130_fd_sc_hd__a211o_4
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24578_ _24080_/CLK _16455_/X HRESETn VGND VGND VPWR VPWR _24578_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ _25165_/Q _14330_/Y _14339_/A VGND VGND VPWR VPWR _25165_/D sky130_fd_sc_hd__o21a_4
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_49_0_HCLK clkbuf_6_24_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_98_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23529_ _24199_/CLK _23529_/D VGND VGND VPWR VPWR _23529_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25404__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _14262_/A VGND VGND VPWR VPWR _14262_/X sky130_fd_sc_hd__buf_2
X_17050_ _17050_/A _17050_/B VGND VGND VPWR VPWR _17051_/C sky130_fd_sc_hd__nand2_4
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24287__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13213_ _13199_/A VGND VGND VPWR VPWR _13260_/A sky130_fd_sc_hd__buf_2
X_16001_ HWDATA[28] VGND VGND VPWR VPWR _16001_/X sky130_fd_sc_hd__buf_2
X_14193_ _20510_/A _14188_/X _13826_/X _14190_/X VGND VGND VPWR VPWR _14193_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24216__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13144_ _13288_/A VGND VGND VPWR VPWR _13397_/A sky130_fd_sc_hd__buf_2
XFILLER_152_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13075_ _12981_/D _13074_/X VGND VGND VPWR VPWR _13079_/B sky130_fd_sc_hd__or2_4
X_17952_ _17949_/A _17952_/B VGND VGND VPWR VPWR _17952_/X sky130_fd_sc_hd__or2_4
X_12026_ _25490_/Q VGND VGND VPWR VPWR _12026_/Y sky130_fd_sc_hd__inv_2
X_16903_ _22870_/A _24276_/Q _16118_/Y _17761_/A VGND VGND VPWR VPWR _16910_/A sky130_fd_sc_hd__o22a_4
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18254__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17883_ _17752_/A _17885_/B _17882_/Y VGND VGND VPWR VPWR _24261_/D sky130_fd_sc_hd__o21a_4
XANTENNA__15924__B _15855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19622_ _19622_/A VGND VGND VPWR VPWR _21193_/B sky130_fd_sc_hd__inv_2
XFILLER_238_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16834_ _16841_/A VGND VGND VPWR VPWR _16834_/X sky130_fd_sc_hd__buf_2
XFILLER_76_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13827__A1_N _13538_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19553_ _22238_/B _19550_/X _11906_/X _19550_/X VGND VGND VPWR VPWR _19553_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21942__A _17709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16765_ _16765_/A VGND VGND VPWR VPWR _16765_/Y sky130_fd_sc_hd__inv_2
X_13977_ _13992_/A VGND VGND VPWR VPWR _14012_/A sky130_fd_sc_hd__buf_2
XANTENNA__25075__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18504_ _24185_/Q _18504_/B VGND VGND VPWR VPWR _18506_/B sky130_fd_sc_hd__or2_4
X_15716_ _12570_/Y _15714_/X _15560_/X _15714_/X VGND VGND VPWR VPWR _15716_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12928_ _12749_/Y _12588_/X VGND VGND VPWR VPWR _12958_/B sky130_fd_sc_hd__or2_4
X_19484_ _23721_/Q VGND VGND VPWR VPWR _22258_/B sky130_fd_sc_hd__inv_2
XFILLER_202_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16568__B1 _16483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25004__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16696_ _16696_/A VGND VGND VPWR VPWR _16696_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18435_ _16205_/Y _24181_/Q _16205_/Y _24181_/Q VGND VGND VPWR VPWR _18438_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_221_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15647_ _15639_/Y _15642_/X _15643_/X _21018_/B _15646_/X VGND VGND VPWR VPWR _24892_/D
+ sky130_fd_sc_hd__a32o_4
X_12859_ _25397_/Q _12859_/B VGND VGND VPWR VPWR _12861_/B sky130_fd_sc_hd__or2_4
XPHY_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23302__A1 _24476_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18366_ _18358_/X _18365_/Y _18350_/A _18357_/Y VGND VGND VPWR VPWR _24201_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22195__D _22194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15578_ _15578_/A VGND VGND VPWR VPWR _15578_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21313__B1 _24717_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17317_ _17314_/C _17305_/X VGND VGND VPWR VPWR _17318_/B sky130_fd_sc_hd__or2_4
X_14529_ scl_oen_o_S4 _14523_/X _14524_/Y _14528_/Y VGND VGND VPWR VPWR _14530_/B
+ sky130_fd_sc_hd__o22a_4
X_18297_ _18296_/X VGND VGND VPWR VPWR _18298_/B sky130_fd_sc_hd__inv_2
XFILLER_147_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12076__A _14262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17248_ _22709_/A VGND VGND VPWR VPWR _17248_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16740__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_6_0_HCLK clkbuf_6_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_17179_ _17179_/A VGND VGND VPWR VPWR _17179_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23100__C _23092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20190_ _20189_/Y _20185_/X _20102_/X _20185_/X VGND VGND VPWR VPWR _20190_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24921__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23939__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22592__A2 _21098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22900_ _22769_/A _22899_/X VGND VGND VPWR VPWR _22900_/X sky130_fd_sc_hd__and2_4
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23880_ _23844_/CLK _19034_/X VGND VGND VPWR VPWR _18046_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_229_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16011__A _24740_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22831_ _23075_/B VGND VGND VPWR VPWR _22831_/X sky130_fd_sc_hd__buf_2
XANTENNA__16271__A2 _15986_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22667__B _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22762_ _17757_/Y _21447_/X _12443_/A _21448_/X VGND VGND VPWR VPWR _22762_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21552__B1 _14158_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21713_ _21711_/X _21712_/X _21058_/X VGND VGND VPWR VPWR _21713_/X sky130_fd_sc_hd__or3_4
X_24501_ _24501_/CLK _24501_/D HRESETn VGND VGND VPWR VPWR _24501_/Q sky130_fd_sc_hd__dfrtp_4
X_25481_ _25479_/CLK _25481_/D HRESETn VGND VGND VPWR VPWR _25481_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22693_ _22469_/X _22689_/X _23062_/A _22692_/X VGND VGND VPWR VPWR _22694_/A sky130_fd_sc_hd__o22a_4
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24798__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21644_ _21215_/X VGND VGND VPWR VPWR _21960_/B sky130_fd_sc_hd__buf_2
X_24432_ _25028_/CLK _24432_/D HRESETn VGND VGND VPWR VPWR _14908_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_185_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24727__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24363_ _24629_/CLK _24363_/D HRESETn VGND VGND VPWR VPWR _23012_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_165_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13793__B1 _13791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ _21575_/A VGND VGND VPWR VPWR _21575_/X sky130_fd_sc_hd__buf_2
XFILLER_193_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23314_ _21520_/X _23313_/X _21522_/X _15980_/A _23152_/X VGND VGND VPWR VPWR _23315_/A
+ sky130_fd_sc_hd__a32o_4
X_20526_ _20526_/A VGND VGND VPWR VPWR _20526_/Y sky130_fd_sc_hd__inv_2
X_24294_ _24297_/CLK _24294_/D HRESETn VGND VGND VPWR VPWR _24294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16731__B1 _16459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15534__B2 _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24380__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23245_ _23213_/A _23245_/B _23245_/C VGND VGND VPWR VPWR _23246_/D sky130_fd_sc_hd__and3_4
XFILLER_153_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20457_ _20603_/A _20449_/X VGND VGND VPWR VPWR _20457_/X sky130_fd_sc_hd__and2_4
XFILLER_4_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23176_ _23176_/A VGND VGND VPWR VPWR _23213_/A sky130_fd_sc_hd__buf_2
X_20388_ _20387_/X VGND VGND VPWR VPWR _20389_/A sky130_fd_sc_hd__inv_2
XFILLER_137_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22127_ _13772_/C _22090_/X _22095_/X _22101_/X _22126_/X VGND VGND VPWR VPWR _22127_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_121_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22058_ _22386_/A _22058_/B VGND VGND VPWR VPWR _22058_/X sky130_fd_sc_hd__or2_4
XFILLER_88_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25515__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13900_ _13903_/A _13907_/B _13907_/A _13887_/Y VGND VGND VPWR VPWR _13900_/X sky130_fd_sc_hd__o22a_4
X_21009_ _23968_/Q _23969_/Q _21010_/B VGND VGND VPWR VPWR _21009_/X sky130_fd_sc_hd__o21a_4
XFILLER_248_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17017__A _17333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14880_ _25019_/Q VGND VGND VPWR VPWR _14880_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18251__A3 _18250_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22858__A _22146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21762__A _14678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13831_ _13536_/Y _13828_/X _13785_/X _13828_/X VGND VGND VPWR VPWR _25259_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18858__A1_N _24571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15470__B1 _15469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16856__A _14777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22335__A2 _22320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19736__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16550_ _16550_/A VGND VGND VPWR VPWR _16550_/Y sky130_fd_sc_hd__inv_2
X_13762_ _21283_/A VGND VGND VPWR VPWR _13807_/C sky130_fd_sc_hd__inv_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_12_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__21543__B1 _24718_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15501_ _24941_/Q VGND VGND VPWR VPWR _15501_/Y sky130_fd_sc_hd__inv_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12713_ _12692_/X _12713_/B _12722_/C VGND VGND VPWR VPWR _12713_/X sky130_fd_sc_hd__and3_4
XFILLER_189_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17211__B2 _17249_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16481_ _24568_/Q VGND VGND VPWR VPWR _16481_/Y sky130_fd_sc_hd__inv_2
X_13693_ _13686_/B _13667_/X _13692_/X _13690_/X _11806_/A VGND VGND VPWR VPWR _25293_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18220_ _18220_/A _18216_/X _18220_/C VGND VGND VPWR VPWR _18220_/X sky130_fd_sc_hd__or3_4
XANTENNA__13280__A _13150_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15432_ _15432_/A VGND VGND VPWR VPWR _15432_/X sky130_fd_sc_hd__buf_2
XANTENNA__22099__A1 _24552_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12644_ _12644_/A _12639_/X VGND VGND VPWR VPWR _12645_/C sky130_fd_sc_hd__nand2_4
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24468__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18151_ _18151_/A _23877_/Q VGND VGND VPWR VPWR _18151_/X sky130_fd_sc_hd__or2_4
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12575_ _12575_/A VGND VGND VPWR VPWR _12655_/A sky130_fd_sc_hd__inv_2
X_15363_ _15352_/A _15357_/X _15362_/Y VGND VGND VPWR VPWR _24994_/D sky130_fd_sc_hd__and3_4
XFILLER_200_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17102_ _17099_/C _17099_/D VGND VGND VPWR VPWR _17103_/B sky130_fd_sc_hd__or2_4
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ _12153_/Y VGND VGND VPWR VPWR _14314_/X sky130_fd_sc_hd__buf_2
X_18082_ _18082_/A VGND VGND VPWR VPWR _18132_/A sky130_fd_sc_hd__buf_2
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15294_ _15106_/Y _15294_/B _15294_/C _15294_/D VGND VGND VPWR VPWR _15294_/X sky130_fd_sc_hd__or4_4
XANTENNA__16722__B1 _16716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15525__B2 _15524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17033_ _24386_/Q VGND VGND VPWR VPWR _17120_/A sky130_fd_sc_hd__inv_2
XFILLER_156_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14245_ _14245_/A VGND VGND VPWR VPWR _14246_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_136_0_HCLK clkbuf_7_68_0_HCLK/X VGND VGND VPWR VPWR _23464_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_125_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24050__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15000__A _24475_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14176_ _12038_/B VGND VGND VPWR VPWR _14177_/B sky130_fd_sc_hd__inv_2
XANTENNA__22271__A1 _21284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_199_0_HCLK clkbuf_7_99_0_HCLK/X VGND VGND VPWR VPWR _24486_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13127_ _20685_/B VGND VGND VPWR VPWR _20688_/B sky130_fd_sc_hd__inv_2
XFILLER_124_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18984_ HWDATA[5] VGND VGND VPWR VPWR _18985_/A sky130_fd_sc_hd__buf_2
XFILLER_124_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18311__A _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13058_ _13087_/A VGND VGND VPWR VPWR _13085_/A sky130_fd_sc_hd__buf_2
X_17935_ _18016_/A VGND VGND VPWR VPWR _17940_/A sky130_fd_sc_hd__buf_2
XFILLER_39_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12009_ _12009_/A VGND VGND VPWR VPWR _12009_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13455__A _21568_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22574__A2 _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17866_ _17866_/A _17866_/B _17865_/X VGND VGND VPWR VPWR _17866_/X sky130_fd_sc_hd__and3_4
XANTENNA__20955__A1_N _20828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18242__A3 _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16693__A1_N _16691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16817_ _14922_/Y _16813_/X HWDATA[19] _16816_/X VGND VGND VPWR VPWR _16817_/X sky130_fd_sc_hd__a2bb2o_4
X_19605_ _19605_/A VGND VGND VPWR VPWR _19605_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17797_ _16906_/Y _17796_/X VGND VGND VPWR VPWR _17800_/B sky130_fd_sc_hd__or2_4
XANTENNA__15461__B1 _14403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19536_ _23702_/Q VGND VGND VPWR VPWR _19536_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15670__A _16368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19142__A _19141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16748_ _24465_/Q VGND VGND VPWR VPWR _16748_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19467_ _23726_/Q VGND VGND VPWR VPWR _21813_/B sky130_fd_sc_hd__inv_2
XFILLER_179_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16679_ _16679_/A VGND VGND VPWR VPWR _16679_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18981__A _18981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13190__A _13285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24891__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18418_ _24167_/Q VGND VGND VPWR VPWR _18567_/A sky130_fd_sc_hd__inv_2
X_19398_ _18073_/B VGND VGND VPWR VPWR _19398_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16961__B1 _16031_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24820__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21837__A1 _14220_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18349_ _13175_/A _18341_/Y _18346_/X VGND VGND VPWR VPWR _18349_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21837__B2 _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24138__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21360_ _13482_/B _21358_/X _12087_/B _21359_/X VGND VGND VPWR VPWR _21360_/X sky130_fd_sc_hd__o22a_4
XFILLER_238_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_32_0_HCLK clkbuf_7_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_32_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20311_ _20306_/X _19573_/X _11760_/X _22400_/A _20310_/X VGND VGND VPWR VPWR _20311_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_7_95_0_HCLK clkbuf_7_95_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_95_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21291_ _21592_/A VGND VGND VPWR VPWR _21598_/A sky130_fd_sc_hd__inv_2
X_23030_ _16108_/Y _22559_/X _22849_/X _11694_/Y _21051_/A VGND VGND VPWR VPWR _23030_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__17269__A1 _17232_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20242_ _20242_/A VGND VGND VPWR VPWR _20243_/A sky130_fd_sc_hd__inv_2
XFILLER_190_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15845__A _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12750__B2 _24785_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20173_ _20173_/A VGND VGND VPWR VPWR _21405_/B sky130_fd_sc_hd__inv_2
XFILLER_170_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_HCLK clkbuf_3_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_24981_ _24980_/CLK _24981_/D HRESETn VGND VGND VPWR VPWR _15405_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_229_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23932_ _23932_/CLK _23932_/D HRESETn VGND VGND VPWR VPWR _20990_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_97_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22678__A _16272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21582__A _21582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23863_ _23808_/CLK _19082_/X VGND VGND VPWR VPWR _23863_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24979__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22814_ _22814_/A _22729_/B VGND VGND VPWR VPWR _22819_/B sky130_fd_sc_hd__or2_4
XFILLER_199_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23794_ _23754_/CLK _19277_/X VGND VGND VPWR VPWR _23794_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20198__A _17952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24908__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25533_ _25533_/CLK _11740_/X HRESETn VGND VGND VPWR VPWR _11737_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20186__A2_N _20180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22745_ _24800_/Q _22630_/B VGND VGND VPWR VPWR _22745_/X sky130_fd_sc_hd__or2_4
XANTENNA__12709__A _12680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22676_ _22676_/A VGND VGND VPWR VPWR _22676_/Y sky130_fd_sc_hd__inv_2
X_25464_ _25382_/CLK _25464_/D HRESETn VGND VGND VPWR VPWR _12167_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_198_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24561__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21627_ _21627_/A VGND VGND VPWR VPWR _22380_/A sky130_fd_sc_hd__buf_2
X_24415_ _24477_/CLK _24415_/D HRESETn VGND VGND VPWR VPWR _24415_/Q sky130_fd_sc_hd__dfrtp_4
X_25395_ _25397_/CLK _12869_/X HRESETn VGND VGND VPWR VPWR _12735_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12360_ _25338_/Q VGND VGND VPWR VPWR _12360_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21558_ _21558_/A _21722_/B VGND VGND VPWR VPWR _21558_/Y sky130_fd_sc_hd__nor2_4
X_24346_ _24346_/CLK _17370_/X HRESETn VGND VGND VPWR VPWR _24346_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20509_ _24002_/Q _20448_/X _20469_/X VGND VGND VPWR VPWR _24002_/D sky130_fd_sc_hd__a21o_4
XFILLER_4_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12291_ _12291_/A VGND VGND VPWR VPWR _12291_/X sky130_fd_sc_hd__buf_2
X_24277_ _25450_/CLK _17823_/X HRESETn VGND VGND VPWR VPWR _24277_/Q sky130_fd_sc_hd__dfrtp_4
X_21489_ _22257_/A VGND VGND VPWR VPWR _21489_/X sky130_fd_sc_hd__buf_2
XFILLER_154_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14030_ _14029_/X VGND VGND VPWR VPWR _14030_/Y sky130_fd_sc_hd__inv_2
X_23228_ _22286_/X _23218_/X _23228_/C _23228_/D VGND VGND VPWR VPWR _23228_/X sky130_fd_sc_hd__or4_4
XFILLER_180_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14191__B1 _13824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_209_0_HCLK clkbuf_7_104_0_HCLK/X VGND VGND VPWR VPWR _24051_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_181_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23159_ _23108_/X _23154_/Y _23155_/X _23158_/X VGND VGND VPWR VPWR _23159_/X sky130_fd_sc_hd__a2bb2o_4
X_15981_ _15981_/A VGND VGND VPWR VPWR _21745_/B sky130_fd_sc_hd__buf_2
XFILLER_67_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17720_ _17720_/A VGND VGND VPWR VPWR _21473_/A sky130_fd_sc_hd__buf_2
XFILLER_48_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14932_ _14932_/A VGND VGND VPWR VPWR _14932_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18785__B _18745_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17651_ _24306_/Q _17651_/B VGND VGND VPWR VPWR _17652_/C sky130_fd_sc_hd__or2_4
X_14863_ _24953_/Q VGND VGND VPWR VPWR _14863_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19709__B1 _19708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16602_ _16600_/Y _16598_/X _16601_/X _16598_/X VGND VGND VPWR VPWR _16602_/X sky130_fd_sc_hd__a2bb2o_4
X_13814_ _13556_/Y _13810_/X _11739_/X _13813_/X VGND VGND VPWR VPWR _13814_/X sky130_fd_sc_hd__a2bb2o_4
X_17582_ _17660_/A _17582_/B _17581_/X VGND VGND VPWR VPWR _17628_/B sky130_fd_sc_hd__or3_4
XFILLER_90_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14794_ _14808_/C _14808_/B _14809_/A VGND VGND VPWR VPWR _14795_/B sky130_fd_sc_hd__or3_4
XFILLER_44_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19321_ _19321_/A VGND VGND VPWR VPWR _19327_/A sky130_fd_sc_hd__inv_2
XFILLER_90_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24649__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16533_ _16532_/Y _16528_/X _16435_/X _16528_/X VGND VGND VPWR VPWR _24549_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13745_ _13745_/A _13736_/Y VGND VGND VPWR VPWR _13745_/X sky130_fd_sc_hd__or2_4
XFILLER_232_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15640__D _14422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19252_ _13723_/A _13741_/D _13743_/X _14683_/X VGND VGND VPWR VPWR _19253_/A sky130_fd_sc_hd__or4_4
X_16464_ HWDATA[28] VGND VGND VPWR VPWR _16464_/X sky130_fd_sc_hd__buf_2
X_13676_ _13676_/A _13676_/B VGND VGND VPWR VPWR _13677_/B sky130_fd_sc_hd__or2_4
XFILLER_204_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16943__B1 _21435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18203_ _17987_/X _18203_/B VGND VGND VPWR VPWR _18203_/X sky130_fd_sc_hd__or2_4
X_15415_ _15410_/X _15415_/B _15402_/X VGND VGND VPWR VPWR _24978_/D sky130_fd_sc_hd__and3_4
X_12627_ _12650_/A VGND VGND VPWR VPWR _12627_/X sky130_fd_sc_hd__buf_2
X_19183_ _23826_/Q VGND VGND VPWR VPWR _19183_/Y sky130_fd_sc_hd__inv_2
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16395_ HWDATA[20] VGND VGND VPWR VPWR _16395_/X sky130_fd_sc_hd__buf_2
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24231__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18134_ _17966_/X _18133_/X _24245_/Q _18024_/X VGND VGND VPWR VPWR _18134_/X sky130_fd_sc_hd__o22a_4
X_15346_ _15331_/A _15331_/B VGND VGND VPWR VPWR _15347_/B sky130_fd_sc_hd__or2_4
XFILLER_129_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12558_ _12684_/A VGND VGND VPWR VPWR _12558_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_19_0_HCLK clkbuf_5_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_39_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18065_ _13597_/A VGND VGND VPWR VPWR _18103_/A sky130_fd_sc_hd__buf_2
XFILLER_8_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15277_ _15269_/A _15273_/X _15276_/Y VGND VGND VPWR VPWR _25010_/D sky130_fd_sc_hd__and3_4
X_12489_ _12252_/X _12491_/B _12488_/Y VGND VGND VPWR VPWR _12489_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15071__A2_N _16363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17016_ _17343_/B VGND VGND VPWR VPWR _17333_/A sky130_fd_sc_hd__buf_2
X_14228_ _14227_/Y _14225_/X _13521_/X _14225_/X VGND VGND VPWR VPWR _14228_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22795__A2 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15665__A _21587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14159_ _14154_/A VGND VGND VPWR VPWR _14159_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18967_ _18964_/Y _18960_/X _18965_/X _18966_/X VGND VGND VPWR VPWR _23902_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25090__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17880__A _17880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17918_ _13528_/X VGND VGND VPWR VPWR _17918_/Y sky130_fd_sc_hd__inv_2
X_18898_ _18896_/Y _18897_/Y _17440_/X _18897_/Y VGND VGND VPWR VPWR _18898_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17849_ _16904_/Y VGND VGND VPWR VPWR _17849_/X sky130_fd_sc_hd__buf_2
XFILLER_66_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20860_ _20859_/X VGND VGND VPWR VPWR _20860_/Y sky130_fd_sc_hd__inv_2
XFILLER_240_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19519_ _23707_/Q VGND VGND VPWR VPWR _21190_/B sky130_fd_sc_hd__inv_2
X_20791_ _15574_/Y _20708_/A _20716_/X _20790_/X VGND VGND VPWR VPWR _20791_/X sky130_fd_sc_hd__o22a_4
XFILLER_50_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24319__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22530_ _22530_/A VGND VGND VPWR VPWR _23301_/B sky130_fd_sc_hd__buf_2
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19600__A _19600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22461_ _11833_/Y _21955_/A _13562_/Y _22515_/A VGND VGND VPWR VPWR _22461_/X sky130_fd_sc_hd__o22a_4
XFILLER_210_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23122__A _16654_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14744__A _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21412_ _22202_/A _21412_/B VGND VGND VPWR VPWR _21412_/X sky130_fd_sc_hd__or2_4
X_24200_ _24257_/CLK _24200_/D HRESETn VGND VGND VPWR VPWR _21979_/A sky130_fd_sc_hd__dfrtp_4
X_25180_ _25479_/CLK _25180_/D HRESETn VGND VGND VPWR VPWR _14289_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22392_ _21515_/Y _22363_/X _13763_/X _22391_/X VGND VGND VPWR VPWR _22392_/Y sky130_fd_sc_hd__a22oi_4
X_24131_ _24139_/CLK _24131_/D HRESETn VGND VGND VPWR VPWR _24131_/Q sky130_fd_sc_hd__dfrtp_4
X_21343_ _21343_/A _21343_/B VGND VGND VPWR VPWR _21343_/X sky130_fd_sc_hd__or2_4
XFILLER_163_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23027__A3 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24062_ _24060_/CLK _20947_/Y HRESETn VGND VGND VPWR VPWR _13635_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23954__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21274_ _21177_/A VGND VGND VPWR VPWR _21274_/X sky130_fd_sc_hd__buf_2
XANTENNA__25178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23013_ _16303_/A _22817_/B _22817_/C VGND VGND VPWR VPWR _23013_/X sky130_fd_sc_hd__and3_4
X_20225_ _20224_/Y _20222_/X _19743_/X _20222_/X VGND VGND VPWR VPWR _23457_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25107__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_182_0_HCLK clkbuf_7_91_0_HCLK/X VGND VGND VPWR VPWR _23958_/CLK sky130_fd_sc_hd__clkbuf_1
X_20156_ _20156_/A VGND VGND VPWR VPWR _22387_/B sky130_fd_sc_hd__inv_2
Xclkbuf_8_39_0_HCLK clkbuf_8_39_0_HCLK/A VGND VGND VPWR VPWR _24257_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_104_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13807__B _13807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22538__A2 _21031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20087_ _20087_/A VGND VGND VPWR VPWR _20088_/A sky130_fd_sc_hd__buf_2
X_24964_ _24073_/CLK _15449_/X HRESETn VGND VGND VPWR VPWR _13892_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23915_ _23853_/CLK _18930_/X VGND VGND VPWR VPWR _23915_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_218_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24895_ _24037_/CLK _24895_/D HRESETn VGND VGND VPWR VPWR _24895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11860_ _11860_/A VGND VGND VPWR VPWR _11860_/Y sky130_fd_sc_hd__inv_2
X_23846_ _23846_/CLK _23846_/D VGND VGND VPWR VPWR _23846_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14779__A2 _14777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24742__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ HWDATA[0] VGND VGND VPWR VPWR _13797_/A sky130_fd_sc_hd__buf_2
XFILLER_198_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20989_ _20988_/X VGND VGND VPWR VPWR _23932_/D sky130_fd_sc_hd__inv_2
X_23777_ _24089_/CLK _19325_/X VGND VGND VPWR VPWR _23777_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _25260_/Q VGND VGND VPWR VPWR _13530_/Y sky130_fd_sc_hd__inv_2
X_25516_ _24679_/CLK _25516_/D HRESETn VGND VGND VPWR VPWR _11797_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22728_ _22800_/B VGND VGND VPWR VPWR _22729_/B sky130_fd_sc_hd__buf_2
XFILLER_40_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13461_ _25324_/Q VGND VGND VPWR VPWR _13461_/Y sky130_fd_sc_hd__inv_2
X_25447_ _25453_/CLK _25447_/D HRESETn VGND VGND VPWR VPWR _25447_/Q sky130_fd_sc_hd__dfrtp_4
X_22659_ _22129_/X _22658_/X _21541_/X _24868_/Q _21542_/X VGND VGND VPWR VPWR _22660_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_201_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15200_ _15064_/X _15167_/B _14995_/X VGND VGND VPWR VPWR _15200_/X sky130_fd_sc_hd__o21a_4
X_12412_ _25456_/Q _12412_/B VGND VGND VPWR VPWR _12412_/X sky130_fd_sc_hd__or2_4
X_16180_ _16180_/A VGND VGND VPWR VPWR _16180_/X sky130_fd_sc_hd__buf_2
XFILLER_139_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13392_ _13392_/A _13392_/B VGND VGND VPWR VPWR _13392_/X sky130_fd_sc_hd__or2_4
X_25378_ _25373_/CLK _12939_/Y HRESETn VGND VGND VPWR VPWR _25378_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15794__A1_N _12316_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15131_ _15130_/Y _24603_/Q _15130_/Y _24603_/Q VGND VGND VPWR VPWR _15136_/B sky130_fd_sc_hd__a2bb2o_4
X_12343_ _13017_/A _24843_/Q _13017_/A _24843_/Q VGND VGND VPWR VPWR _12343_/X sky130_fd_sc_hd__a2bb2o_4
X_24329_ _24326_/CLK _24329_/D HRESETn VGND VGND VPWR VPWR _17426_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22590__B _16368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12274_ _12187_/Y _12428_/B _12201_/Y _12176_/A VGND VGND VPWR VPWR _12274_/X sky130_fd_sc_hd__or4_4
X_15062_ _15062_/A _15214_/B _14921_/A _15062_/D VGND VGND VPWR VPWR _15062_/X sky130_fd_sc_hd__or4_4
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25530__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12714__A1 _12569_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20237__B1 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14013_ _14006_/A _13981_/X VGND VGND VPWR VPWR _14014_/D sky130_fd_sc_hd__or2_4
X_19870_ _19868_/Y _19869_/X _19617_/X _19869_/X VGND VGND VPWR VPWR _19870_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18821_ _18815_/A _18815_/B VGND VGND VPWR VPWR _18822_/C sky130_fd_sc_hd__nand2_4
XANTENNA__12805__A1_N _12804_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18752_ _18752_/A _18752_/B _18751_/X VGND VGND VPWR VPWR _24147_/D sky130_fd_sc_hd__and3_4
XFILLER_95_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15964_ _15930_/Y VGND VGND VPWR VPWR _15964_/X sky130_fd_sc_hd__buf_2
XFILLER_209_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17703_ _13807_/A _17703_/B _21177_/A _21176_/A VGND VGND VPWR VPWR _17703_/X sky130_fd_sc_hd__or4_4
X_14915_ _14913_/A _24438_/Q _15189_/A _14914_/Y VGND VGND VPWR VPWR _14915_/X sky130_fd_sc_hd__o22a_4
XFILLER_64_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18683_ _18683_/A VGND VGND VPWR VPWR _18683_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15895_ _12734_/Y _15892_/X _15619_/X _15892_/X VGND VGND VPWR VPWR _15895_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22111__A _22111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17634_ _17647_/A _17632_/X _17633_/X VGND VGND VPWR VPWR _24312_/D sky130_fd_sc_hd__and3_4
X_14846_ _14838_/X _14845_/Y _14796_/A _14838_/X VGND VGND VPWR VPWR _14846_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20960__A1 _20822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24483__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17565_ _17564_/Y _17511_/Y VGND VGND VPWR VPWR _17584_/C sky130_fd_sc_hd__or2_4
X_14777_ _14777_/A VGND VGND VPWR VPWR _14777_/X sky130_fd_sc_hd__buf_2
X_11989_ _25310_/Q _11977_/A _25310_/Q _11977_/A VGND VGND VPWR VPWR _11998_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19304_ _19303_/Y _19300_/X _19279_/X _19300_/X VGND VGND VPWR VPWR _23785_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24412__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16516_ _16515_/Y _16513_/X _16145_/X _16513_/X VGND VGND VPWR VPWR _16516_/X sky130_fd_sc_hd__a2bb2o_4
X_13728_ _13728_/A _13728_/B _24513_/Q VGND VGND VPWR VPWR _14761_/B sky130_fd_sc_hd__and3_4
X_17496_ _11650_/Y _17564_/A _11650_/Y _17564_/A VGND VGND VPWR VPWR _17497_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17859__B _17849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19235_ _19235_/A VGND VGND VPWR VPWR _22222_/B sky130_fd_sc_hd__inv_2
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16447_ _16446_/X VGND VGND VPWR VPWR _21327_/B sky130_fd_sc_hd__inv_2
XFILLER_149_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13659_ _25299_/Q _13657_/X _13658_/Y VGND VGND VPWR VPWR _25299_/D sky130_fd_sc_hd__o21a_4
XFILLER_220_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19166_ _19162_/Y _19165_/X _19144_/X _19165_/X VGND VGND VPWR VPWR _19166_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16378_ _15140_/Y _16376_/X _16001_/X _16376_/X VGND VGND VPWR VPWR _16378_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_185_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18117_ _17947_/A _18109_/X _18116_/X VGND VGND VPWR VPWR _18117_/X sky130_fd_sc_hd__and3_4
XFILLER_145_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15329_ _15282_/B _15324_/Y _15328_/X VGND VGND VPWR VPWR _15329_/X sky130_fd_sc_hd__or3_4
X_19097_ _19093_/Y _19096_/X _19006_/X _19096_/X VGND VGND VPWR VPWR _23858_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25144__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18048_ _18004_/X _18048_/B VGND VGND VPWR VPWR _18050_/B sky130_fd_sc_hd__or2_4
XFILLER_160_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21397__A _22202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20228__B1 _19746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20010_ _23538_/Q VGND VGND VPWR VPWR _22340_/B sky130_fd_sc_hd__inv_2
Xclkbuf_8_255_0_HCLK clkbuf_8_255_0_HCLK/A VGND VGND VPWR VPWR _24973_/CLK sky130_fd_sc_hd__clkbuf_1
X_19999_ _19998_/Y _19996_/X _19974_/X _19996_/X VGND VGND VPWR VPWR _23543_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21961_ _18263_/X _21959_/X _21960_/X _13774_/Y _21643_/X VGND VGND VPWR VPWR _21962_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_66_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23700_ _24208_/CLK _19544_/X VGND VGND VPWR VPWR _23700_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20912_ _13636_/D _20907_/X _20916_/B VGND VGND VPWR VPWR _20912_/Y sky130_fd_sc_hd__a21oi_4
X_21892_ _22083_/A _19261_/Y VGND VGND VPWR VPWR _21892_/X sky130_fd_sc_hd__or2_4
X_24680_ _23665_/CLK _16175_/X HRESETn VGND VGND VPWR VPWR _13725_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_199_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _24039_/Q _13642_/X _20842_/Y VGND VGND VPWR VPWR _20843_/Y sky130_fd_sc_hd__a21oi_4
X_23631_ _23464_/CLK _23631_/D VGND VGND VPWR VPWR _19749_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24153__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20774_ _22922_/A _20708_/A _20716_/X _20773_/Y VGND VGND VPWR VPWR _20774_/X sky130_fd_sc_hd__o22a_4
X_23562_ _23559_/CLK _19942_/X VGND VGND VPWR VPWR _23562_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21900__B1 _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25301_ _25308_/CLK _25301_/D HRESETn VGND VGND VPWR VPWR _13513_/B sky130_fd_sc_hd__dfstp_4
XFILLER_195_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22513_ _13800_/X _22511_/X _21596_/X _22512_/X VGND VGND VPWR VPWR _22514_/A sky130_fd_sc_hd__o22a_4
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23493_ _23476_/CLK _20129_/X VGND VGND VPWR VPWR _20127_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_149_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22444_ _21022_/A VGND VGND VPWR VPWR _22444_/X sky130_fd_sc_hd__buf_2
X_25232_ _23976_/CLK _14074_/X HRESETn VGND VGND VPWR VPWR _13991_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_183_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22691__A _22435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25359__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22375_ _22387_/A _22375_/B VGND VGND VPWR VPWR _22376_/C sky130_fd_sc_hd__or2_4
X_25163_ _25140_/CLK _25163_/D HRESETn VGND VGND VPWR VPWR _14338_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_191_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21326_ _15662_/A VGND VGND VPWR VPWR _23001_/A sky130_fd_sc_hd__buf_2
X_24114_ _24618_/CLK _18904_/X HRESETn VGND VGND VPWR VPWR _24114_/Q sky130_fd_sc_hd__dfrtp_4
X_25094_ _25098_/CLK _14577_/X HRESETn VGND VGND VPWR VPWR _25094_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15894__B1 _15616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21100__A _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21257_ _21251_/X _21256_/X _14672_/A VGND VGND VPWR VPWR _21257_/X sky130_fd_sc_hd__o21a_4
X_24045_ _24487_/CLK _20876_/X HRESETn VGND VGND VPWR VPWR _24045_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13818__A _15965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20208_ _18070_/B VGND VGND VPWR VPWR _20208_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18832__B1 _16536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21188_ _21205_/A _21188_/B VGND VGND VPWR VPWR _21188_/X sky130_fd_sc_hd__or2_4
XFILLER_77_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24994__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20139_ _20135_/Y _20138_/X _20089_/X _20138_/X VGND VGND VPWR VPWR _23490_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24923__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12961_ _12816_/Y _12963_/B _12960_/Y VGND VGND VPWR VPWR _12961_/X sky130_fd_sc_hd__o21a_4
X_24947_ _24947_/CLK _15490_/X HRESETn VGND VGND VPWR VPWR _12038_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12791__A1_N _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14700_ _14699_/X VGND VGND VPWR VPWR _14701_/A sky130_fd_sc_hd__buf_2
X_11912_ _11910_/Y _11907_/X _11911_/X _11907_/X VGND VGND VPWR VPWR _11912_/X sky130_fd_sc_hd__a2bb2o_4
X_15680_ _15680_/A VGND VGND VPWR VPWR _15681_/A sky130_fd_sc_hd__inv_2
XFILLER_205_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12892_ _12839_/D _12892_/B VGND VGND VPWR VPWR _12892_/X sky130_fd_sc_hd__or2_4
X_24878_ _24866_/CLK _15726_/X HRESETn VGND VGND VPWR VPWR _24878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_206_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14368__B _14425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14631_ _18062_/A _14630_/X _18062_/A _14630_/X VGND VGND VPWR VPWR _25078_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21770__A _22381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11843_ _11843_/A VGND VGND VPWR VPWR _13686_/A sky130_fd_sc_hd__inv_2
X_23829_ _23846_/CLK _23829_/D VGND VGND VPWR VPWR _23829_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _17237_/Y _17348_/A VGND VGND VPWR VPWR _17350_/X sky130_fd_sc_hd__or2_4
X_14562_ _14562_/A VGND VGND VPWR VPWR _14563_/B sky130_fd_sc_hd__inv_2
XPHY_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11774_/A VGND VGND VPWR VPWR _14380_/A sky130_fd_sc_hd__buf_2
XPHY_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ HWDATA[23] VGND VGND VPWR VPWR _16301_/X sky130_fd_sc_hd__buf_2
XFILLER_198_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13501_/Y _13513_/B VGND VGND VPWR VPWR _13513_/X sky130_fd_sc_hd__and2_4
XPHY_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281_ _24368_/Q _17280_/Y VGND VGND VPWR VPWR _17281_/X sky130_fd_sc_hd__or2_4
X_14493_ _25112_/Q _14492_/B _14491_/X _14492_/Y VGND VGND VPWR VPWR _14493_/X sky130_fd_sc_hd__a211o_4
X_19020_ _19020_/A VGND VGND VPWR VPWR _19020_/Y sky130_fd_sc_hd__inv_2
X_16232_ _24660_/Q VGND VGND VPWR VPWR _16232_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14385__B1 _14384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13444_ _13254_/A _13442_/X _13443_/X VGND VGND VPWR VPWR _13444_/X sky130_fd_sc_hd__and3_4
XFILLER_155_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16163_ _21064_/A VGND VGND VPWR VPWR _16163_/Y sky130_fd_sc_hd__inv_2
X_13375_ _13234_/X _13375_/B VGND VGND VPWR VPWR _13375_/X sky130_fd_sc_hd__or2_4
XFILLER_186_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25029__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15114_ _24994_/Q _24598_/Q _15292_/A _15113_/Y VGND VGND VPWR VPWR _15115_/D sky130_fd_sc_hd__o22a_4
XFILLER_170_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12326_ _12324_/A _24838_/Q _12324_/Y _12325_/Y VGND VGND VPWR VPWR _12327_/D sky130_fd_sc_hd__o22a_4
X_16094_ _23225_/A VGND VGND VPWR VPWR _16094_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15045_ _15066_/A _15046_/A _15207_/A _15047_/A VGND VGND VPWR VPWR _15045_/X sky130_fd_sc_hd__a2bb2o_4
X_19922_ _19922_/A VGND VGND VPWR VPWR _19922_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12257_ _25439_/Q VGND VGND VPWR VPWR _12257_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12188_ _22857_/A VGND VGND VPWR VPWR _12188_/Y sky130_fd_sc_hd__inv_2
X_19853_ _19851_/Y _19847_/X _19852_/X _19835_/A VGND VGND VPWR VPWR _19853_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18804_ _18804_/A _18810_/A VGND VGND VPWR VPWR _18812_/B sky130_fd_sc_hd__or2_4
Xclkbuf_8_22_0_HCLK clkbuf_8_22_0_HCLK/A VGND VGND VPWR VPWR _24317_/CLK sky130_fd_sc_hd__clkbuf_1
X_16996_ _16040_/Y _24386_/Q _16040_/Y _24386_/Q VGND VGND VPWR VPWR _17000_/A sky130_fd_sc_hd__a2bb2o_4
X_19784_ _19784_/A VGND VGND VPWR VPWR _19784_/X sky130_fd_sc_hd__buf_2
XFILLER_205_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24664__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_85_0_HCLK clkbuf_8_85_0_HCLK/A VGND VGND VPWR VPWR _25346_/CLK sky130_fd_sc_hd__clkbuf_1
X_15947_ _12245_/Y _15944_/X _15946_/X _15944_/X VGND VGND VPWR VPWR _24768_/D sky130_fd_sc_hd__a2bb2o_4
X_18735_ _18735_/A VGND VGND VPWR VPWR _18735_/X sky130_fd_sc_hd__buf_2
XFILLER_237_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18666_ _16550_/A _18707_/B _16610_/Y _24130_/Q VGND VGND VPWR VPWR _18668_/C sky130_fd_sc_hd__a2bb2o_4
X_15878_ _12780_/Y _15875_/X _11721_/X _15875_/X VGND VGND VPWR VPWR _15878_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14829_ _14812_/C _14797_/X _14812_/C _14797_/X VGND VGND VPWR VPWR _14829_/X sky130_fd_sc_hd__a2bb2o_4
X_17617_ _17564_/Y _17616_/X _17593_/X VGND VGND VPWR VPWR _17617_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_52_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18597_ _18477_/D _18498_/X _18500_/X _18595_/B VGND VGND VPWR VPWR _18598_/A sky130_fd_sc_hd__a211o_4
XFILLER_224_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22875__A1_N _17179_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17548_ _11777_/Y _24294_/Q _25521_/Q _17580_/C VGND VGND VPWR VPWR _17553_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17479_ _17473_/Y _17448_/A _17479_/C VGND VGND VPWR VPWR _18356_/B sky130_fd_sc_hd__and3_4
XFILLER_32_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11711__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19218_ _19218_/A VGND VGND VPWR VPWR _19218_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14376__B1 _13826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20490_ _20485_/X _20490_/B VGND VGND VPWR VPWR _20490_/X sky130_fd_sc_hd__or2_4
XANTENNA__25452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19149_ _19149_/A VGND VGND VPWR VPWR _19149_/X sky130_fd_sc_hd__buf_2
XANTENNA__22942__C _22941_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21110__A1 _24716_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22160_ _24452_/Q _21309_/X _22891_/A VGND VGND VPWR VPWR _22160_/X sky130_fd_sc_hd__o21a_4
XFILLER_246_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21111_ _21111_/A VGND VGND VPWR VPWR _21111_/X sky130_fd_sc_hd__buf_2
XFILLER_160_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14679__B2 _14678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15876__B1 _11715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22091_ _15121_/A _23088_/B VGND VGND VPWR VPWR _22095_/B sky130_fd_sc_hd__or2_4
XFILLER_172_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21042_ _16268_/A _21089_/B VGND VGND VPWR VPWR _21042_/X sky130_fd_sc_hd__and2_4
XFILLER_141_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16891__A2_N _24283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15853__A _22638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21574__B _21574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24801_ _24819_/CLK _15882_/X HRESETn VGND VGND VPWR VPWR _24801_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22993_ _20781_/Y _22992_/X _20920_/Y _21227_/X VGND VGND VPWR VPWR _22993_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24334__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24732_ _24365_/CLK _24732_/D HRESETn VGND VGND VPWR VPWR _16031_/A sky130_fd_sc_hd__dfrtp_4
X_21944_ _21466_/A _21944_/B VGND VGND VPWR VPWR _21944_/X sky130_fd_sc_hd__or2_4
XFILLER_216_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16053__B1 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22686__A _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21590__A _22829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24663_ _24662_/CLK _16224_/X HRESETn VGND VGND VPWR VPWR _22806_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_231_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21875_ _16154_/Y _21030_/A _22654_/B _11772_/Y _21581_/X VGND VGND VPWR VPWR _21875_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_131_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15800__B1 _11688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23627_/CLK _23614_/D VGND VGND VPWR VPWR _13350_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_242_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _20823_/A _20826_/B VGND VGND VPWR VPWR _20827_/A sky130_fd_sc_hd__or2_4
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24594_ _24594_/CLK _24594_/D HRESETn VGND VGND VPWR VPWR _22701_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23545_ _23526_/CLK _19994_/X VGND VGND VPWR VPWR _23545_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20757_ _20784_/A VGND VGND VPWR VPWR _20757_/X sky130_fd_sc_hd__buf_2
XANTENNA__23013__C _22817_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20688_ _20685_/A _20688_/B VGND VGND VPWR VPWR _20716_/A sky130_fd_sc_hd__or2_4
X_23476_ _23476_/CLK _23476_/D VGND VGND VPWR VPWR _20173_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12917__A1 _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25215_ _25224_/CLK _25215_/D HRESETn VGND VGND VPWR VPWR _14088_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_149_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22427_ _22394_/X _22409_/X _22427_/C _22427_/D VGND VGND VPWR VPWR HRDATA[7] sky130_fd_sc_hd__or4_4
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25122__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13160_ _13179_/A _13158_/X _13159_/X VGND VGND VPWR VPWR _13160_/X sky130_fd_sc_hd__and3_4
X_25146_ _25146_/CLK _14393_/X HRESETn VGND VGND VPWR VPWR _20606_/A sky130_fd_sc_hd__dfrtp_4
X_22358_ _21466_/A _22358_/B VGND VGND VPWR VPWR _22358_/X sky130_fd_sc_hd__or2_4
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15867__B1 _24811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12111_ _25469_/Q VGND VGND VPWR VPWR _12111_/Y sky130_fd_sc_hd__inv_2
X_13091_ _13091_/A _13090_/X _13091_/C VGND VGND VPWR VPWR _25340_/D sky130_fd_sc_hd__and3_4
X_21309_ _21309_/A VGND VGND VPWR VPWR _21309_/X sky130_fd_sc_hd__buf_2
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19058__B1 _19057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22289_ _16701_/Y _22416_/B VGND VGND VPWR VPWR _22289_/X sky130_fd_sc_hd__and2_4
X_25077_ _23889_/CLK _14633_/X HRESETn VGND VGND VPWR VPWR _14628_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12042_ _11668_/B VGND VGND VPWR VPWR _12160_/C sky130_fd_sc_hd__buf_2
X_24028_ _24060_/CLK _20799_/X HRESETn VGND VGND VPWR VPWR _20796_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15882__A3 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16850_ _14932_/Y _16845_/X _16849_/X _16845_/X VGND VGND VPWR VPWR _16850_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15801_ _15777_/X _15789_/X _15725_/X _24843_/Q _15787_/X VGND VGND VPWR VPWR _15801_/X
+ sky130_fd_sc_hd__a32o_4
X_16781_ _16781_/A VGND VGND VPWR VPWR _16781_/Y sky130_fd_sc_hd__inv_2
X_13993_ _13986_/X _13987_/X _14019_/C _14019_/D VGND VGND VPWR VPWR _13994_/A sky130_fd_sc_hd__or4_4
XANTENNA__24075__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18520_ _18480_/X _18498_/X _18510_/C VGND VGND VPWR VPWR _18520_/X sky130_fd_sc_hd__o21a_4
X_15732_ _12521_/Y _15728_/X _11715_/X _15731_/X VGND VGND VPWR VPWR _24874_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_218_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12944_ _12952_/A _12944_/B _12944_/C VGND VGND VPWR VPWR _12944_/X sky130_fd_sc_hd__and3_4
XFILLER_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24004__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18451_ _18451_/A _18448_/X _18449_/X _18451_/D VGND VGND VPWR VPWR _18452_/D sky130_fd_sc_hd__or4_4
X_15663_ _15663_/A VGND VGND VPWR VPWR _15663_/X sky130_fd_sc_hd__buf_2
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19781__B2 _19764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12875_ _12796_/Y _12875_/B VGND VGND VPWR VPWR _12885_/B sky130_fd_sc_hd__or2_4
XPHY_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16594__A _24525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17402_ _17384_/X _17398_/X _24339_/Q _21002_/A _17401_/X VGND VGND VPWR VPWR _17402_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14613_/X VGND VGND VPWR VPWR _14614_/Y sky130_fd_sc_hd__inv_2
XPHY_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11826_/A VGND VGND VPWR VPWR _11826_/Y sky130_fd_sc_hd__inv_2
X_18382_ _18381_/Y _18379_/X _24194_/Q _18379_/X VGND VGND VPWR VPWR _24195_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22668__A1 _12418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15593_/Y _15589_/X _11726_/X _15589_/X VGND VGND VPWR VPWR _15594_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17333_/A _17244_/X VGND VGND VPWR VPWR _17333_/X sky130_fd_sc_hd__or2_4
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14544_/X VGND VGND VPWR VPWR _14566_/D sky130_fd_sc_hd__inv_2
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ HWDATA[8] VGND VGND VPWR VPWR _11757_/X sky130_fd_sc_hd__buf_2
XFILLER_159_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12627__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21340__A1 _16534_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17264_ _17343_/B _17228_/X VGND VGND VPWR VPWR _17264_/X sky130_fd_sc_hd__and2_4
X_14476_ _14474_/Y _14475_/X _14384_/X _14475_/X VGND VGND VPWR VPWR _14476_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11688_ HWDATA[24] VGND VGND VPWR VPWR _11688_/X sky130_fd_sc_hd__buf_2
XFILLER_201_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19003_ _19002_/X VGND VGND VPWR VPWR _19011_/A sky130_fd_sc_hd__inv_2
X_16215_ _16190_/X VGND VGND VPWR VPWR _16215_/X sky130_fd_sc_hd__buf_2
XFILLER_174_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13427_ _13285_/A _13427_/B VGND VGND VPWR VPWR _13427_/X sky130_fd_sc_hd__or2_4
X_17195_ _24621_/Q _24350_/Q _16336_/Y _17358_/A VGND VGND VPWR VPWR _17198_/C sky130_fd_sc_hd__o22a_4
XANTENNA__23093__B2 _22846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16146_ _16144_/Y _16142_/X _16145_/X _16142_/X VGND VGND VPWR VPWR _24689_/D sky130_fd_sc_hd__a2bb2o_4
X_13358_ _13390_/A _13356_/X _13357_/X VGND VGND VPWR VPWR _13362_/B sky130_fd_sc_hd__and3_4
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12309_ _12309_/A VGND VGND VPWR VPWR _12309_/Y sky130_fd_sc_hd__inv_2
X_16077_ _16077_/A _15773_/B VGND VGND VPWR VPWR _16077_/X sky130_fd_sc_hd__or2_4
X_13289_ _13289_/A VGND VGND VPWR VPWR _13391_/A sky130_fd_sc_hd__buf_2
XFILLER_142_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24845__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15028_ _15028_/A _15021_/X _15024_/X _15027_/X VGND VGND VPWR VPWR _15028_/X sky130_fd_sc_hd__or4_4
X_19905_ _19900_/A VGND VGND VPWR VPWR _19905_/X sky130_fd_sc_hd__buf_2
X_19836_ _19831_/Y _19835_/X _19807_/X _19835_/X VGND VGND VPWR VPWR _23602_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16999__A1_N _16035_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19767_ _22224_/B _19764_/X _16864_/X _19764_/X VGND VGND VPWR VPWR _23625_/D sky130_fd_sc_hd__a2bb2o_4
X_16979_ _24745_/Q _16978_/A _15995_/Y _16978_/Y VGND VGND VPWR VPWR _16979_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18984__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11706__A _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18718_ _18718_/A VGND VGND VPWR VPWR _24154_/D sky130_fd_sc_hd__inv_2
X_19698_ _13273_/B VGND VGND VPWR VPWR _19698_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18649_ _24149_/Q VGND VGND VPWR VPWR _18739_/A sky130_fd_sc_hd__buf_2
XFILLER_213_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22659__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21660_ _21656_/X _21659_/X _17725_/X VGND VGND VPWR VPWR _21668_/B sky130_fd_sc_hd__o21a_4
XFILLER_101_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22659__B2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20611_ _20611_/A _20505_/X VGND VGND VPWR VPWR _23960_/D sky130_fd_sc_hd__and2_4
X_21591_ _16711_/Y _21745_/B VGND VGND VPWR VPWR _21591_/X sky130_fd_sc_hd__and2_4
XANTENNA__21331__A1 _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16937__A1_N _16154_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20542_ _18886_/X VGND VGND VPWR VPWR _20543_/A sky130_fd_sc_hd__inv_2
X_23330_ _24578_/Q _23172_/X _21339_/X VGND VGND VPWR VPWR _23330_/X sky130_fd_sc_hd__o21a_4
XFILLER_178_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20473_ _20450_/X _20611_/A _14530_/A _20435_/X VGND VGND VPWR VPWR _24082_/D sky130_fd_sc_hd__a211o_4
X_23261_ _23261_/A VGND VGND VPWR VPWR _23261_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15848__A _22816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19288__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14752__A _22202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23084__B2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25000_ _24133_/CLK _15338_/X HRESETn VGND VGND VPWR VPWR _25000_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22212_ _22212_/A _22208_/X _22211_/X VGND VGND VPWR VPWR _22213_/C sky130_fd_sc_hd__or3_4
XFILLER_180_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21095__B1 _21864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23192_ _23192_/A VGND VGND VPWR VPWR _23192_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22143_ _23138_/A VGND VGND VPWR VPWR _22282_/A sky130_fd_sc_hd__buf_2
XFILLER_105_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25200__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24586__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22074_ _22068_/X _22073_/X _14666_/X VGND VGND VPWR VPWR _22074_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__14521__B1 _23393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22595__B1 _24866_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24515__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21025_ _21024_/X VGND VGND VPWR VPWR _22466_/A sky130_fd_sc_hd__buf_2
XFILLER_113_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_1_0_HCLK_A clkbuf_3_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19212__B1 _19144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22976_ _23043_/A _22976_/B VGND VGND VPWR VPWR _22983_/C sky130_fd_sc_hd__and2_4
XFILLER_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16026__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24715_ _24645_/CLK _16076_/X HRESETn VGND VGND VPWR VPWR _21066_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21927_ _21933_/A _21927_/B _21927_/C VGND VGND VPWR VPWR _21927_/X sky130_fd_sc_hd__and3_4
XFILLER_215_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12660_ _12655_/A _12655_/B _12627_/X _12657_/B VGND VGND VPWR VPWR _12661_/A sky130_fd_sc_hd__a211o_4
X_24646_ _24903_/CLK _16269_/X HRESETn VGND VGND VPWR VPWR _21013_/A sky130_fd_sc_hd__dfrtp_4
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _24720_/Q _21336_/X _21118_/X _21857_/X VGND VGND VPWR VPWR _21859_/C sky130_fd_sc_hd__a211o_4
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25374__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _13125_/B VGND VGND VPWR VPWR _20810_/A sky130_fd_sc_hd__inv_2
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12680_/A VGND VGND VPWR VPWR _12648_/A sky130_fd_sc_hd__buf_2
X_24577_ _24080_/CLK _24577_/D HRESETn VGND VGND VPWR VPWR _16456_/A sky130_fd_sc_hd__dfrtp_4
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21789_ _21789_/A VGND VGND VPWR VPWR _21789_/Y sky130_fd_sc_hd__inv_2
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _14329_/X VGND VGND VPWR VPWR _14330_/Y sky130_fd_sc_hd__inv_2
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23528_ _23528_/CLK _20040_/X VGND VGND VPWR VPWR _20038_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20664__A _20664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23040__A _22638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14261_ _25186_/Q VGND VGND VPWR VPWR _14261_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23459_ _24252_/CLK _20218_/X VGND VGND VPWR VPWR _18203_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16000_ _24744_/Q VGND VGND VPWR VPWR _16000_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13212_ _13334_/A _23921_/Q VGND VGND VPWR VPWR _13212_/X sky130_fd_sc_hd__or2_4
XANTENNA__22822__A1 _24733_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14192_ _20516_/A VGND VGND VPWR VPWR _20510_/A sky130_fd_sc_hd__inv_2
XFILLER_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13143_ _13247_/A VGND VGND VPWR VPWR _13288_/A sky130_fd_sc_hd__inv_2
X_25129_ _25117_/CLK _25129_/D HRESETn VGND VGND VPWR VPWR _14083_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_124_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13074_ _13074_/A _13074_/B VGND VGND VPWR VPWR _13074_/X sky130_fd_sc_hd__or2_4
X_17951_ _17940_/A _17951_/B VGND VGND VPWR VPWR _17951_/X sky130_fd_sc_hd__or2_4
XFILLER_152_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24256__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12025_ _12024_/Y _12020_/X _25490_/Q _12020_/X VGND VGND VPWR VPWR _25491_/D sky130_fd_sc_hd__a2bb2o_4
X_16902_ _24276_/Q VGND VGND VPWR VPWR _17761_/A sky130_fd_sc_hd__inv_2
X_17882_ _17752_/A _17885_/B _16952_/X VGND VGND VPWR VPWR _17882_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA_clkbuf_5_30_0_HCLK_A clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19621_ _21496_/B _19616_/X _19620_/X _19616_/X VGND VGND VPWR VPWR _23676_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16833_ _24425_/Q VGND VGND VPWR VPWR _16833_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16764_ _16763_/Y _16760_/X _15746_/X _16760_/X VGND VGND VPWR VPWR _24458_/D sky130_fd_sc_hd__a2bb2o_4
X_19552_ _19552_/A VGND VGND VPWR VPWR _22238_/B sky130_fd_sc_hd__inv_2
XFILLER_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13976_ _25242_/Q VGND VGND VPWR VPWR _14001_/A sky130_fd_sc_hd__buf_2
XFILLER_247_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16017__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15715_ _12534_/Y _15714_/X _15557_/X _15714_/X VGND VGND VPWR VPWR _15715_/X sky130_fd_sc_hd__a2bb2o_4
X_18503_ _18493_/B VGND VGND VPWR VPWR _18504_/B sky130_fd_sc_hd__inv_2
XFILLER_46_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12927_ _12967_/A VGND VGND VPWR VPWR _12952_/A sky130_fd_sc_hd__buf_2
X_16695_ _16694_/Y _16692_/X _16597_/X _16692_/X VGND VGND VPWR VPWR _16695_/X sky130_fd_sc_hd__a2bb2o_4
X_19483_ _22336_/B _19482_/X _11902_/X _19482_/X VGND VGND VPWR VPWR _23722_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_159_0_HCLK clkbuf_7_79_0_HCLK/X VGND VGND VPWR VPWR _23927_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_206_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15646_ _15671_/A _15771_/B VGND VGND VPWR VPWR _15646_/X sky130_fd_sc_hd__or2_4
X_18434_ _16232_/Y _24171_/Q _16232_/Y _24171_/Q VGND VGND VPWR VPWR _18438_/A sky130_fd_sc_hd__a2bb2o_4
X_12858_ _12860_/B VGND VGND VPWR VPWR _12859_/B sky130_fd_sc_hd__inv_2
XFILLER_179_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23302__A2 _22661_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11809_ _11810_/A _11808_/Y _11803_/Y _24230_/Q VGND VGND VPWR VPWR _11809_/X sky130_fd_sc_hd__a2bb2o_4
X_18365_ _18365_/A _18365_/B VGND VGND VPWR VPWR _18365_/Y sky130_fd_sc_hd__nor2_4
XFILLER_221_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15577_ _15574_/Y _15570_/X _11691_/X _15576_/X VGND VGND VPWR VPWR _24916_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21313__A1 _21305_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12789_ _22713_/A VGND VGND VPWR VPWR _12837_/B sky130_fd_sc_hd__inv_2
XANTENNA__25044__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21313__B2 _22523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17316_ _17251_/C _17314_/X _17315_/Y VGND VGND VPWR VPWR _17316_/X sky130_fd_sc_hd__o21a_4
X_14528_ _14528_/A VGND VGND VPWR VPWR _14528_/Y sky130_fd_sc_hd__inv_2
X_18296_ _18296_/A _18303_/B VGND VGND VPWR VPWR _18296_/X sky130_fd_sc_hd__and2_4
XFILLER_202_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17247_ _24356_/Q VGND VGND VPWR VPWR _17329_/A sky130_fd_sc_hd__inv_2
X_14459_ _25122_/Q VGND VGND VPWR VPWR _14459_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17178_ _17170_/X _17173_/X _17176_/X _17178_/D VGND VGND VPWR VPWR _17178_/X sky130_fd_sc_hd__or4_4
XANTENNA__23100__D _23099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16129_ _16124_/A VGND VGND VPWR VPWR _16129_/X sky130_fd_sc_hd__buf_2
XFILLER_115_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19690__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19819_ _19819_/A VGND VGND VPWR VPWR _21752_/B sky130_fd_sc_hd__inv_2
XFILLER_29_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22830_ _20902_/Y _22829_/X _20764_/C _22290_/A VGND VGND VPWR VPWR _22830_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19603__A _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23979__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16271__A3 _16267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_55_0_HCLK clkbuf_7_55_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16008__B1 _15567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22761_ _21879_/X VGND VGND VPWR VPWR _22761_/X sky130_fd_sc_hd__buf_2
XANTENNA__14747__A _14678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21552__B2 _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18219__A _18056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24500_ _24501_/CLK _16666_/X HRESETn VGND VGND VPWR VPWR _24500_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21712_ _17241_/Y _22543_/A _25371_/Q _21423_/A VGND VGND VPWR VPWR _21712_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_212_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25480_ _25479_/CLK _25480_/D HRESETn VGND VGND VPWR VPWR _12074_/A sky130_fd_sc_hd__dfrtp_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23955__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22692_ _12226_/X _22721_/A _17758_/Y _22691_/X VGND VGND VPWR VPWR _22692_/X sky130_fd_sc_hd__o22a_4
XFILLER_197_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ _25028_/CLK _24431_/D HRESETn VGND VGND VPWR VPWR _14936_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_240_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21643_ _21379_/B VGND VGND VPWR VPWR _21643_/X sky130_fd_sc_hd__buf_2
XFILLER_240_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22501__B1 _12772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22683__B _22730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24362_ _24341_/CLK _24362_/D HRESETn VGND VGND VPWR VPWR _17174_/A sky130_fd_sc_hd__dfrtp_4
X_21574_ _21568_/A _21574_/B VGND VGND VPWR VPWR _21575_/A sky130_fd_sc_hd__or2_4
XFILLER_165_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23313_ _23313_/A _21528_/B VGND VGND VPWR VPWR _23313_/X sky130_fd_sc_hd__or2_4
X_20525_ _23967_/Q _20525_/B _20525_/C _20524_/X VGND VGND VPWR VPWR _20526_/A sky130_fd_sc_hd__or4_4
X_24293_ _24947_/CLK _17697_/X HRESETn VGND VGND VPWR VPWR _17521_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_165_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24767__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20456_ _20454_/X _20455_/X VGND VGND VPWR VPWR _20456_/X sky130_fd_sc_hd__or2_4
X_23244_ _14962_/A _23138_/X _22801_/X _23243_/X VGND VGND VPWR VPWR _23245_/C sky130_fd_sc_hd__a211o_4
XFILLER_118_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20387_ _20387_/A _20387_/B _20387_/C VGND VGND VPWR VPWR _20387_/X sky130_fd_sc_hd__or3_4
X_23175_ _23209_/A _23170_/X _23174_/X VGND VGND VPWR VPWR _23175_/X sky130_fd_sc_hd__and3_4
XANTENNA__19681__B1 _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12513__A1_N _25411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22126_ _21345_/Y _22109_/X _22113_/Y _22118_/Y _22125_/X VGND VGND VPWR VPWR _22126_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_133_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22204__A _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22057_ _22385_/A _19812_/Y VGND VGND VPWR VPWR _22059_/B sky130_fd_sc_hd__or2_4
XFILLER_121_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21008_ _21008_/A VGND VGND VPWR VPWR _21010_/B sky130_fd_sc_hd__inv_2
XFILLER_208_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13830_ _13530_/Y _13828_/X _13829_/X _13828_/X VGND VGND VPWR VPWR _25260_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23035__A _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13761_ _13807_/B VGND VGND VPWR VPWR _16721_/B sky130_fd_sc_hd__buf_2
X_22959_ _23094_/A _22958_/X VGND VGND VPWR VPWR _22959_/Y sky130_fd_sc_hd__nor2_4
XFILLER_204_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13481__B1 _13459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15500_ _15498_/Y _15494_/X HADDR[17] _15499_/X VGND VGND VPWR VPWR _15500_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21543__B2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12712_ _25406_/Q _12711_/Y VGND VGND VPWR VPWR _12713_/B sky130_fd_sc_hd__or2_4
X_16480_ _16479_/Y _16475_/X _16391_/X _16475_/X VGND VGND VPWR VPWR _24569_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13692_ _11806_/A _13692_/B VGND VGND VPWR VPWR _13692_/X sky130_fd_sc_hd__or2_4
XFILLER_189_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15431_ _13927_/A _15427_/X _15430_/X VGND VGND VPWR VPWR _24975_/D sky130_fd_sc_hd__o21ai_4
X_12643_ _12505_/Y _12645_/B _12642_/Y VGND VGND VPWR VPWR _12643_/X sky130_fd_sc_hd__o21a_4
X_24629_ _24629_/CLK _16316_/X HRESETn VGND VGND VPWR VPWR _22821_/A sky130_fd_sc_hd__dfrtp_4
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22099__A2 _21064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16970__A1 _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18150_ _18118_/A _18150_/B VGND VGND VPWR VPWR _18152_/B sky130_fd_sc_hd__or2_4
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15362_ _15292_/A _15361_/X VGND VGND VPWR VPWR _15362_/Y sky130_fd_sc_hd__nand2_4
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _24877_/Q VGND VGND VPWR VPWR _12574_/Y sky130_fd_sc_hd__inv_2
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17101_ _16969_/Y _17099_/X _17100_/Y VGND VGND VPWR VPWR _17101_/X sky130_fd_sc_hd__o21a_4
XFILLER_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11795__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ _14318_/A _25170_/Q _25169_/Q VGND VGND VPWR VPWR _14313_/X sky130_fd_sc_hd__a21o_4
XFILLER_196_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18081_ _17947_/A _18072_/X _18080_/X VGND VGND VPWR VPWR _18081_/X sky130_fd_sc_hd__and3_4
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15293_ _15351_/A _15293_/B _15347_/A VGND VGND VPWR VPWR _15301_/A sky130_fd_sc_hd__or3_4
XFILLER_184_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12905__A _12838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14392__A _14392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16722__B2 _16721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17032_ _17032_/A _17004_/Y _17031_/X VGND VGND VPWR VPWR _17032_/X sky130_fd_sc_hd__or3_4
XFILLER_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14244_ _21155_/B VGND VGND VPWR VPWR _14245_/A sky130_fd_sc_hd__buf_2
XFILLER_137_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24437__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14175_ _14174_/Y VGND VGND VPWR VPWR _20496_/A sky130_fd_sc_hd__buf_2
XFILLER_180_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16486__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13126_ _13126_/A _13125_/X VGND VGND VPWR VPWR _20685_/B sky130_fd_sc_hd__or2_4
XFILLER_112_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18983_ _18983_/A VGND VGND VPWR VPWR _18983_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24090__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13057_ _13057_/A VGND VGND VPWR VPWR _25349_/D sky130_fd_sc_hd__inv_2
X_17934_ _17950_/A _17932_/X _17934_/C VGND VGND VPWR VPWR _17934_/X sky130_fd_sc_hd__and3_4
XFILLER_112_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19424__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23220__B2 _21871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12008_ _24098_/Q _12007_/A _12006_/Y _12007_/Y VGND VGND VPWR VPWR _12012_/C sky130_fd_sc_hd__o22a_4
XANTENNA__17419__A2_N _17414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17865_ _16915_/Y _17862_/X VGND VGND VPWR VPWR _17865_/X sky130_fd_sc_hd__or2_4
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19604_ _22240_/B _19599_/X _19603_/X _19599_/X VGND VGND VPWR VPWR _23681_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15951__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16816_ _16799_/A VGND VGND VPWR VPWR _16816_/X sky130_fd_sc_hd__buf_2
XFILLER_94_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17796_ _17764_/A _17795_/X VGND VGND VPWR VPWR _17796_/X sky130_fd_sc_hd__or2_4
XFILLER_93_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19535_ _21960_/A _19531_/X _19534_/X _19531_/X VGND VGND VPWR VPWR _23703_/D sky130_fd_sc_hd__a2bb2o_4
X_13959_ _13929_/Y _13939_/B _13958_/X _13952_/B VGND VGND VPWR VPWR _13959_/X sky130_fd_sc_hd__or4_4
X_16747_ _15047_/Y _16745_/X _16395_/X _16745_/X VGND VGND VPWR VPWR _16747_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13472__B1 _11775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16678_ _16677_/Y _16673_/X _16320_/X _16673_/X VGND VGND VPWR VPWR _16678_/X sky130_fd_sc_hd__a2bb2o_4
X_19466_ _21947_/B _19463_/X _11915_/X _19463_/X VGND VGND VPWR VPWR _23727_/D sky130_fd_sc_hd__a2bb2o_4
X_18417_ _23248_/A _24187_/Q _16189_/Y _18416_/Y VGND VGND VPWR VPWR _18424_/A sky130_fd_sc_hd__o22a_4
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15629_ _21746_/A _15622_/X _15469_/X _15628_/X VGND VGND VPWR VPWR _24896_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19397_ _19394_/Y _19389_/X _19395_/X _19396_/X VGND VGND VPWR VPWR _19397_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12087__A _16181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16782__A HWDATA[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18348_ _13179_/A _18346_/X _18347_/Y VGND VGND VPWR VPWR _18348_/X sky130_fd_sc_hd__o21a_4
XFILLER_147_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21837__A2 _14212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18279_ _18279_/A VGND VGND VPWR VPWR _18279_/X sky130_fd_sc_hd__buf_2
XFILLER_175_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20310_ _20309_/X VGND VGND VPWR VPWR _20310_/X sky130_fd_sc_hd__buf_2
XANTENNA__24860__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21290_ _21290_/A VGND VGND VPWR VPWR _21592_/A sky130_fd_sc_hd__buf_2
XFILLER_163_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24178__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20241_ _20157_/C _13744_/X _13743_/X _14683_/X VGND VGND VPWR VPWR _20242_/A sky130_fd_sc_hd__or4_4
XANTENNA__21847__B _22119_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24107__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20172_ _21630_/B _20171_/X _20106_/X _20171_/X VGND VGND VPWR VPWR _23477_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15819__A3 _16240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19415__B1 _19414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24980_ _24980_/CLK _24980_/D HRESETn VGND VGND VPWR VPWR _24980_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16022__A _24736_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23931_ _23932_/CLK _23931_/D HRESETn VGND VGND VPWR VPWR _23931_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21863__A _21127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23862_ _23806_/CLK _19084_/X VGND VGND VPWR VPWR _23862_/Q sky130_fd_sc_hd__dfxtp_4
X_22813_ _16444_/X VGND VGND VPWR VPWR _23251_/A sky130_fd_sc_hd__buf_2
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23793_ _23754_/CLK _23793_/D VGND VGND VPWR VPWR _23793_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_226_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17729__B1 _17725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22722__B1 _24834_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25532_ _25533_/CLK _11745_/X HRESETn VGND VGND VPWR VPWR _25532_/Q sky130_fd_sc_hd__dfrtp_4
X_22744_ _22629_/A _22744_/B _22743_/X VGND VGND VPWR VPWR _22766_/C sky130_fd_sc_hd__and3_4
XFILLER_198_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16401__B1 _16400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_142_0_HCLK clkbuf_7_71_0_HCLK/X VGND VGND VPWR VPWR _23735_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25463_ _25382_/CLK _12384_/Y HRESETn VGND VGND VPWR VPWR _25463_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_197_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22675_ _22450_/X _22672_/X _22454_/X _22674_/X VGND VGND VPWR VPWR _22676_/A sky130_fd_sc_hd__o22a_4
XFILLER_241_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24414_ _24477_/CLK _16853_/X HRESETn VGND VGND VPWR VPWR _16852_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_240_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24948__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21626_ _21769_/A _21623_/X _21625_/X VGND VGND VPWR VPWR _21626_/X sky130_fd_sc_hd__and3_4
XFILLER_197_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25394_ _25397_/CLK _25394_/D HRESETn VGND VGND VPWR VPWR _25394_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_178_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24345_ _24346_/CLK _24345_/D HRESETn VGND VGND VPWR VPWR _21856_/A sky130_fd_sc_hd__dfrtp_4
X_21557_ _21557_/A _21721_/B VGND VGND VPWR VPWR _21557_/Y sky130_fd_sc_hd__nor2_4
X_20508_ _24001_/Q _20448_/X _20507_/X VGND VGND VPWR VPWR _20508_/X sky130_fd_sc_hd__a21o_4
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12290_ _12290_/A VGND VGND VPWR VPWR _12291_/A sky130_fd_sc_hd__inv_2
X_24276_ _25450_/CLK _24276_/D HRESETn VGND VGND VPWR VPWR _24276_/Q sky130_fd_sc_hd__dfrtp_4
X_21488_ _21484_/X _21488_/B _21488_/C VGND VGND VPWR VPWR _21488_/X sky130_fd_sc_hd__and3_4
XANTENNA__24530__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23227_ _23108_/X _23224_/Y _23155_/X _23226_/X VGND VGND VPWR VPWR _23228_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_181_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20439_ _20438_/X VGND VGND VPWR VPWR _20439_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14940__A _14940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16468__B1 _16467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23158_ _22908_/X _23157_/X _23050_/X _25546_/Q _22910_/X VGND VGND VPWR VPWR _23158_/X
+ sky130_fd_sc_hd__a32o_4
X_22109_ _22109_/A _22109_/B _22109_/C _22108_/X VGND VGND VPWR VPWR _22109_/X sky130_fd_sc_hd__or4_4
X_15980_ _15980_/A VGND VGND VPWR VPWR _15980_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19406__B1 _19360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23089_ _15037_/A _23263_/B _23263_/C VGND VGND VPWR VPWR _23089_/X sky130_fd_sc_hd__and3_4
XANTENNA__22869__A _22145_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14931_ _25010_/Q VGND VGND VPWR VPWR _15273_/A sky130_fd_sc_hd__inv_2
XFILLER_94_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22556__A3 _22135_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21773__A _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22961__B1 _11710_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14862_ _14806_/X _14861_/Y _15468_/A _14806_/X VGND VGND VPWR VPWR _25044_/D sky130_fd_sc_hd__a2bb2o_4
X_17650_ _17638_/B VGND VGND VPWR VPWR _17651_/B sky130_fd_sc_hd__inv_2
XFILLER_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15443__A1 _14269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13813_ _13810_/A VGND VGND VPWR VPWR _13813_/X sky130_fd_sc_hd__buf_2
X_16601_ HWDATA[8] VGND VGND VPWR VPWR _16601_/X sky130_fd_sc_hd__buf_2
XFILLER_217_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17581_ _17581_/A _17581_/B _17581_/C VGND VGND VPWR VPWR _17581_/X sky130_fd_sc_hd__or3_4
XFILLER_235_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14793_ _14859_/A _14859_/B _14859_/C _25044_/Q VGND VGND VPWR VPWR _14808_/B sky130_fd_sc_hd__or4_4
X_16532_ _24549_/Q VGND VGND VPWR VPWR _16532_/Y sky130_fd_sc_hd__inv_2
X_19320_ _19320_/A _13596_/A _19320_/C VGND VGND VPWR VPWR _19321_/A sky130_fd_sc_hd__or3_4
X_13744_ _13739_/Y VGND VGND VPWR VPWR _13744_/X sky130_fd_sc_hd__buf_2
XFILLER_44_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12619__B _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16463_ _24575_/Q VGND VGND VPWR VPWR _16463_/Y sky130_fd_sc_hd__inv_2
X_19251_ _23802_/Q VGND VGND VPWR VPWR _19251_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13675_ _11832_/Y _13675_/B VGND VGND VPWR VPWR _13676_/B sky130_fd_sc_hd__or2_4
XFILLER_232_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23269__B2 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16943__B2 _17880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15414_ _15296_/B _15418_/A VGND VGND VPWR VPWR _15415_/B sky130_fd_sc_hd__nand2_4
X_18202_ _17985_/X _18202_/B VGND VGND VPWR VPWR _18202_/X sky130_fd_sc_hd__or2_4
XANTENNA__24689__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12626_ _12512_/Y _12608_/X _12503_/Y _12626_/D VGND VGND VPWR VPWR _12626_/X sky130_fd_sc_hd__or4_4
X_19182_ _19181_/Y _19177_/X _19138_/X _19170_/A VGND VGND VPWR VPWR _23827_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16394_ _15084_/Y _16393_/X _16020_/X _16393_/X VGND VGND VPWR VPWR _24601_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18133_ _15691_/X _18117_/X _18132_/X _24246_/Q _18022_/X VGND VGND VPWR VPWR _18133_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24618__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15345_ _15281_/A VGND VGND VPWR VPWR _15352_/A sky130_fd_sc_hd__buf_2
X_12557_ _12549_/X _12557_/B _12557_/C _12556_/X VGND VGND VPWR VPWR _12587_/A sky130_fd_sc_hd__or4_4
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18064_ _17966_/X _18063_/X _24247_/Q _18024_/X VGND VGND VPWR VPWR _18064_/X sky130_fd_sc_hd__o22a_4
X_15276_ _15273_/A _15273_/B VGND VGND VPWR VPWR _15276_/Y sky130_fd_sc_hd__nand2_4
XFILLER_156_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12488_ _12252_/X _12491_/B _12382_/X VGND VGND VPWR VPWR _12488_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_172_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17015_ _16987_/X _17014_/X VGND VGND VPWR VPWR _17343_/B sky130_fd_sc_hd__or2_4
XANTENNA__24271__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14227_ _25195_/Q VGND VGND VPWR VPWR _14227_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15946__A HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12193__B1 _12191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24200__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14158_ _25132_/Q VGND VGND VPWR VPWR _14158_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13109_ _13109_/A VGND VGND VPWR VPWR _13111_/A sky130_fd_sc_hd__inv_2
X_14089_ _14103_/C _14088_/X _14089_/C VGND VGND VPWR VPWR _14089_/X sky130_fd_sc_hd__or3_4
X_18966_ _14654_/A VGND VGND VPWR VPWR _18966_/X sky130_fd_sc_hd__buf_2
XANTENNA__25477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17917_ _15907_/Y _17917_/B VGND VGND VPWR VPWR _17917_/Y sky130_fd_sc_hd__nor2_4
X_18897_ _14425_/B _17438_/B VGND VGND VPWR VPWR _18897_/Y sky130_fd_sc_hd__nor2_4
XFILLER_39_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16777__A HWDATA[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17848_ _17810_/A VGND VGND VPWR VPWR _17866_/A sky130_fd_sc_hd__buf_2
XANTENNA__18620__B2 _18760_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17779_ _17779_/A VGND VGND VPWR VPWR _17780_/B sky130_fd_sc_hd__inv_2
XFILLER_82_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19518_ _21492_/B _19515_/X _11927_/X _19515_/X VGND VGND VPWR VPWR _19518_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25167__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20790_ _20789_/Y _20786_/Y _20793_/B VGND VGND VPWR VPWR _20790_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17187__A1 _24619_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19449_ _19449_/A VGND VGND VPWR VPWR _19449_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_215_0_HCLK clkbuf_8_214_0_HCLK/A VGND VGND VPWR VPWR _25021_/CLK sky130_fd_sc_hd__clkbuf_1
X_22460_ _21962_/A VGND VGND VPWR VPWR _22696_/B sky130_fd_sc_hd__buf_2
XFILLER_195_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24359__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21411_ _22197_/A _21411_/B VGND VGND VPWR VPWR _21411_/X sky130_fd_sc_hd__or2_4
XFILLER_194_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22391_ _22228_/A _22370_/Y _22377_/Y _22384_/Y _22390_/Y VGND VGND VPWR VPWR _22391_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24130_ _24139_/CLK _18814_/Y HRESETn VGND VGND VPWR VPWR _24130_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16698__B1 _16601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21342_ _21845_/A _21335_/X _21342_/C VGND VGND VPWR VPWR _21419_/B sky130_fd_sc_hd__and3_4
XFILLER_191_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18857__A1_N _16520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24061_ _24060_/CLK _24061_/D HRESETn VGND VGND VPWR VPWR _20941_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21273_ _14710_/A _21265_/X _21272_/X VGND VGND VPWR VPWR _21273_/X sky130_fd_sc_hd__or3_4
XFILLER_116_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18439__B2 _18400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23012_ _23012_/A _21058_/X VGND VGND VPWR VPWR _23015_/B sky130_fd_sc_hd__or2_4
XFILLER_116_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21443__B1 _24821_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20224_ _20224_/A VGND VGND VPWR VPWR _20224_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21296__C _15660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20155_ _21259_/B _20150_/X _20133_/X _20137_/Y VGND VGND VPWR VPWR _23483_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23994__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23923__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20086_ _20136_/A _13734_/X VGND VGND VPWR VPWR _20087_/A sky130_fd_sc_hd__and2_4
X_24963_ _24073_/CLK _24963_/D HRESETn VGND VGND VPWR VPWR _13935_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23914_ _23391_/CLK _23914_/D VGND VGND VPWR VPWR _23914_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19063__A _19063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24894_ _24035_/CLK _15633_/X HRESETn VGND VGND VPWR VPWR _24894_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_15_0_HCLK_A clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23845_ _23846_/CLK _19134_/X VGND VGND VPWR VPWR _23845_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_25_0_HCLK clkbuf_6_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _25520_/Q VGND VGND VPWR VPWR _11790_/Y sky130_fd_sc_hd__inv_2
X_23776_ _23827_/CLK _19328_/X VGND VGND VPWR VPWR _18048_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20988_ _20987_/A _14084_/Y _20987_/C VGND VGND VPWR VPWR _20988_/X sky130_fd_sc_hd__or3_4
XPHY_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22171__B2 _14209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15131__A2_N _24603_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25515_ _25499_/CLK _25515_/D HRESETn VGND VGND VPWR VPWR _25515_/Q sky130_fd_sc_hd__dfrtp_4
X_22727_ _22530_/A VGND VGND VPWR VPWR _22800_/B sky130_fd_sc_hd__buf_2
XFILLER_213_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24782__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13460_ _13452_/Y _13458_/Y _13459_/X _13458_/Y VGND VGND VPWR VPWR _25325_/D sky130_fd_sc_hd__a2bb2o_4
X_25446_ _25453_/CLK _25446_/D HRESETn VGND VGND VPWR VPWR _12229_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22658_ _24798_/Q _22658_/B VGND VGND VPWR VPWR _22658_/X sky130_fd_sc_hd__or2_4
XFILLER_230_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12411_ _12402_/X VGND VGND VPWR VPWR _12412_/B sky130_fd_sc_hd__inv_2
XANTENNA__24711__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21609_ _22221_/A VGND VGND VPWR VPWR _21609_/X sky130_fd_sc_hd__buf_2
X_13391_ _13391_/A _19226_/A VGND VGND VPWR VPWR _13393_/B sky130_fd_sc_hd__or2_4
X_25377_ _25373_/CLK _12944_/X HRESETn VGND VGND VPWR VPWR _12772_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19875__B1 _19874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22589_ _22588_/X VGND VGND VPWR VPWR _22614_/B sky130_fd_sc_hd__inv_2
XANTENNA__24029__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15130_ _24999_/Q VGND VGND VPWR VPWR _15130_/Y sky130_fd_sc_hd__inv_2
X_12342_ _12342_/A VGND VGND VPWR VPWR _13017_/A sky130_fd_sc_hd__inv_2
X_24328_ _24326_/CLK _17430_/X HRESETn VGND VGND VPWR VPWR _24328_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21768__A _22379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20672__A _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14164__A1 _14158_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15061_ _15061_/A _14944_/Y _15210_/A _15207_/A VGND VGND VPWR VPWR _15063_/C sky130_fd_sc_hd__or4_4
X_12273_ _12273_/A _12273_/B _12272_/Y _12248_/Y VGND VGND VPWR VPWR _12275_/C sky130_fd_sc_hd__or4_4
X_24259_ _24263_/CLK _24259_/D HRESETn VGND VGND VPWR VPWR _16923_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_181_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14670__A _21622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14012_ _14012_/A _13975_/A VGND VGND VPWR VPWR _14034_/C sky130_fd_sc_hd__or2_4
X_18820_ _18793_/A _18820_/B _18819_/Y VGND VGND VPWR VPWR _18820_/X sky130_fd_sc_hd__and3_4
XANTENNA__12190__A _25441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12621__C _12681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18751_ _18613_/X _18749_/A VGND VGND VPWR VPWR _18751_/X sky130_fd_sc_hd__or2_4
X_15963_ _15784_/X _15958_/X _16240_/A _22597_/A _15925_/X VGND VGND VPWR VPWR _15963_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_107_0_HCLK clkbuf_6_53_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_214_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16597__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17702_ _17701_/X VGND VGND VPWR VPWR _24291_/D sky130_fd_sc_hd__inv_2
XFILLER_76_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14914_ _24438_/Q VGND VGND VPWR VPWR _14914_/Y sky130_fd_sc_hd__inv_2
X_15894_ _12763_/Y _15892_/X _15616_/X _15892_/X VGND VGND VPWR VPWR _24792_/D sky130_fd_sc_hd__a2bb2o_4
X_18682_ _18679_/Y _18643_/A _18787_/A _18682_/D VGND VGND VPWR VPWR _18682_/X sky130_fd_sc_hd__or4_4
XFILLER_124_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17633_ _17502_/Y _17630_/X VGND VGND VPWR VPWR _17633_/X sky130_fd_sc_hd__or2_4
X_14845_ _14823_/X _14844_/X _25194_/Q _14830_/X VGND VGND VPWR VPWR _14845_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_90_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14776_ _14775_/Y _14776_/B VGND VGND VPWR VPWR _14777_/A sky130_fd_sc_hd__and2_4
X_17564_ _17564_/A VGND VGND VPWR VPWR _17564_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21950__B _21950_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11988_ _25311_/Q _11985_/X _11986_/Y _11987_/Y VGND VGND VPWR VPWR _11998_/A sky130_fd_sc_hd__o22a_4
X_19303_ _23785_/Q VGND VGND VPWR VPWR _19303_/Y sky130_fd_sc_hd__inv_2
X_13727_ _13727_/A VGND VGND VPWR VPWR _13730_/A sky130_fd_sc_hd__inv_2
X_16515_ _24555_/Q VGND VGND VPWR VPWR _16515_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17495_ _25526_/Q _17574_/D _17494_/Y _24110_/Q VGND VGND VPWR VPWR _17497_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16916__A1 _22494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19234_ _22365_/B _19233_/X _16860_/X _19233_/X VGND VGND VPWR VPWR _23810_/D sky130_fd_sc_hd__a2bb2o_4
X_13658_ _13658_/A VGND VGND VPWR VPWR _13658_/Y sky130_fd_sc_hd__inv_2
X_16446_ _13800_/B _21571_/A _16446_/C _16446_/D VGND VGND VPWR VPWR _16446_/X sky130_fd_sc_hd__or4_4
XFILLER_176_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24452__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12609_ _12512_/Y _12608_/X VGND VGND VPWR VPWR _12630_/B sky130_fd_sc_hd__or2_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16377_ _15104_/Y _16370_/X _15996_/X _16376_/X VGND VGND VPWR VPWR _16377_/X sky130_fd_sc_hd__a2bb2o_4
X_19165_ _19170_/A VGND VGND VPWR VPWR _19165_/X sky130_fd_sc_hd__buf_2
X_13589_ _25073_/Q VGND VGND VPWR VPWR _13596_/A sky130_fd_sc_hd__buf_2
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_45_0_HCLK clkbuf_8_45_0_HCLK/A VGND VGND VPWR VPWR _23425_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_173_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15328_ _15320_/B _15320_/D _15082_/Y VGND VGND VPWR VPWR _15328_/X sky130_fd_sc_hd__o21a_4
X_18116_ _18227_/A _18112_/X _18115_/X VGND VGND VPWR VPWR _18116_/X sky130_fd_sc_hd__or3_4
XFILLER_173_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19096_ _19101_/A VGND VGND VPWR VPWR _19096_/X sky130_fd_sc_hd__buf_2
XFILLER_145_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15259_ _15254_/A _15254_/B _15185_/A _15256_/B VGND VGND VPWR VPWR _15259_/X sky130_fd_sc_hd__a211o_4
X_18047_ _18085_/A _18045_/X _18047_/C VGND VGND VPWR VPWR _18047_/X sky130_fd_sc_hd__and3_4
XANTENNA__19618__B1 _19617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18052__A _18052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13196__A _13289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19998_ _19998_/A VGND VGND VPWR VPWR _19998_/Y sky130_fd_sc_hd__inv_2
X_18949_ _18946_/Y _18947_/X _18948_/X _18947_/X VGND VGND VPWR VPWR _18949_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21960_ _21960_/A _21960_/B VGND VGND VPWR VPWR _21960_/X sky130_fd_sc_hd__or2_4
XFILLER_67_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16604__B1 _16518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20911_ _20911_/A VGND VGND VPWR VPWR _20916_/B sky130_fd_sc_hd__inv_2
X_21891_ _21886_/X _21890_/X _22205_/A VGND VGND VPWR VPWR _21891_/X sky130_fd_sc_hd__o21a_4
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23630_ _23464_/CLK _19752_/X VGND VGND VPWR VPWR _23630_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20842_ _13644_/B VGND VGND VPWR VPWR _20842_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23561_ _25070_/CLK _19944_/X VGND VGND VPWR VPWR _19943_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20773_ _24022_/Q _20768_/X _20777_/B VGND VGND VPWR VPWR _20773_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_223_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16907__B2 _16906_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18227__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25300_ _23853_/CLK _25300_/D HRESETn VGND VGND VPWR VPWR _25300_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22512_ _20727_/Y _22992_/A _20866_/Y _22794_/A VGND VGND VPWR VPWR _22512_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22394__D _22393_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23492_ _23476_/CLK _23492_/D VGND VGND VPWR VPWR _23492_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24193__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25231_ _25230_/CLK _14075_/X HRESETn VGND VGND VPWR VPWR _13991_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22443_ _22781_/A _22443_/B _22443_/C _22442_/Y VGND VGND VPWR VPWR _22443_/X sky130_fd_sc_hd__or4_4
XFILLER_167_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25162_ _25164_/CLK _25162_/D HRESETn VGND VGND VPWR VPWR _12148_/C sky130_fd_sc_hd__dfrtp_4
X_22374_ _22378_/A _20407_/Y VGND VGND VPWR VPWR _22376_/B sky130_fd_sc_hd__or2_4
XFILLER_109_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24113_ _24626_/CLK _24113_/D HRESETn VGND VGND VPWR VPWR _24113_/Q sky130_fd_sc_hd__dfrtp_4
X_21325_ _11704_/A VGND VGND VPWR VPWR _21325_/X sky130_fd_sc_hd__buf_2
XFILLER_191_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25093_ _25089_/CLK _25093_/D HRESETn VGND VGND VPWR VPWR _25093_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12157__B1 SCLK_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25399__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24044_ _24487_/CLK _20869_/Y HRESETn VGND VGND VPWR VPWR _24044_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21256_ _22223_/A _21253_/X _21256_/C VGND VGND VPWR VPWR _21256_/X sky130_fd_sc_hd__and3_4
XFILLER_190_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21069__A1_N _21736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18897__A _14425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25328__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20207_ _20205_/Y _20201_/X _19746_/X _20206_/X VGND VGND VPWR VPWR _20207_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21187_ _21181_/X _21186_/X _17723_/A VGND VGND VPWR VPWR _21187_/X sky130_fd_sc_hd__o21a_4
XFILLER_78_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23953__D sda_i_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16843__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20138_ _20137_/Y VGND VGND VPWR VPWR _20138_/X sky130_fd_sc_hd__buf_2
XFILLER_237_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22212__A _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12960_ _12816_/Y _12963_/B _12854_/X VGND VGND VPWR VPWR _12960_/Y sky130_fd_sc_hd__a21oi_4
X_20069_ _23513_/Q VGND VGND VPWR VPWR _22203_/B sky130_fd_sc_hd__inv_2
X_24946_ _24357_/CLK _15491_/X HRESETn VGND VGND VPWR VPWR _15636_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11911_ _19606_/A VGND VGND VPWR VPWR _11911_/X sky130_fd_sc_hd__buf_2
XANTENNA__22392__B2 _22391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12891_ _12801_/X _12912_/A _12890_/X VGND VGND VPWR VPWR _12892_/B sky130_fd_sc_hd__or3_4
X_24877_ _24874_/CLK _15727_/X HRESETn VGND VGND VPWR VPWR _24877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_233_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14630_ _17950_/A _17943_/A _14630_/C _18009_/A VGND VGND VPWR VPWR _14630_/X sky130_fd_sc_hd__and4_4
XANTENNA__24963__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11842_ _11840_/A _11841_/A _13669_/A _11841_/Y VGND VGND VPWR VPWR _11842_/X sky130_fd_sc_hd__o22a_4
X_23828_ _23844_/CLK _23828_/D VGND VGND VPWR VPWR _23828_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14561_/A _14561_/B VGND VGND VPWR VPWR _14562_/A sky130_fd_sc_hd__or2_4
XPHY_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ HWDATA[4] VGND VGND VPWR VPWR _11774_/A sky130_fd_sc_hd__buf_2
X_23759_ _23767_/CLK _19375_/X VGND VGND VPWR VPWR _23759_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _14290_/A VGND VGND VPWR VPWR _13512_/Y sky130_fd_sc_hd__inv_2
X_16300_ _24635_/Q VGND VGND VPWR VPWR _16300_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _17280_/A VGND VGND VPWR VPWR _17280_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12788__A2_N _24797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _25112_/Q _14492_/B VGND VGND VPWR VPWR _14492_/Y sky130_fd_sc_hd__nor2_4
XPHY_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22882__A _23062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16231_ _16228_/Y _16223_/X _16229_/X _16230_/X VGND VGND VPWR VPWR _24661_/D sky130_fd_sc_hd__a2bb2o_4
X_13443_ _13443_/A _13443_/B VGND VGND VPWR VPWR _13443_/X sky130_fd_sc_hd__or2_4
X_25429_ _25428_/CLK _25429_/D HRESETn VGND VGND VPWR VPWR _25429_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_186_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15582__B1 _15581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17976__A _17999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_4_0_HCLK clkbuf_8_5_0_HCLK/A VGND VGND VPWR VPWR _25510_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_167_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16162_ _16161_/Y _16086_/A _15901_/X _16086_/A VGND VGND VPWR VPWR _16162_/X sky130_fd_sc_hd__a2bb2o_4
X_13374_ _13374_/A _23789_/Q VGND VGND VPWR VPWR _13376_/B sky130_fd_sc_hd__or2_4
XFILLER_6_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15113_ _24598_/Q VGND VGND VPWR VPWR _15113_/Y sky130_fd_sc_hd__inv_2
X_12325_ _24838_/Q VGND VGND VPWR VPWR _12325_/Y sky130_fd_sc_hd__inv_2
X_16093_ _16090_/Y _16086_/X _15996_/X _16092_/X VGND VGND VPWR VPWR _24710_/D sky130_fd_sc_hd__a2bb2o_4
X_15044_ _14883_/Y _24477_/Q _14883_/Y _24477_/Q VGND VGND VPWR VPWR _15049_/B sky130_fd_sc_hd__a2bb2o_4
X_19921_ _19918_/Y _19920_/X _19600_/X _19920_/X VGND VGND VPWR VPWR _19921_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21407__B1 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12256_ _12264_/A _12243_/Y _12266_/C _24752_/Q VGND VGND VPWR VPWR _12259_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25069__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19852_ _19852_/A VGND VGND VPWR VPWR _19852_/X sky130_fd_sc_hd__buf_2
XFILLER_96_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12187_ _12187_/A VGND VGND VPWR VPWR _12187_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18803_ _18803_/A VGND VGND VPWR VPWR _18803_/Y sky130_fd_sc_hd__inv_2
X_19783_ _19783_/A VGND VGND VPWR VPWR _19784_/A sky130_fd_sc_hd__inv_2
XFILLER_122_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16995_ _16995_/A _16995_/B _16993_/X _16995_/D VGND VGND VPWR VPWR _16995_/X sky130_fd_sc_hd__or4_4
XFILLER_95_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18734_ _18734_/A _18734_/B _18734_/C VGND VGND VPWR VPWR _24151_/D sky130_fd_sc_hd__and3_4
XFILLER_95_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15946_ HWDATA[20] VGND VGND VPWR VPWR _15946_/X sky130_fd_sc_hd__buf_2
X_18665_ _18665_/A VGND VGND VPWR VPWR _18707_/B sky130_fd_sc_hd__buf_2
X_15877_ _12753_/Y _15875_/X _11718_/X _15875_/X VGND VGND VPWR VPWR _15877_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17616_ _17511_/Y _17615_/X VGND VGND VPWR VPWR _17616_/X sky130_fd_sc_hd__or2_4
X_14828_ _23993_/D _14827_/X _20664_/A _23993_/D VGND VGND VPWR VPWR _14828_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_221_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18596_ _18592_/B _18596_/B _18593_/C VGND VGND VPWR VPWR _24159_/D sky130_fd_sc_hd__and3_4
XANTENNA__24633__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17547_ _17540_/X _17542_/X _17544_/X _17546_/X VGND VGND VPWR VPWR _17547_/X sky130_fd_sc_hd__or4_4
X_14759_ _14758_/X VGND VGND VPWR VPWR _16165_/B sky130_fd_sc_hd__inv_2
X_17478_ _21220_/A VGND VGND VPWR VPWR _17478_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19217_ _19215_/Y _19211_/X _19125_/X _19216_/X VGND VGND VPWR VPWR _23816_/D sky130_fd_sc_hd__a2bb2o_4
X_16429_ _24584_/Q VGND VGND VPWR VPWR _16429_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17886__A _17880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15573__B1 _11688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19148_ _19148_/A VGND VGND VPWR VPWR _19148_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21110__A2 _21098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19079_ _19074_/A VGND VGND VPWR VPWR _19079_/X sky130_fd_sc_hd__buf_2
XFILLER_161_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25492__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21110_ _24716_/Q _21098_/X _21099_/X _21109_/X VGND VGND VPWR VPWR _21110_/X sky130_fd_sc_hd__a211o_4
X_22090_ _21274_/X _22050_/Y _22055_/X _21510_/A _22089_/X VGND VGND VPWR VPWR _22090_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_160_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21041_ _15660_/A VGND VGND VPWR VPWR _21041_/X sky130_fd_sc_hd__buf_2
XANTENNA__19606__A _19606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22610__A2 _22435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18510__A _18560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16825__B1 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16537__A1_N _16536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24800_ _24800_/CLK _15883_/X HRESETn VGND VGND VPWR VPWR _24800_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22992_ _22992_/A VGND VGND VPWR VPWR _22992_/X sky130_fd_sc_hd__buf_2
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22967__A _21439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24731_ _24365_/CLK _16036_/X HRESETn VGND VGND VPWR VPWR _16035_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21871__A _23171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21943_ _17720_/A _19886_/Y VGND VGND VPWR VPWR _21945_/B sky130_fd_sc_hd__or2_4
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_5_7_0_HCLK_A clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24662_ _24662_/CLK _24662_/D HRESETn VGND VGND VPWR VPWR _22741_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21874_ _21101_/A VGND VGND VPWR VPWR _22654_/B sky130_fd_sc_hd__buf_2
XFILLER_27_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22126__A1 _21345_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14603__A2 _14610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23627_/CLK _23613_/D VGND VGND VPWR VPWR _13382_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__24374__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _20846_/A VGND VGND VPWR VPWR _20825_/X sky130_fd_sc_hd__buf_2
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24593_ _24592_/CLK _24593_/D HRESETn VGND VGND VPWR VPWR _24593_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_196_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13811__B1 _11730_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24303__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11902__A _19600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23544_ _23415_/CLK _23544_/D VGND VGND VPWR VPWR _23544_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20756_ _13121_/C _20750_/X _20755_/Y VGND VGND VPWR VPWR _20756_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__24109__D MSI_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23475_ _23499_/CLK _23475_/D VGND VGND VPWR VPWR _23475_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20687_ _20708_/A VGND VGND VPWR VPWR _20687_/X sky130_fd_sc_hd__buf_2
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25214_ _25211_/CLK _25214_/D HRESETn VGND VGND VPWR VPWR _14102_/C sky130_fd_sc_hd__dfrtp_4
X_22426_ _22286_/X _22419_/Y _22422_/X _22423_/X _22425_/X VGND VGND VPWR VPWR _22427_/D
+ sky130_fd_sc_hd__o32a_4
XFILLER_109_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22207__A _22199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25509__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25145_ _25113_/CLK _25145_/D HRESETn VGND VGND VPWR VPWR _25145_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__13829__A _13829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21111__A _21111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22357_ _21463_/A _22357_/B VGND VGND VPWR VPWR _22357_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_91_0_HCLK clkbuf_8_91_0_HCLK/A VGND VGND VPWR VPWR _25373_/CLK sky130_fd_sc_hd__clkbuf_1
X_12110_ _12154_/A _12107_/X _12076_/X _12107_/X VGND VGND VPWR VPWR _12110_/X sky130_fd_sc_hd__a2bb2o_4
X_21308_ _15851_/X VGND VGND VPWR VPWR _21309_/A sky130_fd_sc_hd__buf_2
XFILLER_152_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13090_ _25340_/Q _13090_/B VGND VGND VPWR VPWR _13090_/X sky130_fd_sc_hd__or2_4
X_25076_ _23890_/CLK _25076_/D HRESETn VGND VGND VPWR VPWR _18026_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_124_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22288_ _11704_/A VGND VGND VPWR VPWR _22416_/B sky130_fd_sc_hd__buf_2
XFILLER_105_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12041_ _12087_/B VGND VGND VPWR VPWR _12058_/B sky130_fd_sc_hd__buf_2
X_24027_ _24060_/CLK _20795_/X HRESETn VGND VGND VPWR VPWR _20793_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_105_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21239_ _21239_/A VGND VGND VPWR VPWR _21884_/A sky130_fd_sc_hd__buf_2
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15800_ _12309_/Y _15796_/X _11688_/X _15796_/X VGND VGND VPWR VPWR _24844_/D sky130_fd_sc_hd__a2bb2o_4
X_13992_ _13992_/A _13975_/A _14022_/B _14006_/A VGND VGND VPWR VPWR _14019_/D sky130_fd_sc_hd__or4_4
X_16780_ _15022_/Y _16774_/X _16778_/X _16779_/X VGND VGND VPWR VPWR _24450_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18569__B1 _18489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22877__A _16672_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12943_ _12834_/A _12941_/A VGND VGND VPWR VPWR _12944_/C sky130_fd_sc_hd__or2_4
X_15731_ _15713_/X VGND VGND VPWR VPWR _15731_/X sky130_fd_sc_hd__buf_2
XFILLER_246_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24929_ _25325_/CLK _15531_/X HRESETn VGND VGND VPWR VPWR _12043_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20376__B1 _19746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18450_ _16251_/Y _18395_/A _16259_/Y _24161_/Q VGND VGND VPWR VPWR _18451_/D sky130_fd_sc_hd__a2bb2o_4
X_12874_ _12804_/Y _12841_/D _12588_/X VGND VGND VPWR VPWR _12875_/B sky130_fd_sc_hd__or3_4
X_15662_ _15662_/A VGND VGND VPWR VPWR _15663_/A sky130_fd_sc_hd__buf_2
XPHY_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17401_/A VGND VGND VPWR VPWR _17401_/X sky130_fd_sc_hd__buf_2
XPHY_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11823_/A _24231_/Q _11823_/Y _11824_/Y VGND VGND VPWR VPWR _11825_/X sky130_fd_sc_hd__o22a_4
X_14613_ _25081_/Q _13623_/X _14612_/X VGND VGND VPWR VPWR _14613_/X sky130_fd_sc_hd__a21o_4
XFILLER_33_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ _15593_/A VGND VGND VPWR VPWR _15593_/Y sky130_fd_sc_hd__inv_2
X_18381_ _24195_/Q VGND VGND VPWR VPWR _18381_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22668__A2 _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12908__A _25385_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20679__A1 _20673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24044__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _13757_/Y _13577_/B VGND VGND VPWR VPWR _14544_/X sky130_fd_sc_hd__or2_4
X_17332_ _17331_/X VGND VGND VPWR VPWR _17332_/Y sky130_fd_sc_hd__inv_2
XFILLER_230_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21876__B1 _24824_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11766_/A VGND VGND VPWR VPWR _11756_/X sky130_fd_sc_hd__buf_2
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18611__A1_N _24525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21340__A2 _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _14468_/A VGND VGND VPWR VPWR _14475_/X sky130_fd_sc_hd__buf_2
X_17263_ _17230_/X _17263_/B _17262_/X VGND VGND VPWR VPWR _24372_/D sky130_fd_sc_hd__and3_4
XFILLER_197_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15555__B1 _15554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _11687_/A VGND VGND VPWR VPWR _11687_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19002_ _19117_/A _19002_/B _19163_/C VGND VGND VPWR VPWR _19002_/X sky130_fd_sc_hd__or3_4
XFILLER_146_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13426_ _13394_/A _13426_/B _13425_/X VGND VGND VPWR VPWR _13434_/B sky130_fd_sc_hd__or3_4
X_16214_ _22927_/A VGND VGND VPWR VPWR _16214_/Y sky130_fd_sc_hd__inv_2
X_17194_ _17193_/Y VGND VGND VPWR VPWR _17358_/A sky130_fd_sc_hd__buf_2
XFILLER_167_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23093__A2 _22718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16145_ HWDATA[8] VGND VGND VPWR VPWR _16145_/X sky130_fd_sc_hd__buf_2
X_13357_ _13389_/A _23853_/Q VGND VGND VPWR VPWR _13357_/X sky130_fd_sc_hd__or2_4
XFILLER_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12308_ _12308_/A VGND VGND VPWR VPWR _12308_/Y sky130_fd_sc_hd__inv_2
X_16076_ _11699_/X _21296_/A _15920_/X _21066_/A _16075_/X VGND VGND VPWR VPWR _16076_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_154_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_119_0_HCLK clkbuf_7_59_0_HCLK/X VGND VGND VPWR VPWR _25409_/CLK sky130_fd_sc_hd__clkbuf_1
X_13288_ _13288_/A VGND VGND VPWR VPWR _13393_/A sky130_fd_sc_hd__buf_2
XFILLER_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15027_ _25025_/Q _15025_/Y _15246_/C _15018_/A VGND VGND VPWR VPWR _15027_/X sky130_fd_sc_hd__a2bb2o_4
X_19904_ _19904_/A VGND VGND VPWR VPWR _22084_/B sky130_fd_sc_hd__inv_2
X_12239_ _12239_/A _12239_/B _12239_/C _12238_/X VGND VGND VPWR VPWR _12260_/B sky130_fd_sc_hd__or4_4
XFILLER_142_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24032__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16807__B1 _15721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19835_ _19835_/A VGND VGND VPWR VPWR _19835_/X sky130_fd_sc_hd__buf_2
XFILLER_84_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24885__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19766_ _19766_/A VGND VGND VPWR VPWR _22224_/B sky130_fd_sc_hd__inv_2
X_16978_ _16978_/A VGND VGND VPWR VPWR _16978_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22787__A _22730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18717_ _18707_/B _18707_/C _18709_/X _18714_/B VGND VGND VPWR VPWR _18718_/A sky130_fd_sc_hd__a211o_4
XANTENNA__24814__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15929_ _15923_/X _15928_/X _15710_/X _23275_/A _15926_/X VGND VGND VPWR VPWR _24778_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19697_ _19696_/Y _19694_/X _19630_/X _19694_/X VGND VGND VPWR VPWR _19697_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_232_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18648_ _16587_/Y _24139_/Q _16587_/Y _24139_/Q VGND VGND VPWR VPWR _18648_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22108__B2 _22119_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20382__A3 _13459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18579_ _18471_/D _18579_/B VGND VGND VPWR VPWR _18581_/B sky130_fd_sc_hd__nand2_4
XFILLER_224_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15794__B1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20610_ _20454_/X _20466_/X _20541_/B VGND VGND VPWR VPWR _23957_/D sky130_fd_sc_hd__o21a_4
XFILLER_221_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11722__A _11682_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21590_ _22829_/A VGND VGND VPWR VPWR _21597_/A sky130_fd_sc_hd__buf_2
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21331__A2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20541_ _14523_/A _20541_/B _14004_/X VGND VGND VPWR VPWR _23928_/D sky130_fd_sc_hd__and3_4
XFILLER_178_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23260_ _21421_/A _23258_/X _22831_/X _23259_/X VGND VGND VPWR VPWR _23261_/A sky130_fd_sc_hd__o22a_4
XFILLER_118_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20472_ _14375_/Y _14484_/X _20437_/C VGND VGND VPWR VPWR _20611_/A sky130_fd_sc_hd__a21o_4
XANTENNA__23084__A2 _21303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22211_ _22226_/A _22211_/B _22211_/C VGND VGND VPWR VPWR _22211_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_15_0_HCLK clkbuf_6_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__22292__B1 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23191_ _23044_/X _23190_/X _23046_/X _24743_/Q _23152_/X VGND VGND VPWR VPWR _23192_/A
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_7_78_0_HCLK clkbuf_7_79_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_78_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__21288__D _21287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22142_ _24346_/Q _22141_/X _23328_/A VGND VGND VPWR VPWR _22157_/A sky130_fd_sc_hd__a21o_4
XFILLER_161_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22073_ _22383_/A _22070_/X _22073_/C VGND VGND VPWR VPWR _22073_/X sky130_fd_sc_hd__and3_4
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21024_ _21151_/A _21568_/A _11668_/A _11676_/B VGND VGND VPWR VPWR _21024_/X sky130_fd_sc_hd__or4_4
XFILLER_102_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14199__B _14187_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24555__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22975_ _22971_/X _22972_/X _22973_/X _12514_/A _22974_/X VGND VGND VPWR VPWR _22976_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20358__B1 _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21926_ _21926_/A _20020_/Y VGND VGND VPWR VPWR _21927_/C sky130_fd_sc_hd__or2_4
X_24714_ _24645_/CLK _24714_/D HRESETn VGND VGND VPWR VPWR _24714_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21751__D _21750_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18971__B1 _18951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24645_ _24645_/CLK _24645_/D HRESETn VGND VGND VPWR VPWR _24645_/Q sky130_fd_sc_hd__dfrtp_4
X_21857_ _24616_/Q _21843_/B _21741_/B VGND VGND VPWR VPWR _21857_/X sky130_fd_sc_hd__and3_4
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _20807_/X VGND VGND VPWR VPWR _20808_/Y sky130_fd_sc_hd__inv_2
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12617_/B VGND VGND VPWR VPWR _12680_/A sky130_fd_sc_hd__buf_2
X_24576_ _24574_/CLK _24576_/D HRESETn VGND VGND VPWR VPWR _24576_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21788_ _21649_/X _21786_/X _21510_/A _21787_/X VGND VGND VPWR VPWR _21789_/A sky130_fd_sc_hd__a211o_4
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23527_ _23575_/CLK _20042_/X VGND VGND VPWR VPWR _20041_/A sky130_fd_sc_hd__dfxtp_4
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20739_ _20738_/Y _20732_/Y _13120_/B VGND VGND VPWR VPWR _20739_/X sky130_fd_sc_hd__o21a_4
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15001__A2 _24475_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _21557_/A _14259_/X _13791_/X _14259_/X VGND VGND VPWR VPWR _14260_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23458_ _23458_/CLK _23458_/D VGND VGND VPWR VPWR _23458_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25343__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13211_ _13289_/A VGND VGND VPWR VPWR _13334_/A sky130_fd_sc_hd__buf_2
XFILLER_109_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22409_ _21501_/X _18274_/A _22403_/X _22407_/X _22408_/X VGND VGND VPWR VPWR _22409_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_125_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14191_ _20496_/A _14188_/X _13824_/X _14190_/X VGND VGND VPWR VPWR _14191_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22283__B1 _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23389_ _23388_/CLK _23389_/D VGND VGND VPWR VPWR _13294_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__12771__B1 _12769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13142_ _13169_/A _13137_/X _13141_/X VGND VGND VPWR VPWR _13142_/X sky130_fd_sc_hd__and3_4
X_25128_ _23927_/CLK _25128_/D HRESETn VGND VGND VPWR VPWR _20539_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_136_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13073_ _13073_/A _13073_/B VGND VGND VPWR VPWR _13074_/B sky130_fd_sc_hd__or2_4
X_17950_ _17950_/A _17950_/B _17950_/C VGND VGND VPWR VPWR _17950_/X sky130_fd_sc_hd__and3_4
X_25059_ _23665_/CLK _25059_/D HRESETn VGND VGND VPWR VPWR _25059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12024_ _12024_/A VGND VGND VPWR VPWR _12024_/Y sky130_fd_sc_hd__inv_2
X_16901_ _16901_/A _16901_/B _16899_/X _16901_/D VGND VGND VPWR VPWR _16920_/B sky130_fd_sc_hd__or4_4
XANTENNA__22586__B2 _22992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17881_ _16917_/Y _17880_/X VGND VGND VPWR VPWR _17885_/B sky130_fd_sc_hd__or2_4
X_19620_ _19620_/A VGND VGND VPWR VPWR _19620_/X sky130_fd_sc_hd__buf_2
XFILLER_239_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16832_ _16831_/Y _16827_/X _15746_/X _16827_/X VGND VGND VPWR VPWR _16832_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24296__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19551_ _22353_/B _19550_/X _11902_/X _19550_/X VGND VGND VPWR VPWR _19551_/X sky130_fd_sc_hd__a2bb2o_4
X_16763_ _16763_/A VGND VGND VPWR VPWR _16763_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13975_ _13975_/A VGND VGND VPWR VPWR _13975_/Y sky130_fd_sc_hd__inv_2
X_18502_ _18502_/A VGND VGND VPWR VPWR _24186_/D sky130_fd_sc_hd__inv_2
XFILLER_206_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24225__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15714_ _15713_/X VGND VGND VPWR VPWR _15714_/X sky130_fd_sc_hd__buf_2
XFILLER_74_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12926_ _12926_/A VGND VGND VPWR VPWR _12926_/Y sky130_fd_sc_hd__inv_2
X_19482_ _19494_/A VGND VGND VPWR VPWR _19482_/X sky130_fd_sc_hd__buf_2
X_16694_ _16694_/A VGND VGND VPWR VPWR _16694_/Y sky130_fd_sc_hd__inv_2
X_18433_ _18433_/A _18433_/B _18431_/X _18432_/X VGND VGND VPWR VPWR _18452_/A sky130_fd_sc_hd__or4_4
XFILLER_179_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15645_ _16268_/A VGND VGND VPWR VPWR _15771_/B sky130_fd_sc_hd__buf_2
XFILLER_221_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12857_ _12857_/A _12857_/B VGND VGND VPWR VPWR _12860_/B sky130_fd_sc_hd__or2_4
XFILLER_206_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12638__A _12592_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11808_ _11808_/A VGND VGND VPWR VPWR _11808_/Y sky130_fd_sc_hd__inv_2
X_18364_ _18360_/Y _18363_/Y _18359_/X _18363_/A VGND VGND VPWR VPWR _18364_/X sky130_fd_sc_hd__o22a_4
X_12788_ _12920_/A _24797_/Q _12786_/Y _24797_/Q VGND VGND VPWR VPWR _12788_/X sky130_fd_sc_hd__a2bb2o_4
X_15576_ _15576_/A VGND VGND VPWR VPWR _15576_/X sky130_fd_sc_hd__buf_2
XANTENNA__24120__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17251_/C _17314_/X _17268_/X VGND VGND VPWR VPWR _17315_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_202_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11739_ _16233_/A VGND VGND VPWR VPWR _11739_/X sky130_fd_sc_hd__buf_2
X_14527_ _14030_/Y _14032_/Y _14527_/C _14003_/X VGND VGND VPWR VPWR _14528_/A sky130_fd_sc_hd__or4_4
X_18295_ _17707_/X _22261_/A VGND VGND VPWR VPWR _18303_/B sky130_fd_sc_hd__and2_4
XFILLER_159_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17246_ _24353_/Q VGND VGND VPWR VPWR _17246_/Y sky130_fd_sc_hd__inv_2
X_14458_ _14457_/Y _14455_/X _14262_/X _14455_/X VGND VGND VPWR VPWR _25123_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14200__B1 _13791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25084__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13409_ _13293_/A _13405_/X _13408_/X VGND VGND VPWR VPWR _13409_/X sky130_fd_sc_hd__or3_4
X_14389_ _16361_/A VGND VGND VPWR VPWR _14389_/X sky130_fd_sc_hd__buf_2
X_17177_ _16360_/Y _17239_/A _16360_/Y _17239_/A VGND VGND VPWR VPWR _17178_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12373__A _12204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25013__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16128_ _24695_/Q VGND VGND VPWR VPWR _16128_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16059_ _14403_/A VGND VGND VPWR VPWR _16059_/X sky130_fd_sc_hd__buf_2
XFILLER_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18060__A _18060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19818_ _19816_/Y _19814_/X _19817_/X _19814_/X VGND VGND VPWR VPWR _23607_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19749_ _19749_/A VGND VGND VPWR VPWR _19749_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17205__B1 _24617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22760_ _22759_/X VGND VGND VPWR VPWR _22760_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14747__B _14739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21552__A2 _14212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21711_ _12252_/X _21531_/X _24261_/Q _21431_/X VGND VGND VPWR VPWR _21711_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22691_ _22435_/A VGND VGND VPWR VPWR _22691_/X sky130_fd_sc_hd__buf_2
XANTENNA__15767__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24430_ _24462_/CLK _16823_/X HRESETn VGND VGND VPWR VPWR _16820_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_240_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21642_ _21642_/A VGND VGND VPWR VPWR _21642_/X sky130_fd_sc_hd__buf_2
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23948__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24361_ _24357_/CLK _24361_/D HRESETn VGND VGND VPWR VPWR _24361_/Q sky130_fd_sc_hd__dfrtp_4
X_21573_ _18385_/Y _21571_/X _12106_/Y _21570_/X VGND VGND VPWR VPWR _21573_/X sky130_fd_sc_hd__o22a_4
XFILLER_221_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14990__B2 _24474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23312_ _22716_/A _23312_/B VGND VGND VPWR VPWR _23319_/C sky130_fd_sc_hd__and2_4
X_20524_ _24076_/Q _20524_/B _24077_/Q VGND VGND VPWR VPWR _20524_/X sky130_fd_sc_hd__or3_4
X_24292_ _24305_/CLK _24292_/D HRESETn VGND VGND VPWR VPWR _17529_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16192__B1 _15996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23243_ _24474_/Q _22661_/X _23178_/X VGND VGND VPWR VPWR _23243_/X sky130_fd_sc_hd__o21a_4
XFILLER_107_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20455_ _20467_/A _20437_/A _20455_/C VGND VGND VPWR VPWR _20455_/X sky130_fd_sc_hd__and3_4
XFILLER_165_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22804__A2 _21871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21596__A _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23174_ _16554_/A _23171_/X _22928_/X _23173_/X VGND VGND VPWR VPWR _23174_/X sky130_fd_sc_hd__a211o_4
XFILLER_118_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20386_ _20386_/A VGND VGND VPWR VPWR _20386_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22125_ _22119_/X _22121_/Y _22123_/Y _22124_/X _21556_/Y VGND VGND VPWR VPWR _22125_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19066__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_102_0_HCLK clkbuf_7_51_0_HCLK/X VGND VGND VPWR VPWR _24623_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24736__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_165_0_HCLK clkbuf_7_82_0_HCLK/X VGND VGND VPWR VPWR _23884_/CLK sky130_fd_sc_hd__clkbuf_1
X_22056_ _22056_/A VGND VGND VPWR VPWR _22385_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_8_0_HCLK clkbuf_7_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21007_ _21007_/A VGND VGND VPWR VPWR _21007_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22220__A _22205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19197__B1 _19106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13760_ _13807_/A VGND VGND VPWR VPWR _16721_/A sky130_fd_sc_hd__buf_2
XFILLER_228_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17314__A _17179_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22958_ _12245_/Y _22718_/X _22719_/X _12354_/Y _22846_/X VGND VGND VPWR VPWR _22958_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_43_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12711_ _12711_/A VGND VGND VPWR VPWR _12711_/Y sky130_fd_sc_hd__inv_2
X_21909_ _21902_/A _20250_/Y VGND VGND VPWR VPWR _21909_/X sky130_fd_sc_hd__or2_4
X_13691_ _13686_/X _13667_/X _13689_/Y _13690_/X _11843_/A VGND VGND VPWR VPWR _13691_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15758__B1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22889_ _23176_/A VGND VGND VPWR VPWR _23005_/A sky130_fd_sc_hd__buf_2
XFILLER_71_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12642_ _12505_/Y _12645_/B _12641_/X VGND VGND VPWR VPWR _12642_/Y sky130_fd_sc_hd__a21oi_4
X_15430_ _15430_/A _15436_/B VGND VGND VPWR VPWR _15430_/X sky130_fd_sc_hd__or2_4
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24628_ _25521_/CLK _24628_/D HRESETn VGND VGND VPWR VPWR _24628_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25524__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ _15361_/A _15367_/B VGND VGND VPWR VPWR _15361_/X sky130_fd_sc_hd__or2_4
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22593__C _22592_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12573_ _12512_/Y _24881_/Q _12575_/A _12572_/Y VGND VGND VPWR VPWR _12573_/X sky130_fd_sc_hd__a2bb2o_4
X_24559_ _24558_/CLK _16506_/X HRESETn VGND VGND VPWR VPWR _24559_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15769__A HWDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17100_ _16969_/Y _17099_/X _17053_/X VGND VGND VPWR VPWR _17100_/Y sky130_fd_sc_hd__a21oi_4
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14312_ _25171_/Q _14294_/A _14296_/X _13480_/A _14295_/A VGND VGND VPWR VPWR _25171_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11795__B2 _11794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15292_ _15292_/A _15361_/A _15292_/C VGND VGND VPWR VPWR _15347_/A sky130_fd_sc_hd__or3_4
X_18080_ _18227_/A _18075_/X _18079_/X VGND VGND VPWR VPWR _18080_/X sky130_fd_sc_hd__or3_4
XFILLER_157_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _14243_/A VGND VGND VPWR VPWR _21155_/B sky130_fd_sc_hd__buf_2
X_17031_ _16984_/Y _17103_/A _17030_/X VGND VGND VPWR VPWR _17031_/X sky130_fd_sc_hd__or3_4
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13289__A _13289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17984__A _18090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14174_ _20503_/A VGND VGND VPWR VPWR _14174_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_61_0_HCLK clkbuf_7_61_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13125_ _13125_/A _13125_/B _13125_/C _20805_/A VGND VGND VPWR VPWR _13125_/X sky130_fd_sc_hd__or4_4
XFILLER_140_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18982_ _18979_/Y _18977_/X _18981_/X _18977_/X VGND VGND VPWR VPWR _23897_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24477__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13056_ _12976_/D _13032_/B _12998_/A _13054_/B VGND VGND VPWR VPWR _13057_/A sky130_fd_sc_hd__a211o_4
X_17933_ _17949_/A _19024_/A VGND VGND VPWR VPWR _17934_/C sky130_fd_sc_hd__or2_4
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12007_ _12007_/A VGND VGND VPWR VPWR _12007_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24406__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21231__B2 _15661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17864_ _16915_/A _17864_/B VGND VGND VPWR VPWR _17866_/B sky130_fd_sc_hd__or2_4
XFILLER_39_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19603_ _19603_/A VGND VGND VPWR VPWR _19603_/X sky130_fd_sc_hd__buf_2
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16815_ _14964_/Y _16813_/X HWDATA[20] _16813_/X VGND VGND VPWR VPWR _16815_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17795_ _16940_/Y _17763_/X _17555_/X VGND VGND VPWR VPWR _17795_/X sky130_fd_sc_hd__or3_4
XFILLER_93_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19534_ _11774_/A VGND VGND VPWR VPWR _19534_/X sky130_fd_sc_hd__buf_2
X_16746_ _15020_/Y _16745_/X _16483_/X _16745_/X VGND VGND VPWR VPWR _24467_/D sky130_fd_sc_hd__a2bb2o_4
X_13958_ _13957_/Y _13958_/B VGND VGND VPWR VPWR _13958_/X sky130_fd_sc_hd__and2_4
XFILLER_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18935__B1 _17415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12909_ _12889_/X _12904_/X _12908_/X VGND VGND VPWR VPWR _25385_/D sky130_fd_sc_hd__and3_4
X_19465_ _19465_/A VGND VGND VPWR VPWR _21947_/B sky130_fd_sc_hd__inv_2
XFILLER_179_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15749__B1 _24866_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16677_ _24495_/Q VGND VGND VPWR VPWR _16677_/Y sky130_fd_sc_hd__inv_2
X_13889_ _13943_/A VGND VGND VPWR VPWR _13934_/B sky130_fd_sc_hd__inv_2
XFILLER_62_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18416_ _24187_/Q VGND VGND VPWR VPWR _18416_/Y sky130_fd_sc_hd__inv_2
X_15628_ _15608_/A VGND VGND VPWR VPWR _15628_/X sky130_fd_sc_hd__buf_2
X_19396_ _19388_/Y VGND VGND VPWR VPWR _19396_/X sky130_fd_sc_hd__buf_2
XFILLER_61_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18347_ _18344_/X VGND VGND VPWR VPWR _18347_/Y sky130_fd_sc_hd__inv_2
X_15559_ _15559_/A VGND VGND VPWR VPWR _15559_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18278_ _19455_/A VGND VGND VPWR VPWR _18280_/A sky130_fd_sc_hd__buf_2
X_17229_ _17228_/X VGND VGND VPWR VPWR _17341_/A sky130_fd_sc_hd__buf_2
XFILLER_238_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13199__A _13199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19112__B1 _19067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20240_ _23450_/Q VGND VGND VPWR VPWR _20240_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20171_ _20158_/Y VGND VGND VPWR VPWR _20171_/X sky130_fd_sc_hd__buf_2
XFILLER_171_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_238_0_HCLK clkbuf_8_239_0_HCLK/A VGND VGND VPWR VPWR _25050_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24147__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23930_ _25100_/CLK _20991_/X HRESETn VGND VGND VPWR VPWR _23930_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23861_ _23806_/CLK _19087_/X VGND VGND VPWR VPWR _19085_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_123_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22812_ _22781_/X _22784_/X _22793_/Y _22811_/X VGND VGND VPWR VPWR HRDATA[16] sky130_fd_sc_hd__a211o_4
XFILLER_226_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23792_ _23464_/CLK _23792_/D VGND VGND VPWR VPWR _19281_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_65_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18926__B1 _16849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22722__A1 _24762_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22722__B2 _21833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22743_ _16582_/A _21098_/X _21738_/X _22742_/X VGND VGND VPWR VPWR _22743_/X sky130_fd_sc_hd__a211o_4
X_25531_ _25524_/CLK _25531_/D HRESETn VGND VGND VPWR VPWR _25531_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25462_ _25382_/CLK _12389_/X HRESETn VGND VGND VPWR VPWR _12204_/A sky130_fd_sc_hd__dfrtp_4
X_22674_ _16587_/Y _22821_/B _21582_/X _22673_/X VGND VGND VPWR VPWR _22674_/X sky130_fd_sc_hd__o22a_4
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24413_ _24413_/CLK _16857_/X HRESETn VGND VGND VPWR VPWR _24413_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_241_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21625_ _22379_/A _19911_/Y VGND VGND VPWR VPWR _21625_/X sky130_fd_sc_hd__or2_4
X_25393_ _24809_/CLK _25393_/D HRESETn VGND VGND VPWR VPWR _12878_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_21_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11910__A _19610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24344_ _24172_/CLK _17376_/X HRESETn VGND VGND VPWR VPWR _17241_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_166_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21556_ _21556_/A VGND VGND VPWR VPWR _21556_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20507_ _25152_/Q _14484_/X _20505_/X _20466_/X _20506_/X VGND VGND VPWR VPWR _20507_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24988__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24275_ _24275_/CLK _24275_/D HRESETn VGND VGND VPWR VPWR _16921_/A sky130_fd_sc_hd__dfrtp_4
X_21487_ _21487_/A _19983_/Y VGND VGND VPWR VPWR _21488_/C sky130_fd_sc_hd__or2_4
XFILLER_148_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12726__B1 _12627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23226_ _22552_/X _23225_/X _23050_/X _17541_/A _22555_/X VGND VGND VPWR VPWR _23226_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24917__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20438_ _13965_/X _20605_/A _20436_/X _20437_/X VGND VGND VPWR VPWR _20438_/X sky130_fd_sc_hd__or4_4
XFILLER_106_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_48_0_HCLK clkbuf_5_24_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_97_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_23157_ _23157_/A _23156_/X VGND VGND VPWR VPWR _23157_/X sky130_fd_sc_hd__or2_4
X_20369_ _20369_/A _21215_/A VGND VGND VPWR VPWR _20369_/X sky130_fd_sc_hd__or2_4
XFILLER_162_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22108_ _14467_/Y _21721_/B _25107_/Q _22119_/B VGND VGND VPWR VPWR _22108_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24570__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23088_ _24604_/Q _23088_/B VGND VGND VPWR VPWR _23091_/B sky130_fd_sc_hd__or2_4
XANTENNA__12460__B _12191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13151__B1 _13150_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14930_ _25017_/Q _24423_/Q _15251_/A _14929_/Y VGND VGND VPWR VPWR _14930_/X sky130_fd_sc_hd__o22a_4
X_22039_ _21954_/A _22018_/Y _22025_/Y _22032_/Y _22038_/Y VGND VGND VPWR VPWR _22039_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19524__A _16721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22961__B2 _21051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14861_ _14860_/X VGND VGND VPWR VPWR _14861_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15979__B1 _21088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16600_ _16600_/A VGND VGND VPWR VPWR _16600_/Y sky130_fd_sc_hd__inv_2
X_13812_ _22695_/A _13810_/X _11735_/X _13810_/X VGND VGND VPWR VPWR _25269_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_180_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_HCLK clkbuf_4_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_17580_ _17530_/Y _17578_/Y _17580_/C _17580_/D VGND VGND VPWR VPWR _17581_/C sky130_fd_sc_hd__or4_4
X_14792_ _25055_/Q VGND VGND VPWR VPWR _14814_/C sky130_fd_sc_hd__inv_2
XFILLER_75_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22885__A _23172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20319__A3 _18257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16531_ _16530_/Y _16528_/X _16353_/X _16528_/X VGND VGND VPWR VPWR _24550_/D sky130_fd_sc_hd__a2bb2o_4
X_13743_ _13732_/X VGND VGND VPWR VPWR _13743_/X sky130_fd_sc_hd__buf_2
XANTENNA__17979__A _18054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19250_ _21240_/B _19245_/X _19091_/X _19232_/Y VGND VGND VPWR VPWR _23803_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16462_ _16458_/Y _16454_/X _16459_/X _16461_/X VGND VGND VPWR VPWR _24576_/D sky130_fd_sc_hd__a2bb2o_4
X_13674_ _11814_/Y _13673_/X VGND VGND VPWR VPWR _13675_/B sky130_fd_sc_hd__or2_4
XFILLER_188_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23269__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18201_ _18095_/A _18199_/X _18201_/C VGND VGND VPWR VPWR _18205_/B sky130_fd_sc_hd__and3_4
XFILLER_232_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15413_ _15411_/Y _15413_/B _15402_/X VGND VGND VPWR VPWR _24979_/D sky130_fd_sc_hd__and3_4
X_12625_ _12648_/A _12625_/B _12624_/X VGND VGND VPWR VPWR _25430_/D sky130_fd_sc_hd__and3_4
X_19181_ _23827_/Q VGND VGND VPWR VPWR _19181_/Y sky130_fd_sc_hd__inv_2
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15499__A _15489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16393_ _16387_/A VGND VGND VPWR VPWR _16393_/X sky130_fd_sc_hd__buf_2
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18132_ _18132_/A _18132_/B _18132_/C VGND VGND VPWR VPWR _18132_/X sky130_fd_sc_hd__and3_4
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12556_ _12555_/Y _24869_/Q _12555_/Y _24869_/Q VGND VGND VPWR VPWR _12556_/X sky130_fd_sc_hd__a2bb2o_4
X_15344_ _15343_/X VGND VGND VPWR VPWR _24998_/D sky130_fd_sc_hd__inv_2
XANTENNA__16156__B1 _15466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18063_ _15691_/X _18043_/X _18062_/X _24248_/Q _18022_/X VGND VGND VPWR VPWR _18063_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12211_/Y _12493_/B VGND VGND VPWR VPWR _12491_/B sky130_fd_sc_hd__or2_4
X_15275_ _14976_/X _15273_/X _15274_/Y VGND VGND VPWR VPWR _15275_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15903__B1 _24785_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17014_ _16995_/X _17000_/X _17008_/X _17014_/D VGND VGND VPWR VPWR _17014_/X sky130_fd_sc_hd__or4_4
X_14226_ _14224_/Y _14225_/X _13791_/X _14225_/X VGND VGND VPWR VPWR _14226_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24658__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12193__A1 _25441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14157_ _14100_/X _14156_/Y _25133_/Q _14100_/X VGND VGND VPWR VPWR _14157_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13108_ _20781_/A _13108_/B _13108_/C _13108_/D VGND VGND VPWR VPWR _13122_/B sky130_fd_sc_hd__or4_4
X_14088_ _14102_/C _14087_/X _14088_/C VGND VGND VPWR VPWR _14088_/X sky130_fd_sc_hd__or3_4
X_18965_ _18965_/A VGND VGND VPWR VPWR _18965_/X sky130_fd_sc_hd__buf_2
XFILLER_113_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15131__B2 _24603_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24240__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13039_ _13038_/X VGND VGND VPWR VPWR _25355_/D sky130_fd_sc_hd__inv_2
X_17916_ _15680_/A _14764_/X _15908_/X _17915_/X VGND VGND VPWR VPWR _17917_/B sky130_fd_sc_hd__a211o_4
XFILLER_239_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18896_ _20994_/A VGND VGND VPWR VPWR _18896_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17847_ _17847_/A VGND VGND VPWR VPWR _17847_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_68_0_HCLK clkbuf_7_34_0_HCLK/X VGND VGND VPWR VPWR _24275_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__13482__A _16181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17778_ _16945_/X _17768_/D VGND VGND VPWR VPWR _17779_/A sky130_fd_sc_hd__or2_4
XFILLER_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18908__B1 HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19517_ _19517_/A VGND VGND VPWR VPWR _21492_/B sky130_fd_sc_hd__inv_2
X_16729_ _16725_/A VGND VGND VPWR VPWR _16730_/A sky130_fd_sc_hd__buf_2
XFILLER_207_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19448_ _19446_/Y _19447_/X _19357_/X _19447_/X VGND VGND VPWR VPWR _19448_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15737__A3 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19379_ _18136_/B VGND VGND VPWR VPWR _19379_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14945__B2 _24428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21410_ _14688_/A _21408_/X _21409_/X VGND VGND VPWR VPWR _21410_/X sky130_fd_sc_hd__and3_4
XFILLER_176_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22390_ _21773_/X _22389_/X _14710_/A VGND VGND VPWR VPWR _22390_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__21712__A2_N _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21140__B1 _14171_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21341_ _24516_/Q _21336_/X _15663_/A _21340_/X VGND VGND VPWR VPWR _21342_/C sky130_fd_sc_hd__a211o_4
XANTENNA__21691__A1 _13783_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24060_ _24060_/CLK _20938_/X HRESETn VGND VGND VPWR VPWR _24060_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24399__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21272_ _21268_/X _21271_/X _14672_/A VGND VGND VPWR VPWR _21272_/X sky130_fd_sc_hd__o21a_4
X_23011_ _23251_/A _23008_/X _23010_/X VGND VGND VPWR VPWR _23011_/X sky130_fd_sc_hd__and3_4
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20223_ _20219_/Y _20222_/X _18250_/X _20222_/X VGND VGND VPWR VPWR _23458_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21443__A1 _21305_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24328__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21443__B2 _22523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16033__A _16038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20154_ _23483_/Q VGND VGND VPWR VPWR _21259_/B sky130_fd_sc_hd__inv_2
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15872__A _15861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20085_ _23506_/Q VGND VGND VPWR VPWR _22375_/B sky130_fd_sc_hd__inv_2
X_24962_ _24959_/CLK _24962_/D HRESETn VGND VGND VPWR VPWR _13916_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_245_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23913_ _23452_/CLK _18937_/X VGND VGND VPWR VPWR _13208_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_217_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24893_ _24035_/CLK _15635_/X HRESETn VGND VGND VPWR VPWR _15634_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11905__A _19606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23844_ _23844_/CLK _19136_/X VGND VGND VPWR VPWR _23844_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__23963__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23775_ _24089_/CLK _23775_/D VGND VGND VPWR VPWR _23775_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17799__A _24283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20987_ _20987_/A _20987_/B _20987_/C VGND VGND VPWR VPWR _23931_/D sky130_fd_sc_hd__and3_4
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20706__B1 _20696_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22171__A2 _21349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25514_ _24679_/CLK _11885_/X HRESETn VGND VGND VPWR VPWR _25514_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22726_ _22726_/A _22726_/B _22717_/X _22725_/Y VGND VGND VPWR VPWR HRDATA[14] sky130_fd_sc_hd__or4_4
XFILLER_159_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22657_ _21087_/A VGND VGND VPWR VPWR _22658_/B sky130_fd_sc_hd__buf_2
X_25445_ _25453_/CLK _25445_/D HRESETn VGND VGND VPWR VPWR _25445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11736__A1_N _11732_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12410_ _12410_/A VGND VGND VPWR VPWR _12410_/Y sky130_fd_sc_hd__inv_2
X_21608_ _21769_/A _21605_/X _21607_/X VGND VGND VPWR VPWR _21608_/X sky130_fd_sc_hd__and3_4
X_13390_ _13390_/A _13390_/B _13390_/C VGND VGND VPWR VPWR _13394_/B sky130_fd_sc_hd__and3_4
XFILLER_185_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_11_0_HCLK clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_22588_ _22521_/B _22585_/X _22423_/X _22587_/X VGND VGND VPWR VPWR _22588_/X sky130_fd_sc_hd__o22a_4
X_25376_ _25369_/CLK _25376_/D HRESETn VGND VGND VPWR VPWR _12755_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_223_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21131__B1 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12341_ _12340_/Y _24833_/Q _12340_/Y _24833_/Q VGND VGND VPWR VPWR _12341_/X sky130_fd_sc_hd__a2bb2o_4
X_21539_ _21087_/A VGND VGND VPWR VPWR _22130_/B sky130_fd_sc_hd__buf_2
X_24327_ _24976_/CLK _24327_/D HRESETn VGND VGND VPWR VPWR _24327_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15060_ _14898_/A VGND VGND VPWR VPWR _15210_/A sky130_fd_sc_hd__inv_2
XFILLER_181_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24751__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12272_ _25454_/Q VGND VGND VPWR VPWR _12272_/Y sky130_fd_sc_hd__inv_2
X_24258_ _24263_/CLK _17889_/X HRESETn VGND VGND VPWR VPWR _21059_/A sky130_fd_sc_hd__dfrtp_4
X_14011_ _14022_/B VGND VGND VPWR VPWR _14011_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23209_ _23209_/A _23206_/X _23208_/X VGND VGND VPWR VPWR _23214_/C sky130_fd_sc_hd__and3_4
XANTENNA__24069__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22631__B1 _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24189_ _24188_/CLK _24189_/D HRESETn VGND VGND VPWR VPWR _24189_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22599__B _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18750_ _24147_/Q _18749_/Y VGND VGND VPWR VPWR _18752_/B sky130_fd_sc_hd__or2_4
XANTENNA__19254__A _19253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15962_ _15955_/X _15958_/X _16236_/A _24760_/Q _15956_/X VGND VGND VPWR VPWR _15962_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_110_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_221_0_HCLK clkbuf_7_110_0_HCLK/X VGND VGND VPWR VPWR _25028_/CLK sky130_fd_sc_hd__clkbuf_1
X_17701_ _17580_/D _17602_/X _17604_/X _17698_/Y VGND VGND VPWR VPWR _17701_/X sky130_fd_sc_hd__a211o_4
XFILLER_248_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14913_ _14913_/A VGND VGND VPWR VPWR _15189_/A sky130_fd_sc_hd__inv_2
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18681_ _18681_/A VGND VGND VPWR VPWR _18682_/D sky130_fd_sc_hd__inv_2
XANTENNA__11686__B1 _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15893_ _12757_/Y _15889_/X _15754_/X _15892_/X VGND VGND VPWR VPWR _24793_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14398__A _14408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17632_ _17502_/A _17631_/Y VGND VGND VPWR VPWR _17632_/X sky130_fd_sc_hd__or2_4
XFILLER_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14844_ _14796_/A _14796_/B _14796_/A _14796_/B VGND VGND VPWR VPWR _14844_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17563_ _17563_/A VGND VGND VPWR VPWR _17563_/Y sky130_fd_sc_hd__inv_2
X_14775_ _14775_/A VGND VGND VPWR VPWR _14775_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11987_ _11985_/X VGND VGND VPWR VPWR _11987_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19302_ _19297_/Y _19300_/X _19301_/X _19300_/X VGND VGND VPWR VPWR _19302_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16514_ _16512_/Y _16508_/X _16141_/X _16513_/X VGND VGND VPWR VPWR _16514_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_232_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13726_ _13726_/A _14758_/A VGND VGND VPWR VPWR _13726_/X sky130_fd_sc_hd__or2_4
XANTENNA__18905__A3 HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17494_ _17494_/A VGND VGND VPWR VPWR _17494_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16377__B1 _15996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16916__A2 _16915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19233_ _19232_/Y VGND VGND VPWR VPWR _19233_/X sky130_fd_sc_hd__buf_2
X_16445_ _16444_/X VGND VGND VPWR VPWR _22629_/A sky130_fd_sc_hd__buf_2
XFILLER_32_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13657_ _23375_/Q _20826_/B VGND VGND VPWR VPWR _13657_/X sky130_fd_sc_hd__and2_4
XFILLER_176_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15022__A _15022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12608_ _12608_/A _12638_/C _12595_/X _12607_/X VGND VGND VPWR VPWR _12608_/X sky130_fd_sc_hd__or4_4
X_19164_ _19163_/X VGND VGND VPWR VPWR _19170_/A sky130_fd_sc_hd__inv_2
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24839__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16376_ _16387_/A VGND VGND VPWR VPWR _16376_/X sky130_fd_sc_hd__buf_2
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13588_ _19026_/D VGND VGND VPWR VPWR _13588_/X sky130_fd_sc_hd__buf_2
XFILLER_129_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18115_ _17968_/X _18113_/X _18114_/X VGND VGND VPWR VPWR _18115_/X sky130_fd_sc_hd__and3_4
XFILLER_145_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15327_ _15338_/A _15327_/B _15326_/X VGND VGND VPWR VPWR _15327_/X sky130_fd_sc_hd__and3_4
X_12539_ _25403_/Q VGND VGND VPWR VPWR _12717_/A sky130_fd_sc_hd__inv_2
X_19095_ _19094_/X VGND VGND VPWR VPWR _19101_/A sky130_fd_sc_hd__inv_2
XFILLER_144_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24492__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18046_ _18222_/A _18046_/B VGND VGND VPWR VPWR _18047_/C sky130_fd_sc_hd__or2_4
X_15258_ _15269_/A _15256_/X _15257_/X VGND VGND VPWR VPWR _15258_/X sky130_fd_sc_hd__and3_4
XFILLER_172_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12166__B2 _22597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24421__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14209_ _14209_/A VGND VGND VPWR VPWR _14209_/X sky130_fd_sc_hd__buf_2
X_15189_ _15189_/A _15188_/X VGND VGND VPWR VPWR _15190_/A sky130_fd_sc_hd__or2_4
XFILLER_98_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_31_0_HCLK clkbuf_6_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19997_ _22020_/B _19991_/X _19970_/X _19996_/X VGND VGND VPWR VPWR _23544_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18948_ _19063_/A VGND VGND VPWR VPWR _18948_/X sky130_fd_sc_hd__buf_2
XFILLER_228_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22925__B2 _21315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18879_ _23945_/Q _20580_/B VGND VGND VPWR VPWR _18880_/B sky130_fd_sc_hd__or2_4
X_20910_ _13650_/X _13637_/D VGND VGND VPWR VPWR _20911_/A sky130_fd_sc_hd__or2_4
X_21890_ _21911_/A _21890_/B _21889_/X VGND VGND VPWR VPWR _21890_/X sky130_fd_sc_hd__and3_4
XFILLER_243_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13418__B2 _11950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16080__A2 _21587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20841_ _20840_/X VGND VGND VPWR VPWR _20841_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18508__A _18823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23560_ _25070_/CLK _19947_/X VGND VGND VPWR VPWR _19945_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20772_ _20771_/X VGND VGND VPWR VPWR _20777_/B sky130_fd_sc_hd__inv_2
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16907__A2 _16906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22511_ _12009_/Y _13456_/X _12080_/Y _12058_/B VGND VGND VPWR VPWR _22511_/X sky130_fd_sc_hd__o22a_4
XFILLER_23_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23491_ _23499_/CLK _20134_/X VGND VGND VPWR VPWR _23491_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22442_ _22442_/A VGND VGND VPWR VPWR _22442_/Y sky130_fd_sc_hd__inv_2
X_25230_ _25230_/CLK _14076_/X HRESETn VGND VGND VPWR VPWR _13991_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_195_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21869__A _21047_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25161_ _25211_/CLK _14347_/X HRESETn VGND VGND VPWR VPWR MSO_S3 sky130_fd_sc_hd__dfrtp_4
XANTENNA__24509__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22373_ _22373_/A _22371_/X _22372_/X VGND VGND VPWR VPWR _22373_/X sky130_fd_sc_hd__and3_4
XFILLER_191_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_113_0_HCLK clkbuf_6_56_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_227_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_24112_ _24315_/CLK _24112_/D HRESETn VGND VGND VPWR VPWR _24112_/Q sky130_fd_sc_hd__dfrtp_4
X_21324_ _15120_/A _22932_/A VGND VGND VPWR VPWR _21333_/B sky130_fd_sc_hd__or2_4
X_25092_ _25089_/CLK _25092_/D HRESETn VGND VGND VPWR VPWR _13566_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12157__A1 _12111_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24043_ _24486_/CLK _24043_/D HRESETn VGND VGND VPWR VPWR _24043_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24162__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21255_ _22199_/A _20111_/Y VGND VGND VPWR VPWR _21256_/C sky130_fd_sc_hd__or2_4
XFILLER_190_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20206_ _20200_/Y VGND VGND VPWR VPWR _20206_/X sky130_fd_sc_hd__buf_2
XANTENNA__18897__B _17438_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21186_ _21204_/A _21184_/X _21185_/X VGND VGND VPWR VPWR _21186_/X sky130_fd_sc_hd__and3_4
X_20137_ _20137_/A VGND VGND VPWR VPWR _20137_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19074__A _19074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25368__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20068_ _20065_/Y _20067_/X _19807_/X _20067_/X VGND VGND VPWR VPWR _20068_/X sky130_fd_sc_hd__a2bb2o_4
X_24945_ _24357_/CLK _15492_/X HRESETn VGND VGND VPWR VPWR _13453_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22392__A2 _22363_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11910_ _19610_/A VGND VGND VPWR VPWR _11910_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12890_ _22667_/A _12920_/A _12588_/X _12835_/X VGND VGND VPWR VPWR _12890_/X sky130_fd_sc_hd__or4_4
X_24876_ _24874_/CLK _24876_/D HRESETn VGND VGND VPWR VPWR _12514_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_51_0_HCLK clkbuf_8_51_0_HCLK/A VGND VGND VPWR VPWR _25292_/CLK sky130_fd_sc_hd__clkbuf_1
X_11841_ _11841_/A VGND VGND VPWR VPWR _11841_/Y sky130_fd_sc_hd__inv_2
X_23827_ _23827_/CLK _23827_/D VGND VGND VPWR VPWR _23827_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11772_/A VGND VGND VPWR VPWR _11772_/Y sky130_fd_sc_hd__inv_2
X_14560_ _14576_/B VGND VGND VPWR VPWR _14561_/B sky130_fd_sc_hd__inv_2
XFILLER_199_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16359__B1 _16358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12093__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23758_ _23767_/CLK _23758_/D VGND VGND VPWR VPWR _19376_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20155__B2 _20137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24951__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _12013_/C _20964_/B _13510_/X VGND VGND VPWR VPWR _25306_/D sky130_fd_sc_hd__a21o_4
XPHY_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22709_ _22709_/A _21235_/A VGND VGND VPWR VPWR _22709_/X sky130_fd_sc_hd__or2_4
XPHY_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _23957_/Q VGND VGND VPWR VPWR _14491_/X sky130_fd_sc_hd__buf_2
XFILLER_198_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23689_ _23706_/CLK _19579_/X VGND VGND VPWR VPWR _19578_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16239_/A VGND VGND VPWR VPWR _16230_/X sky130_fd_sc_hd__buf_2
X_13442_ _13220_/X _13442_/B VGND VGND VPWR VPWR _13442_/X sky130_fd_sc_hd__or2_4
X_25428_ _25428_/CLK _12634_/X HRESETn VGND VGND VPWR VPWR _12503_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_201_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24932__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13373_ _13219_/X _13371_/X _13372_/X VGND VGND VPWR VPWR _13373_/X sky130_fd_sc_hd__and3_4
X_16161_ _21435_/A VGND VGND VPWR VPWR _16161_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15777__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25359_ _25390_/CLK _13023_/X HRESETn VGND VGND VPWR VPWR _12308_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_154_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_5_24_0_HCLK_A clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15112_ _24994_/Q VGND VGND VPWR VPWR _15292_/A sky130_fd_sc_hd__inv_2
X_12324_ _12324_/A VGND VGND VPWR VPWR _12324_/Y sky130_fd_sc_hd__inv_2
X_16092_ _16111_/A VGND VGND VPWR VPWR _16092_/X sky130_fd_sc_hd__buf_2
XFILLER_154_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16531__B1 _16353_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13297__A _13334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12255_ _12254_/Y _23275_/A _12254_/Y _23275_/A VGND VGND VPWR VPWR _12255_/X sky130_fd_sc_hd__a2bb2o_4
X_15043_ _15249_/A _16765_/A _25012_/Q _15022_/Y VGND VGND VPWR VPWR _15049_/A sky130_fd_sc_hd__a2bb2o_4
X_19920_ _19932_/A VGND VGND VPWR VPWR _19920_/X sky130_fd_sc_hd__buf_2
XFILLER_79_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19851_ _19851_/A VGND VGND VPWR VPWR _19851_/Y sky130_fd_sc_hd__inv_2
X_12186_ _12186_/A _12180_/X _12186_/C _12185_/X VGND VGND VPWR VPWR _12186_/X sky130_fd_sc_hd__or4_4
Xclkbuf_5_18_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18802_ _18797_/A _18797_/B _18724_/X _18798_/Y VGND VGND VPWR VPWR _18803_/A sky130_fd_sc_hd__a211o_4
XFILLER_95_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19782_ _23618_/Q VGND VGND VPWR VPWR _19782_/Y sky130_fd_sc_hd__inv_2
X_16994_ _16037_/Y _17029_/A _16037_/Y _17029_/A VGND VGND VPWR VPWR _16995_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23218__B _23217_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18733_ _18733_/A _18733_/B VGND VGND VPWR VPWR _18734_/C sky130_fd_sc_hd__or2_4
XFILLER_110_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15945_ _12181_/Y _15944_/X _15581_/X _15944_/X VGND VGND VPWR VPWR _15945_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21019__A _15697_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25038__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18664_ _16544_/Y _24156_/Q _16544_/Y _24156_/Q VGND VGND VPWR VPWR _18668_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15876_ _12767_/Y _15872_/X _11715_/X _15875_/X VGND VGND VPWR VPWR _15876_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_221_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17615_ _17563_/Y _17615_/B VGND VGND VPWR VPWR _17615_/X sky130_fd_sc_hd__or2_4
X_14827_ _14798_/C _14812_/X _14814_/A _14814_/B VGND VGND VPWR VPWR _14827_/X sky130_fd_sc_hd__o22a_4
XFILLER_224_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18595_ _18595_/A _18595_/B VGND VGND VPWR VPWR _18596_/B sky130_fd_sc_hd__or2_4
XFILLER_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15270__B1 _15185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13760__A _13807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17546_ _25542_/Q _17545_/Y _11710_/Y _17543_/A VGND VGND VPWR VPWR _17546_/X sky130_fd_sc_hd__a2bb2o_4
X_14758_ _14758_/A _14758_/B _14757_/X VGND VGND VPWR VPWR _14758_/X sky130_fd_sc_hd__or3_4
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13709_ _13673_/X _13707_/Y _13708_/X _13701_/X _11810_/A VGND VGND VPWR VPWR _25287_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_189_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17477_ _18900_/A _17472_/X _17476_/X VGND VGND VPWR VPWR _24324_/D sky130_fd_sc_hd__a21oi_4
XFILLER_232_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14689_ _21911_/A VGND VGND VPWR VPWR _21757_/A sky130_fd_sc_hd__buf_2
XFILLER_60_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19216_ _19224_/A VGND VGND VPWR VPWR _19216_/X sky130_fd_sc_hd__buf_2
X_16428_ _15121_/Y _16426_/X _16062_/X _16426_/X VGND VGND VPWR VPWR _24585_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24673__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23096__B1 _11687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16770__B1 _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19147_ _19146_/Y _19143_/X _19122_/X _19143_/X VGND VGND VPWR VPWR _23841_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24602__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16359_ _16357_/Y _16278_/X _16358_/X _16278_/X VGND VGND VPWR VPWR _16359_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22843__B1 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19078_ _23864_/Q VGND VGND VPWR VPWR _22067_/B sky130_fd_sc_hd__inv_2
X_18029_ _18104_/A _23760_/Q VGND VGND VPWR VPWR _18030_/C sky130_fd_sc_hd__or2_4
XFILLER_246_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21040_ _21128_/B VGND VGND VPWR VPWR _21040_/X sky130_fd_sc_hd__buf_2
XFILLER_114_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24070__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22991_ _23060_/A _22991_/B VGND VGND VPWR VPWR _22991_/Y sky130_fd_sc_hd__nor2_4
XFILLER_27_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24730_ _24365_/CLK _16039_/X HRESETn VGND VGND VPWR VPWR _24730_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21942_ _17709_/A _21940_/X _21942_/C VGND VGND VPWR VPWR _21942_/X sky130_fd_sc_hd__and3_4
XANTENNA__20385__A1 _23393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_38_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_77_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21873_ _11664_/B VGND VGND VPWR VPWR _22435_/A sky130_fd_sc_hd__buf_2
X_24661_ _24592_/CLK _24661_/D HRESETn VGND VGND VPWR VPWR _22705_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22126__A2 _22109_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19527__B1 _19414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _20824_/A VGND VGND VPWR VPWR _20846_/A sky130_fd_sc_hd__buf_2
X_23612_ _23627_/CLK _19799_/X VGND VGND VPWR VPWR _13414_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24592_ _24592_/CLK _24592_/D HRESETn VGND VGND VPWR VPWR _16415_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20755_ _20754_/X VGND VGND VPWR VPWR _20755_/Y sky130_fd_sc_hd__inv_2
X_23543_ _23415_/CLK _23543_/D VGND VGND VPWR VPWR _19998_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23474_ _23490_/CLK _23474_/D VGND VGND VPWR VPWR _20177_/A sky130_fd_sc_hd__dfxtp_4
X_20686_ _20686_/A VGND VGND VPWR VPWR _20708_/A sky130_fd_sc_hd__buf_2
XANTENNA__16761__B1 _15741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_HCLK clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22425_ _12762_/A _22299_/X _22424_/X VGND VGND VPWR VPWR _22425_/X sky130_fd_sc_hd__a21o_4
X_25213_ _23951_/CLK _14157_/X HRESETn VGND VGND VPWR VPWR _14087_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__24343__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22356_ _22352_/X _22355_/X _21686_/X VGND VGND VPWR VPWR _22356_/Y sky130_fd_sc_hd__o21ai_4
X_25144_ _25113_/CLK _14404_/X HRESETn VGND VGND VPWR VPWR _14117_/A sky130_fd_sc_hd__dfstp_4
XFILLER_191_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21307_ _21859_/A VGND VGND VPWR VPWR _22712_/A sky130_fd_sc_hd__buf_2
X_25075_ _23890_/CLK _25075_/D HRESETn VGND VGND VPWR VPWR _13590_/A sky130_fd_sc_hd__dfrtp_4
X_22287_ _21597_/A VGND VGND VPWR VPWR _22287_/X sky130_fd_sc_hd__buf_2
XFILLER_136_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ _21574_/B VGND VGND VPWR VPWR _12087_/B sky130_fd_sc_hd__buf_2
X_24026_ _24501_/CLK _20792_/Y HRESETn VGND VGND VPWR VPWR _20789_/A sky130_fd_sc_hd__dfrtp_4
X_21238_ _21262_/A _21238_/B VGND VGND VPWR VPWR _21238_/X sky130_fd_sc_hd__or2_4
XANTENNA__18266__B1 _16778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22223__A _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17317__A _17314_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13845__A _23995_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21169_ _16265_/Y _15662_/A _16180_/A _21168_/X VGND VGND VPWR VPWR _21175_/B sky130_fd_sc_hd__a211o_4
XFILLER_172_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13991_ _13991_/A _13991_/B _25233_/Q _13991_/D VGND VGND VPWR VPWR _14006_/A sky130_fd_sc_hd__or4_4
XFILLER_218_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15730_ _12572_/Y _15728_/X _11711_/X _15728_/X VGND VGND VPWR VPWR _15730_/X sky130_fd_sc_hd__a2bb2o_4
X_12942_ _12772_/A _12941_/Y VGND VGND VPWR VPWR _12944_/B sky130_fd_sc_hd__or2_4
X_24928_ _25325_/CLK _15532_/X HRESETn VGND VGND VPWR VPWR _11667_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_207_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20678__A _20678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15661_ _15661_/A VGND VGND VPWR VPWR _15662_/A sky130_fd_sc_hd__buf_2
XFILLER_206_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12873_ _12873_/A VGND VGND VPWR VPWR _25394_/D sky130_fd_sc_hd__inv_2
X_24859_ _24855_/CLK _24859_/D HRESETn VGND VGND VPWR VPWR _24859_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15252__B1 _15185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18148__A _18052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _17399_/X VGND VGND VPWR VPWR _17401_/A sky130_fd_sc_hd__buf_2
XFILLER_233_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14612_ _14619_/A _14607_/Y _14611_/Y VGND VGND VPWR VPWR _14612_/X sky130_fd_sc_hd__a21o_4
XPHY_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _24231_/Q VGND VGND VPWR VPWR _11824_/Y sky130_fd_sc_hd__inv_2
X_18380_ _18378_/Y _18374_/X _24195_/Q _18379_/X VGND VGND VPWR VPWR _24196_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12066__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15591_/Y _15589_/X _11721_/X _15589_/X VGND VGND VPWR VPWR _24910_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14395__B _14425_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17248_/Y _17304_/X _17276_/X _17327_/Y VGND VGND VPWR VPWR _17331_/X sky130_fd_sc_hd__a211o_4
XFILLER_42_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14543_ _25098_/Q VGND VGND VPWR VPWR _14543_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21876__A1 _24752_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _25528_/Q VGND VGND VPWR VPWR _11755_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21876__B2 _23138_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _17261_/Y _17258_/X VGND VGND VPWR VPWR _17262_/X sky130_fd_sc_hd__or2_4
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14474_ _25116_/Q VGND VGND VPWR VPWR _14474_/Y sky130_fd_sc_hd__inv_2
X_11686_ _11650_/Y _11684_/X _11685_/X _11684_/X VGND VGND VPWR VPWR _11686_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16752__B1 _16400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19001_ _13606_/A _19116_/B _14648_/A VGND VGND VPWR VPWR _19163_/C sky130_fd_sc_hd__or3_4
XFILLER_146_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16213_ _16212_/Y _16210_/X _15946_/X _16210_/X VGND VGND VPWR VPWR _16213_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24084__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13425_ _13393_/A _13425_/B _13425_/C VGND VGND VPWR VPWR _13425_/X sky130_fd_sc_hd__and3_4
XANTENNA__21302__A _22829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17193_ _24350_/Q VGND VGND VPWR VPWR _17193_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23093__A3 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24013__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16144_ _16144_/A VGND VGND VPWR VPWR _16144_/Y sky130_fd_sc_hd__inv_2
X_13356_ _13388_/A _19061_/A VGND VGND VPWR VPWR _13356_/X sky130_fd_sc_hd__or2_4
XANTENNA__16504__B1 _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12307_ _12305_/A _24828_/Q _13073_/A _12306_/Y VGND VGND VPWR VPWR _12314_/B sky130_fd_sc_hd__o22a_4
XFILLER_114_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18608__A2_N _24142_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16075_ _16077_/A _15771_/B VGND VGND VPWR VPWR _16075_/X sky130_fd_sc_hd__or2_4
XFILLER_142_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13287_ _13390_/A _13285_/X _13287_/C VGND VGND VPWR VPWR _13293_/B sky130_fd_sc_hd__and3_4
XFILLER_114_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15026_ _15026_/A VGND VGND VPWR VPWR _15246_/C sky130_fd_sc_hd__inv_2
X_19903_ _19902_/Y _19900_/X _19810_/X _19900_/X VGND VGND VPWR VPWR _19903_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_216_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12238_ _12443_/A _24763_/Q _12443_/A _24763_/Q VGND VGND VPWR VPWR _12238_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12169_ _22276_/A VGND VGND VPWR VPWR _12169_/Y sky130_fd_sc_hd__inv_2
X_19834_ _19833_/X VGND VGND VPWR VPWR _19835_/A sky130_fd_sc_hd__inv_2
X_16977_ _16977_/A _16972_/X _16977_/C _16976_/X VGND VGND VPWR VPWR _16977_/X sky130_fd_sc_hd__or4_4
X_19765_ _19761_/Y _19764_/X _16860_/X _19764_/X VGND VGND VPWR VPWR _23626_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19757__B1 _19711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15491__B1 HADDR[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15928_ _15958_/A VGND VGND VPWR VPWR _15928_/X sky130_fd_sc_hd__buf_2
X_18716_ _18734_/A _18714_/X _18715_/X VGND VGND VPWR VPWR _24155_/D sky130_fd_sc_hd__and3_4
X_19696_ _13233_/B VGND VGND VPWR VPWR _19696_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18647_ _18647_/A _18647_/B _18645_/X _18647_/D VGND VGND VPWR VPWR _18647_/X sky130_fd_sc_hd__or4_4
XFILLER_224_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15859_ _15843_/X _15850_/X _15710_/X _24815_/Q _15857_/X VGND VGND VPWR VPWR _24815_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_224_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24854__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18578_ _18572_/A _18566_/B _18578_/C VGND VGND VPWR VPWR _18578_/X sky130_fd_sc_hd__and3_4
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17529_ _17529_/A VGND VGND VPWR VPWR _17580_/C sky130_fd_sc_hd__inv_2
XFILLER_178_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20540_ _24332_/Q _23965_/Q VGND VGND VPWR VPWR _23961_/D sky130_fd_sc_hd__and2_4
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20471_ _24069_/D VGND VGND VPWR VPWR _20471_/X sky130_fd_sc_hd__buf_2
XFILLER_119_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22210_ _22210_/A _20161_/Y VGND VGND VPWR VPWR _22211_/C sky130_fd_sc_hd__or2_4
X_23190_ _23190_/A _21528_/B VGND VGND VPWR VPWR _23190_/X sky130_fd_sc_hd__or2_4
XFILLER_173_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22141_ _21859_/A VGND VGND VPWR VPWR _22141_/X sky130_fd_sc_hd__buf_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19617__A _19617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18521__A _18823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22072_ _22387_/A _22072_/B VGND VGND VPWR VPWR _22073_/C sky130_fd_sc_hd__or2_4
X_21023_ _12083_/A VGND VGND VPWR VPWR _21151_/A sky130_fd_sc_hd__buf_2
XFILLER_86_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16274__A2 _15986_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19748__B1 _19746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22974_ _21080_/X VGND VGND VPWR VPWR _22974_/X sky130_fd_sc_hd__buf_2
XFILLER_83_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24713_ _24645_/CLK _16080_/X HRESETn VGND VGND VPWR VPWR _24713_/Q sky130_fd_sc_hd__dfrtp_4
X_21925_ _22343_/A _19864_/Y VGND VGND VPWR VPWR _21927_/B sky130_fd_sc_hd__or2_4
XFILLER_216_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12048__B1 _11793_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24595__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24644_ _24903_/CLK _16274_/X HRESETn VGND VGND VPWR VPWR _24644_/Q sky130_fd_sc_hd__dfrtp_4
X_21856_ _21856_/A _21235_/A VGND VGND VPWR VPWR _21859_/B sky130_fd_sc_hd__or2_4
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21858__A1 _24720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24524__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _15563_/Y _20708_/A _20780_/A _20806_/Y VGND VGND VPWR VPWR _20807_/X sky130_fd_sc_hd__o22a_4
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21787_ _21787_/A _21511_/X VGND VGND VPWR VPWR _21787_/X sky130_fd_sc_hd__and2_4
X_24575_ _24574_/CLK _16465_/X HRESETn VGND VGND VPWR VPWR _24575_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_125_0_HCLK clkbuf_7_62_0_HCLK/X VGND VGND VPWR VPWR _25403_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23526_ _23526_/CLK _20044_/X VGND VGND VPWR VPWR _20043_/A sky130_fd_sc_hd__dfxtp_4
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_188_0_HCLK clkbuf_7_94_0_HCLK/X VGND VGND VPWR VPWR _25113_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20738_ _20738_/A VGND VGND VPWR VPWR _20738_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16734__B1 _16467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21122__A _22992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20669_ _14215_/Y _20615_/A _20629_/A _20668_/Y VGND VGND VPWR VPWR _20670_/A sky130_fd_sc_hd__a211o_4
X_23457_ _23456_/CLK _23457_/D VGND VGND VPWR VPWR _20224_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12744__A _25394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ _13422_/A VGND VGND VPWR VPWR _13300_/A sky130_fd_sc_hd__buf_2
XFILLER_167_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22408_ _24265_/Q _21111_/X _21525_/A VGND VGND VPWR VPWR _22408_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22283__A1 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14190_ _14190_/A VGND VGND VPWR VPWR _14190_/X sky130_fd_sc_hd__buf_2
XANTENNA__22283__B2 _22282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23388_ _23388_/CLK _20399_/X VGND VGND VPWR VPWR _13331_/B sky130_fd_sc_hd__dfxtp_4
X_13141_ _13168_/A _13141_/B VGND VGND VPWR VPWR _13141_/X sky130_fd_sc_hd__or2_4
X_25127_ _23927_/CLK _25127_/D HRESETn VGND VGND VPWR VPWR _14447_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_136_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22339_ _22343_/A _22339_/B VGND VGND VPWR VPWR _22341_/B sky130_fd_sc_hd__or2_4
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16583__A1_N _16582_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25383__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13072_ _13072_/A _13072_/B VGND VGND VPWR VPWR _13073_/B sky130_fd_sc_hd__or2_4
X_25058_ _23665_/CLK _14779_/X HRESETn VGND VGND VPWR VPWR _14769_/B sky130_fd_sc_hd__dfrtp_4
X_12023_ _12022_/Y _12020_/X _12024_/A _12020_/X VGND VGND VPWR VPWR _25492_/D sky130_fd_sc_hd__a2bb2o_4
X_16900_ _16163_/Y _21059_/A _16163_/Y _21059_/A VGND VGND VPWR VPWR _16901_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_183_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19987__B1 _19874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24009_ _24900_/CLK _20715_/Y HRESETn VGND VGND VPWR VPWR _13116_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17880_ _17880_/A _17850_/X VGND VGND VPWR VPWR _17880_/X sky130_fd_sc_hd__or2_4
XFILLER_151_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16831_ _16831_/A VGND VGND VPWR VPWR _16831_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25302__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15473__B1 _15472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19550_ _19549_/Y VGND VGND VPWR VPWR _19550_/X sky130_fd_sc_hd__buf_2
X_16762_ _15014_/Y _16760_/X _15743_/X _16760_/X VGND VGND VPWR VPWR _16762_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13974_ _14005_/A _14005_/B VGND VGND VPWR VPWR _13975_/A sky130_fd_sc_hd__or2_4
X_18501_ _18440_/Y _18499_/X _18500_/X _18495_/B VGND VGND VPWR VPWR _18502_/A sky130_fd_sc_hd__a211o_4
X_15713_ _15759_/A VGND VGND VPWR VPWR _15713_/X sky130_fd_sc_hd__buf_2
XFILLER_207_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12925_ _12920_/A _12919_/X _12872_/A _12921_/Y VGND VGND VPWR VPWR _12926_/A sky130_fd_sc_hd__a211o_4
X_19481_ _19480_/X VGND VGND VPWR VPWR _19494_/A sky130_fd_sc_hd__inv_2
XFILLER_74_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17214__B2 _17347_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16693_ _16691_/Y _16692_/X _16420_/X _16692_/X VGND VGND VPWR VPWR _16693_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12919__A _12617_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18432_ _16228_/Y _18465_/A _16228_/Y _18465_/A VGND VGND VPWR VPWR _18432_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15644_ _15644_/A VGND VGND VPWR VPWR _16268_/A sky130_fd_sc_hd__buf_2
XFILLER_234_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_21_0_HCLK clkbuf_7_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12856_ _12855_/X VGND VGND VPWR VPWR _25398_/D sky130_fd_sc_hd__inv_2
XANTENNA__23299__B1 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12638__B _12606_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24265__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_84_0_HCLK clkbuf_7_85_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_84_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11806_/Y _22620_/A _11806_/Y _22620_/A VGND VGND VPWR VPWR _11813_/B sky130_fd_sc_hd__a2bb2o_4
X_18363_ _18363_/A VGND VGND VPWR VPWR _18363_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15550_/Y VGND VGND VPWR VPWR _15576_/A sky130_fd_sc_hd__buf_2
X_12787_ _12786_/Y VGND VGND VPWR VPWR _12920_/A sky130_fd_sc_hd__buf_2
XFILLER_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13609__A1_N _18060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _17179_/Y _17200_/Y _17314_/C _17305_/X VGND VGND VPWR VPWR _17314_/X sky130_fd_sc_hd__or4_4
XANTENNA__21313__A3 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14526_ _13973_/X _14525_/Y _13984_/X VGND VGND VPWR VPWR _14527_/C sky130_fd_sc_hd__o21a_4
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ HWDATA[13] VGND VGND VPWR VPWR _16233_/A sky130_fd_sc_hd__buf_2
X_18294_ _21208_/A VGND VGND VPWR VPWR _22261_/A sky130_fd_sc_hd__buf_2
XFILLER_186_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22128__A _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ _17336_/A VGND VGND VPWR VPWR _17245_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21032__A _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14457_ _25123_/Q VGND VGND VPWR VPWR _14457_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11669_ _21133_/A _21133_/B VGND VGND VPWR VPWR _13765_/A sky130_fd_sc_hd__or2_4
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _13268_/X _13406_/X _13407_/X VGND VGND VPWR VPWR _13408_/X sky130_fd_sc_hd__and3_4
X_17176_ _24633_/Q _17249_/C _23190_/A _17175_/Y VGND VGND VPWR VPWR _17176_/X sky130_fd_sc_hd__a2bb2o_4
X_14388_ _14388_/A VGND VGND VPWR VPWR _14388_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12373__B _12264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16127_ _16126_/Y _16124_/X _11730_/X _16124_/X VGND VGND VPWR VPWR _16127_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_183_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15965__A _15965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17173__A2_N _17347_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13339_ _13264_/X _13339_/B VGND VGND VPWR VPWR _13339_/X sky130_fd_sc_hd__or2_4
XFILLER_127_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16058_ _16038_/A VGND VGND VPWR VPWR _16058_/X sky130_fd_sc_hd__buf_2
XANTENNA__23223__B1 _24744_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25053__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15009_ _25017_/Q _15008_/A _15251_/A _15008_/Y VGND VGND VPWR VPWR _15009_/X sky130_fd_sc_hd__o22a_4
XFILLER_130_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22798__A _22798_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19817_ _16867_/X VGND VGND VPWR VPWR _19817_/X sky130_fd_sc_hd__buf_2
XANTENNA__16796__A _16796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15464__B1 _14407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19748_ _19745_/Y _19740_/X _19746_/X _19747_/X VGND VGND VPWR VPWR _23632_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19679_ _19677_/Y _19673_/X _19633_/X _19678_/X VGND VGND VPWR VPWR _23656_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21710_ _21532_/X _21706_/Y _22712_/A _21709_/X VGND VGND VPWR VPWR _21710_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19900__A _19900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22690_ _23129_/A VGND VGND VPWR VPWR _23062_/A sky130_fd_sc_hd__buf_2
XANTENNA__15767__B2 _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21641_ _21621_/X _21640_/X _21501_/X VGND VGND VPWR VPWR _21641_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_197_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21572_ _13498_/Y _21570_/X _12026_/Y _21571_/X VGND VGND VPWR VPWR _21572_/X sky130_fd_sc_hd__o22a_4
X_24360_ _24629_/CLK _17316_/X HRESETn VGND VGND VPWR VPWR _24360_/Q sky130_fd_sc_hd__dfrtp_4
X_20523_ _20523_/A _20523_/B _20521_/X _20522_/X VGND VGND VPWR VPWR _20523_/X sky130_fd_sc_hd__or4_4
X_23311_ _21868_/X _23310_/X _22477_/X _24886_/Q _21871_/X VGND VGND VPWR VPWR _23312_/B
+ sky130_fd_sc_hd__a32o_4
X_24291_ _24305_/CLK _24291_/D HRESETn VGND VGND VPWR VPWR _24291_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23988__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20454_ _20445_/A _20449_/X VGND VGND VPWR VPWR _20454_/X sky130_fd_sc_hd__and2_4
X_23242_ _23242_/A _23301_/B VGND VGND VPWR VPWR _23245_/B sky130_fd_sc_hd__or2_4
X_23173_ _16469_/A _23172_/X _23133_/X VGND VGND VPWR VPWR _23173_/X sky130_fd_sc_hd__o21a_4
XFILLER_133_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15875__A _15861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20385_ _23393_/Q _20384_/Y _20986_/A _20384_/A VGND VGND VPWR VPWR _23393_/D sky130_fd_sc_hd__o22a_4
XFILLER_134_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22124_ _20517_/A _21849_/X _23962_/Q _21364_/B VGND VGND VPWR VPWR _22124_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13395__A _13285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22055_ _25260_/Q _22051_/X _13771_/A _22054_/Y VGND VGND VPWR VPWR _22055_/X sky130_fd_sc_hd__a211o_4
XFILLER_121_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21006_ _21006_/A _21006_/B _21006_/C VGND VGND VPWR VPWR _21007_/A sky130_fd_sc_hd__or3_4
XFILLER_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24776__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24705__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22957_ _22824_/X _22948_/Y _22952_/Y _22956_/X VGND VGND VPWR VPWR _22957_/X sky130_fd_sc_hd__a211o_4
XFILLER_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12710_ _12693_/X _12708_/Y _12722_/C VGND VGND VPWR VPWR _25407_/D sky130_fd_sc_hd__and3_4
X_21908_ _21904_/X _21907_/X _22205_/A VGND VGND VPWR VPWR _21908_/X sky130_fd_sc_hd__o21a_4
X_13690_ _13664_/Y VGND VGND VPWR VPWR _13690_/X sky130_fd_sc_hd__buf_2
X_22888_ _16444_/X _22883_/X _22887_/X VGND VGND VPWR VPWR _22895_/C sky130_fd_sc_hd__and3_4
XFILLER_31_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12641_ _12650_/A VGND VGND VPWR VPWR _12641_/X sky130_fd_sc_hd__buf_2
X_24627_ _24623_/CLK _24627_/D HRESETn VGND VGND VPWR VPWR _24627_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21839_ _21836_/X _21839_/B _21838_/X VGND VGND VPWR VPWR _21839_/X sky130_fd_sc_hd__and3_4
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ _15366_/A _15370_/B VGND VGND VPWR VPWR _15367_/B sky130_fd_sc_hd__or2_4
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _24875_/Q VGND VGND VPWR VPWR _12572_/Y sky130_fd_sc_hd__inv_2
X_24558_ _24558_/CLK _24558_/D HRESETn VGND VGND VPWR VPWR _16507_/A sky130_fd_sc_hd__dfrtp_4
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16707__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ _14295_/A _14310_/X _25318_/Q _14294_/A VGND VGND VPWR VPWR _14311_/X sky130_fd_sc_hd__o22a_4
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23509_ _23525_/CLK _23509_/D VGND VGND VPWR VPWR _23509_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15291_ _15291_/A _15366_/A _15356_/A _15125_/Y VGND VGND VPWR VPWR _15292_/C sky130_fd_sc_hd__or4_4
XFILLER_184_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24489_ _24487_/CLK _16693_/X HRESETn VGND VGND VPWR VPWR _24489_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17030_ _16969_/Y _17099_/C _17030_/C _17030_/D VGND VGND VPWR VPWR _17030_/X sky130_fd_sc_hd__or4_4
XFILLER_156_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14242_ _25192_/Q VGND VGND VPWR VPWR _14242_/Y sky130_fd_sc_hd__inv_2
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15785__A _11681_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14173_ _14172_/X VGND VGND VPWR VPWR _25210_/D sky130_fd_sc_hd__inv_2
X_13124_ _20796_/A _20793_/A _13124_/C _20793_/B VGND VGND VPWR VPWR _20805_/A sky130_fd_sc_hd__or4_4
XFILLER_124_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18981_ _18981_/A VGND VGND VPWR VPWR _18981_/X sky130_fd_sc_hd__buf_2
XFILLER_180_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13055_ _13048_/A _13051_/B _13055_/C VGND VGND VPWR VPWR _13055_/X sky130_fd_sc_hd__and3_4
X_17932_ _18016_/A _17932_/B VGND VGND VPWR VPWR _17932_/X sky130_fd_sc_hd__or2_4
X_12006_ _24098_/Q VGND VGND VPWR VPWR _12006_/Y sky130_fd_sc_hd__inv_2
X_17863_ _17862_/X VGND VGND VPWR VPWR _17864_/B sky130_fd_sc_hd__inv_2
X_19602_ _23681_/Q VGND VGND VPWR VPWR _22240_/B sky130_fd_sc_hd__inv_2
X_16814_ _14899_/Y _16813_/X _16483_/X _16813_/X VGND VGND VPWR VPWR _24435_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17794_ _17794_/A VGND VGND VPWR VPWR _17794_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22130__B _22130_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16745_ _16730_/A VGND VGND VPWR VPWR _16745_/X sky130_fd_sc_hd__buf_2
X_19533_ _23703_/Q VGND VGND VPWR VPWR _21960_/A sky130_fd_sc_hd__inv_2
XANTENNA__21027__A _21027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24446__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13957_ _13957_/A VGND VGND VPWR VPWR _13957_/Y sky130_fd_sc_hd__inv_2
X_12908_ _25385_/Q _12907_/Y VGND VGND VPWR VPWR _12908_/X sky130_fd_sc_hd__or2_4
X_19464_ _22026_/B _19458_/X _11911_/X _19463_/X VGND VGND VPWR VPWR _19464_/X sky130_fd_sc_hd__a2bb2o_4
X_16676_ _16675_/Y _16673_/X _16402_/X _16673_/X VGND VGND VPWR VPWR _16676_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13888_ _13888_/A VGND VGND VPWR VPWR _13943_/A sky130_fd_sc_hd__buf_2
XANTENNA__16946__B1 _16154_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15627_ _24896_/Q VGND VGND VPWR VPWR _21746_/A sky130_fd_sc_hd__inv_2
X_18415_ _18408_/X _18415_/B _18412_/X _18415_/D VGND VGND VPWR VPWR _18415_/X sky130_fd_sc_hd__or4_4
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12839_ _12793_/Y _12786_/Y _12837_/X _12839_/D VGND VGND VPWR VPWR _12839_/X sky130_fd_sc_hd__or4_4
X_19395_ _18985_/A VGND VGND VPWR VPWR _19395_/X sky130_fd_sc_hd__buf_2
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18346_ _13157_/X _18341_/A VGND VGND VPWR VPWR _18346_/X sky130_fd_sc_hd__and2_4
XFILLER_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15558_ _15556_/Y _15553_/X _15557_/X _15553_/X VGND VGND VPWR VPWR _15558_/X sky130_fd_sc_hd__a2bb2o_4
X_14509_ _14491_/X _14508_/X _25120_/Q _14506_/X VGND VGND VPWR VPWR _25108_/D sky130_fd_sc_hd__o22a_4
X_18277_ _18276_/X VGND VGND VPWR VPWR _19597_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_171_0_HCLK clkbuf_7_85_0_HCLK/X VGND VGND VPWR VPWR _24089_/CLK sky130_fd_sc_hd__clkbuf_1
X_15489_ _15489_/A VGND VGND VPWR VPWR _15489_/X sky130_fd_sc_hd__buf_2
XANTENNA__17371__B1 _17284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17228_ _17228_/A _17228_/B VGND VGND VPWR VPWR _17228_/X sky130_fd_sc_hd__or2_4
XANTENNA__21697__A _21548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_28_0_HCLK clkbuf_8_29_0_HCLK/A VGND VGND VPWR VPWR _23411_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_190_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17159_ _16990_/A _17159_/B VGND VGND VPWR VPWR _17159_/X sky130_fd_sc_hd__or2_4
XFILLER_190_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20170_ _23477_/Q VGND VGND VPWR VPWR _21630_/B sky130_fd_sc_hd__inv_2
XANTENNA__12112__A1_N _12111_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14488__A1 _23393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11728__A _25535_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12742__A1_N _12741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17415__A _14400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23860_ _23859_/CLK _23860_/D VGND VGND VPWR VPWR _19088_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_85_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22811_ _22796_/Y _23072_/A _22811_/C _22811_/D VGND VGND VPWR VPWR _22811_/X sky130_fd_sc_hd__or4_4
XFILLER_84_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24187__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23791_ _23464_/CLK _23791_/D VGND VGND VPWR VPWR _19285_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_226_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25530_ _24626_/CLK _25530_/D HRESETn VGND VGND VPWR VPWR _25530_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19630__A _18981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24116__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22742_ _24562_/Q _22534_/X _22536_/X VGND VGND VPWR VPWR _22742_/X sky130_fd_sc_hd__o21a_4
XFILLER_225_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23152__A _21232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25461_ _25453_/CLK _25461_/D HRESETn VGND VGND VPWR VPWR _12264_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_241_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22673_ _16503_/Y _22816_/A VGND VGND VPWR VPWR _22673_/X sky130_fd_sc_hd__and2_4
X_24412_ _24413_/CLK _16861_/X HRESETn VGND VGND VPWR VPWR _24412_/Q sky130_fd_sc_hd__dfrtp_4
X_21624_ _22199_/A VGND VGND VPWR VPWR _22379_/A sky130_fd_sc_hd__buf_2
X_25392_ _24809_/CLK _25392_/D HRESETn VGND VGND VPWR VPWR _25392_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24343_ _24346_/CLK _24343_/D HRESETn VGND VGND VPWR VPWR _24343_/Q sky130_fd_sc_hd__dfrtp_4
X_21555_ _21720_/A _21555_/B VGND VGND VPWR VPWR _21601_/A sky130_fd_sc_hd__nor2_4
X_20506_ _20462_/A _14053_/A _20467_/A _20506_/D VGND VGND VPWR VPWR _20506_/X sky130_fd_sc_hd__and4_4
XFILLER_166_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21486_ _22262_/A VGND VGND VPWR VPWR _21487_/A sky130_fd_sc_hd__buf_2
X_24274_ _25450_/CLK _24274_/D HRESETn VGND VGND VPWR VPWR _24274_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20437_ _20437_/A _20445_/A _20437_/C VGND VGND VPWR VPWR _20437_/X sky130_fd_sc_hd__or3_4
X_23225_ _23225_/A _23156_/X VGND VGND VPWR VPWR _23225_/X sky130_fd_sc_hd__or2_4
XANTENNA__21400__A _22213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20368_ _19523_/Y VGND VGND VPWR VPWR _20368_/X sky130_fd_sc_hd__buf_2
X_23156_ _22145_/B VGND VGND VPWR VPWR _23156_/X sky130_fd_sc_hd__buf_2
XANTENNA__18862__B1 _16527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22107_ _22107_/A VGND VGND VPWR VPWR _22109_/C sky130_fd_sc_hd__inv_2
X_23087_ _23087_/A VGND VGND VPWR VPWR _23087_/Y sky130_fd_sc_hd__inv_2
X_20299_ _20299_/A VGND VGND VPWR VPWR _21672_/B sky130_fd_sc_hd__inv_2
X_22038_ _21489_/X _22037_/X _17730_/X VGND VGND VPWR VPWR _22038_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__19524__B _16721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22961__A2 _22559_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14860_ _14817_/X _14808_/B _25044_/Q _14859_/X VGND VGND VPWR VPWR _14860_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15979__A1 _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15979__B2 _15925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13811_ _22734_/A _13810_/X _11730_/X _13810_/X VGND VGND VPWR VPWR _25270_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_217_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14791_ scl_oen_o_S5 _21006_/B _20261_/B VGND VGND VPWR VPWR _14802_/B sky130_fd_sc_hd__and3_4
X_23989_ _25052_/CLK scl_i_S5 HRESETn VGND VGND VPWR VPWR _23989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16530_ _16530_/A VGND VGND VPWR VPWR _16530_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13742_ _19072_/C _13734_/X _20066_/A VGND VGND VPWR VPWR _13742_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__19540__A _11785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16928__B1 _16128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23062__A _23062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16461_ _16470_/A VGND VGND VPWR VPWR _16461_/X sky130_fd_sc_hd__buf_2
XFILLER_71_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13673_ _11810_/Y _13673_/B VGND VGND VPWR VPWR _13673_/X sky130_fd_sc_hd__or2_4
XFILLER_231_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18200_ _18017_/A _18200_/B VGND VGND VPWR VPWR _18201_/C sky130_fd_sc_hd__or2_4
XANTENNA__23269__A3 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15412_ _15296_/A _15410_/X VGND VGND VPWR VPWR _15413_/B sky130_fd_sc_hd__or2_4
XFILLER_188_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25133__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12624_ _12624_/A _12624_/B VGND VGND VPWR VPWR _12624_/X sky130_fd_sc_hd__or2_4
X_19180_ _19179_/Y _19177_/X _19067_/X _19177_/X VGND VGND VPWR VPWR _23828_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16392_ _15144_/Y _16387_/X _16391_/X _16387_/X VGND VGND VPWR VPWR _24602_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12414__B1 _12240_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25196__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18131_ _18099_/A _18131_/B _18131_/C VGND VGND VPWR VPWR _18132_/C sky130_fd_sc_hd__or3_4
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15343_ _15282_/B _15340_/B _15342_/X VGND VGND VPWR VPWR _15343_/X sky130_fd_sc_hd__or3_4
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12555_ _25415_/Q VGND VGND VPWR VPWR _12555_/Y sky130_fd_sc_hd__inv_2
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17353__B1 _17284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_244_0_HCLK clkbuf_7_122_0_HCLK/X VGND VGND VPWR VPWR _24477_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18062_ _18062_/A _18062_/B _18062_/C VGND VGND VPWR VPWR _18062_/X sky130_fd_sc_hd__and3_4
XFILLER_184_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15274_ _14976_/X _15273_/X _15169_/X VGND VGND VPWR VPWR _15274_/Y sky130_fd_sc_hd__a21oi_4
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ _12492_/A _12456_/X VGND VGND VPWR VPWR _12493_/B sky130_fd_sc_hd__or2_4
XANTENNA__22406__A _22821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17013_ _17009_/X _17010_/X _17011_/X _17013_/D VGND VGND VPWR VPWR _17014_/D sky130_fd_sc_hd__or4_4
X_14225_ _14213_/A VGND VGND VPWR VPWR _14225_/X sky130_fd_sc_hd__buf_2
XANTENNA__16404__A _16404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14156_ _14155_/X VGND VGND VPWR VPWR _14156_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14216__A1_N _14215_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13107_ _13107_/A _20767_/A _13107_/C _24022_/Q VGND VGND VPWR VPWR _13108_/D sky130_fd_sc_hd__or4_4
XANTENNA__24698__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14087_ _14154_/A _14162_/A _14160_/A _14087_/D VGND VGND VPWR VPWR _14087_/X sky130_fd_sc_hd__or4_4
X_18964_ _18114_/B VGND VGND VPWR VPWR _18964_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12556__A2_N _24869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13038_ _12357_/Y _13032_/X _12998_/A _13035_/B VGND VGND VPWR VPWR _13038_/X sky130_fd_sc_hd__a211o_4
X_17915_ _15904_/B _14764_/X _14608_/Y VGND VGND VPWR VPWR _17915_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24627__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18895_ _24001_/Q _14524_/Y _20992_/A _14523_/A VGND VGND VPWR VPWR _24118_/D sky130_fd_sc_hd__o22a_4
XFILLER_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17846_ _17756_/Y _17841_/B _17793_/A _17843_/B VGND VGND VPWR VPWR _17847_/A sky130_fd_sc_hd__a211o_4
XFILLER_239_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24280__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14989_ _14989_/A VGND VGND VPWR VPWR _15168_/B sky130_fd_sc_hd__buf_2
X_17777_ _17776_/X VGND VGND VPWR VPWR _24288_/D sky130_fd_sc_hd__inv_2
XANTENNA__24335__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19516_ _21681_/B _19515_/X _11924_/X _19515_/X VGND VGND VPWR VPWR _23709_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16728_ _15012_/Y _16726_/X _16373_/X _16726_/X VGND VGND VPWR VPWR _24476_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16659_ _24502_/Q VGND VGND VPWR VPWR _16659_/Y sky130_fd_sc_hd__inv_2
X_19447_ _19447_/A VGND VGND VPWR VPWR _19447_/X sky130_fd_sc_hd__buf_2
XFILLER_50_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25486__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_54_0_HCLK clkbuf_6_54_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_54_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19378_ _19376_/Y _19372_/X _19377_/X _19372_/X VGND VGND VPWR VPWR _23758_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18329_ _17452_/A VGND VGND VPWR VPWR _19273_/A sky130_fd_sc_hd__buf_2
XANTENNA__21140__B2 _21365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21340_ _16534_/A _21337_/X _21339_/X VGND VGND VPWR VPWR _21340_/X sky130_fd_sc_hd__o21a_4
XFILLER_147_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21271_ _22223_/A _21269_/X _21270_/X VGND VGND VPWR VPWR _21271_/X sky130_fd_sc_hd__and3_4
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19097__B1 _19006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20222_ _20227_/A VGND VGND VPWR VPWR _20222_/X sky130_fd_sc_hd__buf_2
X_23010_ _16564_/A _22730_/X _15663_/X _23009_/X VGND VGND VPWR VPWR _23010_/X sky130_fd_sc_hd__a211o_4
XANTENNA__18844__B1 _16503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20153_ _21401_/B _20150_/X _20109_/X _20150_/X VGND VGND VPWR VPWR _23484_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24368__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20084_ _20083_/Y _20079_/X _19852_/X _20067_/A VGND VGND VPWR VPWR _20084_/X sky130_fd_sc_hd__a2bb2o_4
X_24961_ _24959_/CLK _15453_/X HRESETn VGND VGND VPWR VPWR _13903_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23912_ _23912_/CLK _23912_/D VGND VGND VPWR VPWR _18938_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_100_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24892_ _24907_/CLK _24892_/D HRESETn VGND VGND VPWR VPWR _21018_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_246_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23843_ _23844_/CLK _19139_/X VGND VGND VPWR VPWR _23843_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19360__A _19360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19021__B1 _18951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23774_ _23774_/CLK _19332_/X VGND VGND VPWR VPWR _18121_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _20986_/A VGND VGND VPWR VPWR _20987_/A sky130_fd_sc_hd__inv_2
XPHY_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25513_ _24679_/CLK _11887_/X HRESETn VGND VGND VPWR VPWR _11849_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_225_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22725_ _22725_/A _22724_/X VGND VGND VPWR VPWR _22725_/Y sky130_fd_sc_hd__nor2_4
XFILLER_26_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25444_ _25444_/CLK _25444_/D HRESETn VGND VGND VPWR VPWR _25444_/Q sky130_fd_sc_hd__dfrtp_4
X_22656_ _21077_/X _22656_/B VGND VGND VPWR VPWR _22665_/C sky130_fd_sc_hd__and2_4
XANTENNA__23932__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21607_ _21756_/A _21607_/B VGND VGND VPWR VPWR _21607_/X sky130_fd_sc_hd__or2_4
X_25375_ _25375_/CLK _12950_/X HRESETn VGND VGND VPWR VPWR _12762_/A sky130_fd_sc_hd__dfrtp_4
X_22587_ _17237_/Y _22543_/X _22586_/X VGND VGND VPWR VPWR _22587_/X sky130_fd_sc_hd__o21a_4
XFILLER_138_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12340_ _12340_/A VGND VGND VPWR VPWR _12340_/Y sky130_fd_sc_hd__inv_2
X_24326_ _24326_/CLK _17434_/X HRESETn VGND VGND VPWR VPWR _17433_/A sky130_fd_sc_hd__dfrtp_4
X_21538_ _21537_/X VGND VGND VPWR VPWR _22279_/A sky130_fd_sc_hd__buf_2
XFILLER_154_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15897__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21130__A _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12271_ _12197_/Y _12257_/Y _12271_/C _12270_/X VGND VGND VPWR VPWR _12271_/X sky130_fd_sc_hd__or4_4
X_24257_ _24257_/CLK _24257_/D HRESETn VGND VGND VPWR VPWR _17890_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_11_0_HCLK clkbuf_7_5_0_HCLK/X VGND VGND VPWR VPWR _23487_/CLK sky130_fd_sc_hd__clkbuf_1
X_21469_ _21460_/X _21468_/X _17725_/X VGND VGND VPWR VPWR _21469_/X sky130_fd_sc_hd__o21a_4
XANTENNA__12752__A _25386_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14010_ _13975_/A _14005_/Y _14006_/Y _13975_/Y _14009_/Y VGND VGND VPWR VPWR _14010_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23208_ _24542_/Q _23171_/X _22839_/X _23207_/X VGND VGND VPWR VPWR _23208_/X sky130_fd_sc_hd__a211o_4
XFILLER_181_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_74_0_HCLK clkbuf_8_74_0_HCLK/A VGND VGND VPWR VPWR _25538_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_135_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24188_ _24188_/CLK _18491_/Y HRESETn VGND VGND VPWR VPWR _24188_/Q sky130_fd_sc_hd__dfrtp_4
X_23139_ _16737_/A _23002_/X _22891_/X VGND VGND VPWR VPWR _23139_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24791__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15961_ _15955_/X _15958_/X _16233_/A _24761_/Q _15956_/X VGND VGND VPWR VPWR _15961_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_122_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23057__A _16659_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24720__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14912_ _25016_/Q _24422_/Q _15002_/A _14911_/Y VGND VGND VPWR VPWR _14919_/B sky130_fd_sc_hd__o22a_4
X_17700_ _17696_/B _17700_/B _17688_/C VGND VGND VPWR VPWR _24292_/D sky130_fd_sc_hd__and3_4
XFILLER_191_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24038__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15892_ _15889_/A VGND VGND VPWR VPWR _15892_/X sky130_fd_sc_hd__buf_2
X_18680_ _24130_/Q VGND VGND VPWR VPWR _18787_/A sky130_fd_sc_hd__inv_2
XFILLER_248_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16074__B1 _15475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14843_ _14840_/X _14842_/Y _25195_/Q _14840_/X VGND VGND VPWR VPWR _25050_/D sky130_fd_sc_hd__a2bb2o_4
X_17631_ _17630_/X VGND VGND VPWR VPWR _17631_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14624__B2 _14610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15821__B1 _13818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17562_ _17561_/Y _17494_/Y VGND VGND VPWR VPWR _17597_/A sky130_fd_sc_hd__or2_4
XANTENNA__19012__B1 _18985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14774_ _25059_/Q _14771_/X _14768_/A _14773_/Y VGND VGND VPWR VPWR _25059_/D sky130_fd_sc_hd__o22a_4
X_11986_ _25311_/Q VGND VGND VPWR VPWR _11986_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22698__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16513_ _16521_/A VGND VGND VPWR VPWR _16513_/X sky130_fd_sc_hd__buf_2
X_19301_ _19006_/A VGND VGND VPWR VPWR _19301_/X sky130_fd_sc_hd__buf_2
X_13725_ _13725_/A VGND VGND VPWR VPWR _14758_/A sky130_fd_sc_hd__inv_2
XFILLER_204_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17493_ _24297_/Q VGND VGND VPWR VPWR _17574_/D sky130_fd_sc_hd__inv_2
XFILLER_204_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12927__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16444_ _21845_/A VGND VGND VPWR VPWR _16444_/X sky130_fd_sc_hd__buf_2
X_19232_ _19232_/A VGND VGND VPWR VPWR _19232_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13656_ _20823_/B VGND VGND VPWR VPWR _20826_/B sky130_fd_sc_hd__inv_2
XFILLER_32_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12607_ _12599_/X _12606_/X VGND VGND VPWR VPWR _12607_/X sky130_fd_sc_hd__or2_4
X_19163_ _19320_/A _19163_/B _19163_/C VGND VGND VPWR VPWR _19163_/X sky130_fd_sc_hd__or3_4
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _16375_/A VGND VGND VPWR VPWR _16387_/A sky130_fd_sc_hd__buf_2
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13587_ _14648_/A VGND VGND VPWR VPWR _19026_/D sky130_fd_sc_hd__inv_2
XFILLER_9_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ _18146_/A _18114_/B VGND VGND VPWR VPWR _18114_/X sky130_fd_sc_hd__or2_4
XFILLER_219_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15326_ _15326_/A _15324_/A VGND VGND VPWR VPWR _15326_/X sky130_fd_sc_hd__or2_4
X_12538_ _25410_/Q _24864_/Q _12696_/A _12537_/Y VGND VGND VPWR VPWR _12545_/B sky130_fd_sc_hd__o22a_4
X_19094_ _19209_/A _19094_/B _19094_/C VGND VGND VPWR VPWR _19094_/X sky130_fd_sc_hd__or3_4
XFILLER_129_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22136__A _24898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15888__B1 _24796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18045_ _18118_/A _18045_/B VGND VGND VPWR VPWR _18045_/X sky130_fd_sc_hd__or2_4
XFILLER_145_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15257_ _15251_/A _15254_/X VGND VGND VPWR VPWR _15257_/X sky130_fd_sc_hd__or2_4
XANTENNA__24879__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12469_ _12468_/X VGND VGND VPWR VPWR _12469_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14208_ _14208_/A VGND VGND VPWR VPWR _14209_/A sky130_fd_sc_hd__buf_2
XANTENNA__24808__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15188_ _15065_/A _15187_/X VGND VGND VPWR VPWR _15188_/X sky130_fd_sc_hd__or2_4
XFILLER_126_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22622__B2 _21317_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14139_ _14090_/A _14089_/X _14090_/A _14089_/X VGND VGND VPWR VPWR _14139_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19996_ _19990_/Y VGND VGND VPWR VPWR _19996_/X sky130_fd_sc_hd__buf_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24461__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18947_ _18947_/A VGND VGND VPWR VPWR _18947_/X sky130_fd_sc_hd__buf_2
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22925__A2 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18878_ _23944_/Q _18877_/X VGND VGND VPWR VPWR _20580_/B sky130_fd_sc_hd__or2_4
XFILLER_228_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17829_ _16921_/A _17829_/B VGND VGND VPWR VPWR _17830_/C sky130_fd_sc_hd__or2_4
XFILLER_243_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15812__B1 _24836_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20840_ _16708_/Y _20825_/X _20834_/X _20839_/X VGND VGND VPWR VPWR _20840_/X sky130_fd_sc_hd__o22a_4
XFILLER_81_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22689__B2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20771_ _20754_/A _13108_/D VGND VGND VPWR VPWR _20771_/X sky130_fd_sc_hd__or2_4
XFILLER_23_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22510_ _16272_/X _22509_/X VGND VGND VPWR VPWR _22528_/A sky130_fd_sc_hd__nor2_4
XANTENNA__11741__A _25532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23490_ _23490_/CLK _23490_/D VGND VGND VPWR VPWR _23490_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14918__A2 _14917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15040__B2 _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22441_ _22721_/A _22439_/X _21446_/X _22440_/X VGND VGND VPWR VPWR _22442_/A sky130_fd_sc_hd__o22a_4
XFILLER_167_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18524__A _18560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25160_ _23938_/CLK _14350_/X HRESETn VGND VGND VPWR VPWR _25160_/Q sky130_fd_sc_hd__dfrtp_4
X_22372_ _22365_/A _19071_/Y VGND VGND VPWR VPWR _22372_/X sky130_fd_sc_hd__or2_4
XFILLER_176_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24111_ _25538_/CLK _18907_/X HRESETn VGND VGND VPWR VPWR _17541_/A sky130_fd_sc_hd__dfrtp_4
X_21323_ _21323_/A VGND VGND VPWR VPWR _22932_/A sky130_fd_sc_hd__buf_2
X_25091_ _25091_/CLK _14584_/X HRESETn VGND VGND VPWR VPWR _13563_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_190_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16044__A _24727_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13354__A1 _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21254_ _21239_/A VGND VGND VPWR VPWR _22199_/A sky130_fd_sc_hd__buf_2
X_24042_ _24486_/CLK _20860_/Y HRESETn VGND VGND VPWR VPWR _24042_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24549__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20205_ _18033_/B VGND VGND VPWR VPWR _20205_/Y sky130_fd_sc_hd__inv_2
X_21185_ _21189_/A _21185_/B VGND VGND VPWR VPWR _21185_/X sky130_fd_sc_hd__or2_4
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20136_ _20136_/A _19898_/D _19803_/X VGND VGND VPWR VPWR _20137_/A sky130_fd_sc_hd__or3_4
XFILLER_77_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22377__B1 _14666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24131__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20067_ _20067_/A VGND VGND VPWR VPWR _20067_/X sky130_fd_sc_hd__buf_2
X_24944_ _25510_/CLK _24944_/D HRESETn VGND VGND VPWR VPWR _11670_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16056__B1 _16055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24875_ _24874_/CLK _15730_/X HRESETn VGND VGND VPWR VPWR _24875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_245_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11840_ _11840_/A VGND VGND VPWR VPWR _13669_/A sky130_fd_sc_hd__inv_2
X_23826_ _24089_/CLK _23826_/D VGND VGND VPWR VPWR _23826_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23324__B _16792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25337__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11768_/Y _11766_/X _11770_/X _11766_/X VGND VGND VPWR VPWR _11771_/X sky130_fd_sc_hd__a2bb2o_4
X_23757_ _23767_/CLK _19381_/X VGND VGND VPWR VPWR _18136_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _12010_/X _13506_/A VGND VGND VPWR VPWR _24097_/D sky130_fd_sc_hd__and2_4
XFILLER_54_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16219__A _22814_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13507_/Y _13509_/X VGND VGND VPWR VPWR _13510_/X sky130_fd_sc_hd__and2_4
XFILLER_202_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22708_ _22708_/A _22705_/X _22708_/C VGND VGND VPWR VPWR _22708_/X sky130_fd_sc_hd__and3_4
XFILLER_186_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _25111_/Q _14490_/B _14490_/C VGND VGND VPWR VPWR _14492_/B sky130_fd_sc_hd__or3_4
XPHY_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23688_ _23706_/CLK _19582_/X VGND VGND VPWR VPWR _19580_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13441_ _13293_/A _13437_/X _13441_/C VGND VGND VPWR VPWR _13441_/X sky130_fd_sc_hd__or3_4
X_25427_ _25428_/CLK _25427_/D HRESETn VGND VGND VPWR VPWR _25427_/Q sky130_fd_sc_hd__dfrtp_4
X_22639_ _22149_/X _22638_/X _22134_/A _25532_/Q _22554_/X VGND VGND VPWR VPWR _22639_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21104__A1 _24645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16160_ _16159_/Y _16155_/X _15976_/X _16155_/X VGND VGND VPWR VPWR _24683_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13372_ _13260_/A _13372_/B VGND VGND VPWR VPWR _13372_/X sky130_fd_sc_hd__or2_4
X_25358_ _25387_/CLK _25358_/D HRESETn VGND VGND VPWR VPWR _12342_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15111_ _24978_/Q _15110_/A _15296_/B _15110_/Y VGND VGND VPWR VPWR _15111_/X sky130_fd_sc_hd__o22a_4
XFILLER_154_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12323_ _12321_/A _24822_/Q _12321_/Y _12322_/Y VGND VGND VPWR VPWR _12327_/C sky130_fd_sc_hd__o22a_4
X_24309_ _25533_/CLK _17645_/X HRESETn VGND VGND VPWR VPWR _17523_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13578__A _15694_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16091_ _16084_/X VGND VGND VPWR VPWR _16111_/A sky130_fd_sc_hd__buf_2
XANTENNA__24972__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25289_ _24236_/CLK _13704_/X HRESETn VGND VGND VPWR VPWR _11832_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_119_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15042_ _15042_/A _15038_/X _15040_/X _15041_/X VGND VGND VPWR VPWR _15042_/X sky130_fd_sc_hd__or4_4
XFILLER_181_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12254_ _25463_/Q VGND VGND VPWR VPWR _12254_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24901__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16889__A _22190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19850_ _19849_/Y _19847_/X _19827_/X _19847_/X VGND VGND VPWR VPWR _23596_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24219__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12185_ _12184_/Y _21088_/A _12184_/Y _21088_/A VGND VGND VPWR VPWR _12185_/X sky130_fd_sc_hd__a2bb2o_4
X_18801_ _18793_/A _18801_/B _18801_/C VGND VGND VPWR VPWR _18801_/X sky130_fd_sc_hd__and3_4
X_19781_ _21243_/B _19776_/X _19091_/X _19764_/A VGND VGND VPWR VPWR _23619_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16993_ _16042_/Y _17034_/A _16042_/Y _17034_/A VGND VGND VPWR VPWR _16993_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18732_ _18732_/A _18732_/B VGND VGND VPWR VPWR _18734_/B sky130_fd_sc_hd__or2_4
X_15944_ _15931_/X VGND VGND VPWR VPWR _15944_/X sky130_fd_sc_hd__buf_2
XFILLER_48_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15875_ _15861_/X VGND VGND VPWR VPWR _15875_/X sky130_fd_sc_hd__buf_2
X_18663_ _16613_/Y _18683_/A _24516_/Q _18815_/A VGND VGND VPWR VPWR _18663_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14826_ _14826_/A VGND VGND VPWR VPWR _23993_/D sky130_fd_sc_hd__buf_2
X_17614_ _17614_/A _17628_/B _17545_/Y _17571_/X VGND VGND VPWR VPWR _17615_/B sky130_fd_sc_hd__or4_4
XFILLER_221_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18594_ _18587_/B VGND VGND VPWR VPWR _18595_/B sky130_fd_sc_hd__inv_2
XFILLER_224_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25078__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14757_ _25059_/Q _14769_/B _25060_/Q VGND VGND VPWR VPWR _14757_/X sky130_fd_sc_hd__and3_4
X_17545_ _24313_/Q VGND VGND VPWR VPWR _17545_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11969_ _11932_/B _11962_/X VGND VGND VPWR VPWR _11973_/A sky130_fd_sc_hd__and2_4
XANTENNA__16129__A _16124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25007__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13708_ _13666_/Y VGND VGND VPWR VPWR _13708_/X sky130_fd_sc_hd__buf_2
X_17476_ _17476_/A VGND VGND VPWR VPWR _17476_/X sky130_fd_sc_hd__buf_2
XFILLER_205_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14688_ _14688_/A VGND VGND VPWR VPWR _21911_/A sky130_fd_sc_hd__buf_2
XFILLER_204_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19215_ _23816_/Q VGND VGND VPWR VPWR _19215_/Y sky130_fd_sc_hd__inv_2
X_13639_ _24036_/Q _24035_/Q VGND VGND VPWR VPWR _13640_/B sky130_fd_sc_hd__nor2_4
X_16427_ _15072_/Y _16426_/X _16059_/X _16426_/X VGND VGND VPWR VPWR _24586_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23096__B2 _21051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16358_ _18951_/A VGND VGND VPWR VPWR _16358_/X sky130_fd_sc_hd__buf_2
X_19146_ _23841_/Q VGND VGND VPWR VPWR _19146_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15309_ _15338_/A _15307_/X _15308_/X VGND VGND VPWR VPWR _25007_/D sky130_fd_sc_hd__and3_4
XFILLER_118_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16289_ _23190_/A VGND VGND VPWR VPWR _16289_/Y sky130_fd_sc_hd__inv_2
X_19077_ _22215_/B _19074_/X _16864_/X _19074_/X VGND VGND VPWR VPWR _19077_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18028_ _14639_/A VGND VGND VPWR VPWR _18104_/A sky130_fd_sc_hd__buf_2
XFILLER_145_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24642__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18275__A1 _13772_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16286__B1 _15996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22313__B _22327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19979_ _19979_/A VGND VGND VPWR VPWR _21677_/B sky130_fd_sc_hd__inv_2
XFILLER_247_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22990_ _22786_/X _22988_/X _22789_/X _22989_/X VGND VGND VPWR VPWR _22991_/B sky130_fd_sc_hd__o22a_4
XFILLER_28_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21941_ _21466_/A _21941_/B VGND VGND VPWR VPWR _21942_/C sky130_fd_sc_hd__or2_4
XFILLER_227_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24660_ _24592_/CLK _16234_/X HRESETn VGND VGND VPWR VPWR _24660_/Q sky130_fd_sc_hd__dfrtp_4
X_21872_ _24789_/Q _21868_/X _23075_/C _24859_/Q _21871_/X VGND VGND VPWR VPWR _21872_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_243_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _23627_/CLK _23611_/D VGND VGND VPWR VPWR _13446_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__25430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _20823_/A _20823_/B VGND VGND VPWR VPWR _20824_/A sky130_fd_sc_hd__or2_4
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24591_ _24591_/CLK _24591_/D HRESETn VGND VGND VPWR VPWR _24591_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23542_ _23678_/CLK _20001_/X VGND VGND VPWR VPWR _23542_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20754_ _20754_/A VGND VGND VPWR VPWR _20754_/X sky130_fd_sc_hd__buf_2
XFILLER_168_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23473_ _23497_/CLK _23473_/D VGND VGND VPWR VPWR _23473_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20685_ _20685_/A _20685_/B VGND VGND VPWR VPWR _20686_/A sky130_fd_sc_hd__or2_4
XFILLER_210_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14782__A _18052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_24_0_HCLK clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_24_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25212_ _23951_/CLK _14165_/Y HRESETn VGND VGND VPWR VPWR _14154_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_195_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22424_ _20862_/A _22287_/X _13117_/A _21317_/X VGND VGND VPWR VPWR _22424_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25143_ _23958_/CLK _14409_/X HRESETn VGND VGND VPWR VPWR _20592_/A sky130_fd_sc_hd__dfstp_4
X_22355_ _22024_/A _22353_/X _22354_/X VGND VGND VPWR VPWR _22355_/X sky130_fd_sc_hd__and3_4
XFILLER_163_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21306_ _21303_/X _21305_/X _21306_/C VGND VGND VPWR VPWR _21306_/X sky130_fd_sc_hd__and3_4
XANTENNA__24383__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25074_ _23875_/CLK _14655_/Y HRESETn VGND VGND VPWR VPWR _13615_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15867__A3 _15719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22286_ _21099_/X VGND VGND VPWR VPWR _22286_/X sky130_fd_sc_hd__buf_2
XFILLER_151_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22598__B1 _24831_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24025_ _24060_/CLK _20788_/X HRESETn VGND VGND VPWR VPWR _13108_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__24312__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21237_ _25061_/Q VGND VGND VPWR VPWR _21262_/A sky130_fd_sc_hd__buf_2
XFILLER_78_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21168_ _15666_/A _21168_/B _21168_/C VGND VGND VPWR VPWR _21168_/X sky130_fd_sc_hd__and3_4
XANTENNA__17542__A1_N _11772_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_148_0_HCLK clkbuf_7_74_0_HCLK/X VGND VGND VPWR VPWR _25098_/CLK sky130_fd_sc_hd__clkbuf_1
X_20119_ _20118_/Y _20116_/X _20092_/X _20116_/X VGND VGND VPWR VPWR _20119_/X sky130_fd_sc_hd__a2bb2o_4
X_13990_ _13990_/A _13978_/A _13990_/C _13989_/X VGND VGND VPWR VPWR _14019_/C sky130_fd_sc_hd__or4_4
X_21099_ _22525_/A VGND VGND VPWR VPWR _21099_/X sky130_fd_sc_hd__buf_2
XANTENNA__25518__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12941_ _12941_/A VGND VGND VPWR VPWR _12941_/Y sky130_fd_sc_hd__inv_2
X_24927_ _25325_/CLK _24927_/D HRESETn VGND VGND VPWR VPWR _12050_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15660_ _15660_/A VGND VGND VPWR VPWR _15661_/A sky130_fd_sc_hd__buf_2
XANTENNA__17333__A _17333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12872_ _12872_/A _12872_/B _12871_/X VGND VGND VPWR VPWR _12873_/A sky130_fd_sc_hd__or3_4
X_24858_ _24855_/CLK _15765_/X HRESETn VGND VGND VPWR VPWR _24858_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_233_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15252__A1 _15246_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14610_/X VGND VGND VPWR VPWR _14611_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _11823_/A VGND VGND VPWR VPWR _11823_/Y sky130_fd_sc_hd__inv_2
X_23809_ _24413_/CLK _19236_/X VGND VGND VPWR VPWR _19235_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _24910_/Q VGND VGND VPWR VPWR _15591_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24789_ _24886_/CLK _24789_/D HRESETn VGND VGND VPWR VPWR _24789_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17338_/A _17328_/X _17330_/C VGND VGND VPWR VPWR _17330_/X sky130_fd_sc_hd__and3_4
XFILLER_81_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ HREADY HSEL VGND VGND VPWR VPWR _14542_/Y sky130_fd_sc_hd__nand2_4
XFILLER_202_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11752_/Y _11744_/X _11753_/X _11744_/X VGND VGND VPWR VPWR _11754_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21876__A2 _22136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15004__B2 _15003_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16201__B1 _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17261_/A VGND VGND VPWR VPWR _17261_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _21715_/A _14468_/X _14392_/X _14468_/X VGND VGND VPWR VPWR _25117_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ HWDATA[25] VGND VGND VPWR VPWR _11685_/X sky130_fd_sc_hd__buf_2
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16212_ _22939_/A VGND VGND VPWR VPWR _16212_/Y sky130_fd_sc_hd__inv_2
X_19000_ _17932_/B VGND VGND VPWR VPWR _19000_/Y sky130_fd_sc_hd__inv_2
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ _13392_/A _13424_/B VGND VGND VPWR VPWR _13425_/C sky130_fd_sc_hd__or2_4
X_17192_ _23253_/A _17273_/A _16283_/Y _17191_/Y VGND VGND VPWR VPWR _17192_/X sky130_fd_sc_hd__o22a_4
XFILLER_174_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16143_ _16140_/Y _16136_/X _16141_/X _16142_/X VGND VGND VPWR VPWR _16143_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13355_ _13186_/X _13354_/X _25329_/Q _13245_/X VGND VGND VPWR VPWR _13355_/X sky130_fd_sc_hd__o22a_4
XFILLER_6_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ _24828_/Q VGND VGND VPWR VPWR _12306_/Y sky130_fd_sc_hd__inv_2
X_16074_ _16073_/Y _15990_/A _15475_/X _15990_/A VGND VGND VPWR VPWR _16074_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15858__A3 _15702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13286_ _13389_/A _23855_/Q VGND VGND VPWR VPWR _13287_/C sky130_fd_sc_hd__or2_4
XFILLER_108_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15025_ _15025_/A VGND VGND VPWR VPWR _15025_/Y sky130_fd_sc_hd__inv_2
X_19902_ _19902_/A VGND VGND VPWR VPWR _19902_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24053__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12237_ _12273_/A VGND VGND VPWR VPWR _12443_/A sky130_fd_sc_hd__buf_2
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23250__A1 _24544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_44_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_44_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12541__A2 _24857_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19833_ _13732_/X _14683_/X _20136_/A _19898_/D VGND VGND VPWR VPWR _19833_/X sky130_fd_sc_hd__or4_4
XFILLER_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12168_ _12376_/A _23307_/A _12376_/A _23307_/A VGND VGND VPWR VPWR _12168_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19206__B1 _19138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19764_ _19764_/A VGND VGND VPWR VPWR _19764_/X sky130_fd_sc_hd__buf_2
X_12099_ _25474_/Q VGND VGND VPWR VPWR _12099_/Y sky130_fd_sc_hd__inv_2
X_16976_ _24723_/Q _24380_/Q _16054_/Y _16975_/Y VGND VGND VPWR VPWR _16976_/X sky130_fd_sc_hd__o22a_4
XFILLER_232_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18715_ _18707_/A _18713_/A VGND VGND VPWR VPWR _18715_/X sky130_fd_sc_hd__or2_4
X_15927_ _15923_/X _15887_/X _15702_/X _23307_/A _15926_/X VGND VGND VPWR VPWR _24779_/D
+ sky130_fd_sc_hd__a32o_4
X_19695_ _19691_/Y _19694_/X _19652_/X _19694_/X VGND VGND VPWR VPWR _23650_/D sky130_fd_sc_hd__a2bb2o_4
X_18646_ _16584_/Y _24140_/Q _16584_/Y _24140_/Q VGND VGND VPWR VPWR _18647_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15858_ _15843_/X _15850_/X _15702_/X _24816_/Q _15857_/X VGND VGND VPWR VPWR _15858_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_80_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14809_ _14809_/A _14809_/B _25047_/Q VGND VGND VPWR VPWR _14810_/B sky130_fd_sc_hd__or3_4
XFILLER_80_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18577_ _18577_/A _18577_/B VGND VGND VPWR VPWR _18578_/C sky130_fd_sc_hd__nand2_4
XANTENNA__12387__A _12204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15789_ _15783_/X VGND VGND VPWR VPWR _15789_/X sky130_fd_sc_hd__buf_2
XANTENNA__22513__B1 _21596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17528_ _25537_/Q _17646_/A _11768_/Y _17530_/A VGND VGND VPWR VPWR _17528_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24894__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17459_ _17459_/A _17487_/A VGND VGND VPWR VPWR _17472_/C sky130_fd_sc_hd__or2_4
XFILLER_177_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24823__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20470_ _20447_/C _20469_/X VGND VGND VPWR VPWR _20470_/X sky130_fd_sc_hd__or2_4
X_19129_ _19128_/Y _19126_/X _19057_/X _19126_/X VGND VGND VPWR VPWR _19129_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22140_ _22140_/A _22140_/B VGND VGND VPWR VPWR _22158_/C sky130_fd_sc_hd__and2_4
XFILLER_133_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22071_ _22199_/A VGND VGND VPWR VPWR _22387_/A sky130_fd_sc_hd__buf_2
XANTENNA__17418__A _14403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19445__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12850__A _12588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21022_ _21022_/A VGND VGND VPWR VPWR _22632_/A sky130_fd_sc_hd__buf_2
XANTENNA__13665__B _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22595__A3 _22135_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11740__B1 _11739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16274__A3 _16267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19633__A _18985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_1_0_HCLK clkbuf_5_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23155__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22973_ _21427_/A VGND VGND VPWR VPWR _22973_/X sky130_fd_sc_hd__buf_2
XFILLER_216_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13493__B1 _11770_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22752__B1 _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24712_ _24681_/CLK _24712_/D HRESETn VGND VGND VPWR VPWR _23316_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11689__A1_N _11687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21924_ _21924_/A VGND VGND VPWR VPWR _22343_/A sky130_fd_sc_hd__buf_2
XFILLER_216_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22994__A _23062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16431__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24643_ _24641_/CLK _24643_/D HRESETn VGND VGND VPWR VPWR _23313_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21855_ _21720_/A _21851_/X _21854_/X VGND VGND VPWR VPWR _21855_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_231_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22504__B1 _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _24030_/Q _20802_/X _20810_/B VGND VGND VPWR VPWR _20806_/Y sky130_fd_sc_hd__a21oi_4
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24574_ _24574_/CLK _16468_/X HRESETn VGND VGND VPWR VPWR _24574_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21858__A2 _21336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21786_ _21642_/X _21785_/X _13559_/Y _21642_/X VGND VGND VPWR VPWR _21786_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23525_ _23525_/CLK _23525_/D VGND VGND VPWR VPWR _23525_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20737_ _20731_/X _20733_/Y _15607_/A _20736_/X VGND VGND VPWR VPWR _20737_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23456_ _23456_/CLK _20228_/X VGND VGND VPWR VPWR _20226_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24564__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20668_ _17396_/A _17396_/B _17398_/A VGND VGND VPWR VPWR _20668_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22407_ _25527_/Q _22282_/X _21034_/X _22406_/X VGND VGND VPWR VPWR _22407_/X sky130_fd_sc_hd__a211o_4
XFILLER_167_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23387_ _23916_/CLK _20402_/X VGND VGND VPWR VPWR _23387_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_137_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20599_ _14394_/Y _18888_/A _18871_/A _18885_/A VGND VGND VPWR VPWR _20600_/B sky130_fd_sc_hd__o22a_4
XFILLER_125_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13140_ _13421_/A VGND VGND VPWR VPWR _13168_/A sky130_fd_sc_hd__buf_2
X_25126_ _23927_/CLK _25126_/D HRESETn VGND VGND VPWR VPWR _25126_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22338_ _21937_/A _22336_/X _22337_/X VGND VGND VPWR VPWR _22338_/X sky130_fd_sc_hd__and3_4
XFILLER_164_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13071_ _12979_/D _13091_/A VGND VGND VPWR VPWR _13072_/B sky130_fd_sc_hd__or2_4
X_25057_ _23735_/CLK _25057_/D HRESETn VGND VGND VPWR VPWR _25057_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19436__B1 _19414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22269_ _11808_/Y _21503_/X _21510_/A VGND VGND VPWR VPWR _22269_/X sky130_fd_sc_hd__a21o_4
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12022_ _12022_/A VGND VGND VPWR VPWR _12022_/Y sky130_fd_sc_hd__inv_2
X_24008_ _24037_/CLK _20712_/Y HRESETn VGND VGND VPWR VPWR _20709_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19987__B2 _19962_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11731__B1 _11730_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16830_ _16829_/Y _16827_/X _15743_/X _16827_/X VGND VGND VPWR VPWR _16830_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19543__A _19360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25352__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13973_ _13967_/Y _13969_/Y _14007_/C _14007_/D VGND VGND VPWR VPWR _13973_/X sky130_fd_sc_hd__and4_4
X_16761_ _16759_/Y _16755_/X _15741_/X _16760_/X VGND VGND VPWR VPWR _16761_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14687__A _22196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18500_ _18823_/B VGND VGND VPWR VPWR _18500_/X sky130_fd_sc_hd__buf_2
XFILLER_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12924_ _12889_/X _12924_/B _12924_/C VGND VGND VPWR VPWR _12924_/X sky130_fd_sc_hd__and3_4
X_15712_ _15736_/A VGND VGND VPWR VPWR _15759_/A sky130_fd_sc_hd__inv_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16692_ _16692_/A VGND VGND VPWR VPWR _16692_/X sky130_fd_sc_hd__buf_2
X_19480_ _19939_/A _18279_/X _19479_/X VGND VGND VPWR VPWR _19480_/X sky130_fd_sc_hd__or3_4
XFILLER_246_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18431_ _16235_/Y _18470_/A _16235_/Y _18470_/A VGND VGND VPWR VPWR _18431_/X sky130_fd_sc_hd__a2bb2o_4
X_12855_ _12845_/C _12852_/X _12847_/B _12854_/X VGND VGND VPWR VPWR _12855_/X sky130_fd_sc_hd__a211o_4
X_15643_ _13797_/A VGND VGND VPWR VPWR _15643_/X sky130_fd_sc_hd__buf_2
XFILLER_62_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17998__A _18095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _11806_/A VGND VGND VPWR VPWR _11806_/Y sky130_fd_sc_hd__inv_2
XPHY_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15574_ _15574_/A VGND VGND VPWR VPWR _15574_/Y sky130_fd_sc_hd__inv_2
X_18362_ _21983_/A _17476_/X _18361_/A _17480_/X VGND VGND VPWR VPWR _18363_/A sky130_fd_sc_hd__o22a_4
X_12786_ _25380_/Q VGND VGND VPWR VPWR _12786_/Y sky130_fd_sc_hd__inv_2
XPHY_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14525_/A VGND VGND VPWR VPWR _14525_/Y sky130_fd_sc_hd__inv_2
X_17313_ _17313_/A VGND VGND VPWR VPWR _24361_/D sky130_fd_sc_hd__inv_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11737_/A VGND VGND VPWR VPWR _11737_/Y sky130_fd_sc_hd__inv_2
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _24214_/Q VGND VGND VPWR VPWR _18296_/A sky130_fd_sc_hd__buf_2
XANTENNA__23231__C _22140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12935__A _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _14454_/Y _14455_/X _14384_/X _14455_/X VGND VGND VPWR VPWR _25124_/D sky130_fd_sc_hd__a2bb2o_4
X_17244_ _17185_/Y _17165_/Y _17240_/X _17243_/X VGND VGND VPWR VPWR _17244_/X sky130_fd_sc_hd__or4_4
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _11668_/A _11668_/B VGND VGND VPWR VPWR _11676_/A sky130_fd_sc_hd__or2_4
XFILLER_168_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _13234_/X _13407_/B VGND VGND VPWR VPWR _13407_/X sky130_fd_sc_hd__or2_4
X_17175_ _24368_/Q VGND VGND VPWR VPWR _17175_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24234__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14387_ _14386_/Y _14383_/X _14262_/X _14372_/X VGND VGND VPWR VPWR _14387_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16126_ _22753_/A VGND VGND VPWR VPWR _16126_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16489__B1 _16397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12373__C _12254_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13338_ _13434_/A _13338_/B _13337_/X VGND VGND VPWR VPWR _13338_/X sky130_fd_sc_hd__and3_4
XFILLER_127_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16690__A1_N _16689_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16057_ _24722_/Q VGND VGND VPWR VPWR _16057_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17238__A _21856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13269_ _13374_/A _19281_/A VGND VGND VPWR VPWR _13271_/B sky130_fd_sc_hd__or2_4
XANTENNA__19427__B1 _19357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16142__A _16124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15008_ _15008_/A VGND VGND VPWR VPWR _15008_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21234__B1 _21232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19816_ _19816_/A VGND VGND VPWR VPWR _19816_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25093__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_131_0_HCLK clkbuf_7_65_0_HCLK/X VGND VGND VPWR VPWR _23458_/CLK sky130_fd_sc_hd__clkbuf_1
X_19747_ _19740_/A VGND VGND VPWR VPWR _19747_/X sky130_fd_sc_hd__buf_2
X_16959_ _16009_/Y _24398_/Q _16009_/Y _24398_/Q VGND VGND VPWR VPWR _16959_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_194_0_HCLK clkbuf_7_97_0_HCLK/X VGND VGND VPWR VPWR _24654_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__25022__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19678_ _19672_/Y VGND VGND VPWR VPWR _19678_/X sky130_fd_sc_hd__buf_2
XANTENNA__12829__B _12759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18629_ _16571_/A _24145_/Q _16571_/Y _18693_/C VGND VGND VPWR VPWR _18637_/A sky130_fd_sc_hd__o22a_4
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21640_ _14711_/X _21632_/X _21639_/X VGND VGND VPWR VPWR _21640_/X sky130_fd_sc_hd__or3_4
XFILLER_212_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11789__B1 _25521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21571_ _21571_/A VGND VGND VPWR VPWR _21571_/X sky130_fd_sc_hd__buf_2
XANTENNA__12845__A _12769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23310_ _24816_/Q _23278_/B VGND VGND VPWR VPWR _23310_/X sky130_fd_sc_hd__or2_4
XFILLER_177_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20522_ _20522_/A _20448_/X VGND VGND VPWR VPWR _20522_/X sky130_fd_sc_hd__and2_4
XFILLER_165_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24290_ _24227_/CLK _24290_/D HRESETn VGND VGND VPWR VPWR _17704_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23241_ _22708_/A _23238_/X _23240_/X VGND VGND VPWR VPWR _23246_/C sky130_fd_sc_hd__and3_4
XFILLER_181_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20453_ _20444_/A _20450_/X _20453_/C _20453_/D VGND VGND VPWR VPWR _20453_/X sky130_fd_sc_hd__and4_4
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23172_ _23172_/A VGND VGND VPWR VPWR _23172_/X sky130_fd_sc_hd__buf_2
X_20384_ _20384_/A VGND VGND VPWR VPWR _20384_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22123_ _22122_/X VGND VGND VPWR VPWR _22123_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23957__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22054_ _22053_/X VGND VGND VPWR VPWR _22054_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20183__A2_N _20180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21005_ _21006_/A _14790_/A _21006_/C VGND VGND VPWR VPWR _21005_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_90_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_90_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15455__A1 _14269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11924__A _19617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22956_ _22844_/A _22956_/B _22956_/C VGND VGND VPWR VPWR _22956_/X sky130_fd_sc_hd__and3_4
XANTENNA__17314__C _17314_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21907_ _21911_/A _21905_/X _21906_/X VGND VGND VPWR VPWR _21907_/X sky130_fd_sc_hd__and3_4
XFILLER_244_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22887_ _16574_/A _22884_/X _22801_/X _22886_/X VGND VGND VPWR VPWR _22887_/X sky130_fd_sc_hd__a211o_4
XFILLER_71_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12640_ _12644_/A _12639_/X VGND VGND VPWR VPWR _12645_/B sky130_fd_sc_hd__or2_4
X_24626_ _24626_/CLK _16326_/X HRESETn VGND VGND VPWR VPWR _22710_/A sky130_fd_sc_hd__dfrtp_4
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21838_ _20517_/B _14183_/X _14254_/Y _14246_/A VGND VGND VPWR VPWR _21838_/X sky130_fd_sc_hd__o22a_4
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24745__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ _12569_/Y _24859_/Q _25429_/Q _12570_/Y VGND VGND VPWR VPWR _12577_/B sky130_fd_sc_hd__a2bb2o_4
X_24557_ _24555_/CLK _16511_/X HRESETn VGND VGND VPWR VPWR _16510_/A sky130_fd_sc_hd__dfrtp_4
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21769_ _21769_/A _21767_/X _21769_/C VGND VGND VPWR VPWR _21769_/X sky130_fd_sc_hd__and3_4
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _25172_/Q _14288_/Y _25171_/Q _14296_/A VGND VGND VPWR VPWR _14310_/X sky130_fd_sc_hd__o22a_4
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23508_ _23525_/CLK _23508_/D VGND VGND VPWR VPWR _20081_/A sky130_fd_sc_hd__dfxtp_4
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15290_ _24997_/Q VGND VGND VPWR VPWR _15351_/A sky130_fd_sc_hd__inv_2
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24488_ _24487_/CLK _16695_/X HRESETn VGND VGND VPWR VPWR _16694_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_183_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14241_ _14235_/Y _14240_/Y sda_oen_o_S5 _14235_/Y VGND VGND VPWR VPWR _14241_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23439_ _23534_/CLK _20273_/X VGND VGND VPWR VPWR _20271_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__15391__B1 _15334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14172_ _14161_/X _14170_/Y _14118_/X _14171_/Y _14115_/X VGND VGND VPWR VPWR _14172_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__11952__B1 _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13123_ _13122_/X VGND VGND VPWR VPWR _20793_/B sky130_fd_sc_hd__buf_2
X_25109_ _25109_/CLK _25109_/D HRESETn VGND VGND VPWR VPWR _20601_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13586__A _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19409__B1 _19408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18980_ HWDATA[6] VGND VGND VPWR VPWR _18981_/A sky130_fd_sc_hd__buf_2
XANTENNA__12490__A _12211_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25533__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13054_ _25350_/Q _13054_/B VGND VGND VPWR VPWR _13055_/C sky130_fd_sc_hd__or2_4
X_17931_ _13617_/X VGND VGND VPWR VPWR _17947_/A sky130_fd_sc_hd__buf_2
XFILLER_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12005_ _24097_/Q _12002_/A VGND VGND VPWR VPWR _12007_/A sky130_fd_sc_hd__and2_4
X_17862_ _17849_/X _17862_/B VGND VGND VPWR VPWR _17862_/X sky130_fd_sc_hd__or2_4
XANTENNA__15805__A1_N _12354_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19601_ _19596_/Y _19599_/X _19600_/X _19599_/X VGND VGND VPWR VPWR _23682_/D sky130_fd_sc_hd__a2bb2o_4
X_16813_ _16799_/A VGND VGND VPWR VPWR _16813_/X sky130_fd_sc_hd__buf_2
XANTENNA__21308__A _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17793_ _17793_/A _17787_/Y _17792_/X VGND VGND VPWR VPWR _17794_/A sky130_fd_sc_hd__or3_4
Xclkbuf_8_204_0_HCLK clkbuf_8_205_0_HCLK/A VGND VGND VPWR VPWR _24597_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19532_ _19530_/Y _19526_/X _19395_/X _19531_/X VGND VGND VPWR VPWR _23704_/D sky130_fd_sc_hd__a2bb2o_4
X_16744_ _16743_/Y _16739_/X _16391_/X _16739_/X VGND VGND VPWR VPWR _16744_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21027__B _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13956_ _13956_/A VGND VGND VPWR VPWR _13956_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12907_ _12907_/A VGND VGND VPWR VPWR _12907_/Y sky130_fd_sc_hd__inv_2
X_19463_ _19457_/Y VGND VGND VPWR VPWR _19463_/X sky130_fd_sc_hd__buf_2
X_13887_ _13907_/B VGND VGND VPWR VPWR _13887_/Y sky130_fd_sc_hd__inv_2
X_16675_ _24496_/Q VGND VGND VPWR VPWR _16675_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16946__B2 _24262_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18414_ _24654_/Q _24165_/Q _16249_/Y _18577_/A VGND VGND VPWR VPWR _18415_/D sky130_fd_sc_hd__o22a_4
X_12838_ _12838_/A _12838_/B _12766_/Y _12838_/D VGND VGND VPWR VPWR _12839_/D sky130_fd_sc_hd__or4_4
X_15626_ _15625_/Y _15622_/X _15466_/X _15622_/X VGND VGND VPWR VPWR _24897_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24486__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19394_ _18036_/B VGND VGND VPWR VPWR _19394_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18336__B _17448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18345_ _13162_/X _18344_/X _18342_/X VGND VGND VPWR VPWR _18345_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24415__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ _25397_/Q VGND VGND VPWR VPWR _12769_/Y sky130_fd_sc_hd__inv_2
X_15557_ HWDATA[29] VGND VGND VPWR VPWR _15557_/X sky130_fd_sc_hd__buf_2
XFILLER_187_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19896__B1 _19874_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14508_ _25108_/Q _14500_/X _25107_/Q _14502_/X VGND VGND VPWR VPWR _14508_/X sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_2_1_0_HCLK_A clkbuf_1_0_1_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15488_ _15541_/A _15486_/X HADDR[23] _15486_/X VGND VGND VPWR VPWR _15488_/X sky130_fd_sc_hd__a2bb2o_4
X_18276_ _24219_/Q VGND VGND VPWR VPWR _18276_/X sky130_fd_sc_hd__buf_2
X_17227_ _17227_/A _17227_/B _17221_/X _17227_/D VGND VGND VPWR VPWR _17228_/B sky130_fd_sc_hd__or4_4
X_14439_ _14166_/Y _14437_/X _14262_/X _14437_/X VGND VGND VPWR VPWR _14439_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21697__B _21601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12196__B1 _12194_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17158_ _17124_/X VGND VGND VPWR VPWR _17159_/B sky130_fd_sc_hd__inv_2
XFILLER_155_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16109_ _16108_/Y _16104_/X _15942_/X _16104_/X VGND VGND VPWR VPWR _24703_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17089_ _17031_/X _17097_/B VGND VGND VPWR VPWR _17090_/B sky130_fd_sc_hd__or2_4
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12499__B2 _24866_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22602__A _22602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_14_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__22955__B1 _22098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15437__A1 _14269_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23136__C _23135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22707__B1 _21730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22810_ _16444_/X _22806_/X _22810_/C VGND VGND VPWR VPWR _22811_/D sky130_fd_sc_hd__and3_4
XFILLER_72_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23790_ _23464_/CLK _23790_/D VGND VGND VPWR VPWR _23790_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22741_ _22741_/A _22532_/B VGND VGND VPWR VPWR _22744_/B sky130_fd_sc_hd__or2_4
XFILLER_26_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_1_HCLK clkbuf_1_0_1_HCLK/A VGND VGND VPWR VPWR clkbuf_1_0_1_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_25460_ _25453_/CLK _25460_/D HRESETn VGND VGND VPWR VPWR _12170_/A sky130_fd_sc_hd__dfrtp_4
X_22672_ _16829_/Y _22294_/X _21582_/X _22671_/X VGND VGND VPWR VPWR _22672_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24411_ _23610_/CLK _24411_/D HRESETn VGND VGND VPWR VPWR _24411_/Q sky130_fd_sc_hd__dfrtp_4
X_21623_ _22381_/A _21623_/B VGND VGND VPWR VPWR _21623_/X sky130_fd_sc_hd__or2_4
XANTENNA__24156__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25391_ _24809_/CLK _25391_/D HRESETn VGND VGND VPWR VPWR _12796_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_200_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16047__A _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24342_ _24172_/CLK _17380_/X HRESETn VGND VGND VPWR VPWR _17202_/A sky130_fd_sc_hd__dfrtp_4
X_21554_ _21549_/X _21551_/Y _21554_/C _21553_/X VGND VGND VPWR VPWR _21555_/B sky130_fd_sc_hd__and4_4
XFILLER_221_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20505_ _14053_/A _20449_/X VGND VGND VPWR VPWR _20505_/X sky130_fd_sc_hd__and2_4
X_24273_ _24278_/CLK _17837_/X HRESETn VGND VGND VPWR VPWR _17757_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19639__B1 _19587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21485_ _21809_/A _19893_/Y VGND VGND VPWR VPWR _21488_/B sky130_fd_sc_hd__or2_4
XFILLER_147_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23224_ _23223_/X VGND VGND VPWR VPWR _23224_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12726__A2 _12626_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20436_ _20444_/A _20440_/A VGND VGND VPWR VPWR _20436_/X sky130_fd_sc_hd__or2_4
XFILLER_106_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23155_ _22194_/A VGND VGND VPWR VPWR _23155_/X sky130_fd_sc_hd__buf_2
XANTENNA__11919__A _11897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20367_ _21179_/B _20362_/X _19874_/A _20349_/Y VGND VGND VPWR VPWR _23402_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22106_ _22105_/Y _21349_/A _14405_/Y _21351_/X VGND VGND VPWR VPWR _22107_/A sky130_fd_sc_hd__o22a_4
X_23086_ _21421_/A _23084_/Y _22831_/X _23085_/X VGND VGND VPWR VPWR _23087_/A sky130_fd_sc_hd__o22a_4
X_20298_ _21807_/B _20293_/X _19977_/X _20293_/X VGND VGND VPWR VPWR _23429_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21749__B2 _21598_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22037_ _22024_/A _22033_/X _22034_/X _22035_/X _22036_/X VGND VGND VPWR VPWR _22037_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_48_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16510__A _16510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22961__A3 _15855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24997__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11654__A _14364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13810_ _13810_/A VGND VGND VPWR VPWR _13810_/X sky130_fd_sc_hd__buf_2
X_14790_ _14790_/A VGND VGND VPWR VPWR _21006_/B sky130_fd_sc_hd__inv_2
XANTENNA__24926__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23988_ _25050_/CLK _23988_/D HRESETn VGND VGND VPWR VPWR _17399_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_217_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13741_ _13745_/A _13737_/X _20157_/C _13741_/D VGND VGND VPWR VPWR _20066_/A sky130_fd_sc_hd__or4_4
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22939_ _22939_/A _22729_/B VGND VGND VPWR VPWR _22939_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_34_0_HCLK clkbuf_8_35_0_HCLK/A VGND VGND VPWR VPWR _24413_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_204_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_18_0_HCLK_A clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13672_ _11823_/Y _13672_/B VGND VGND VPWR VPWR _13673_/B sky130_fd_sc_hd__or2_4
X_16460_ _16453_/A VGND VGND VPWR VPWR _16470_/A sky130_fd_sc_hd__buf_2
XFILLER_243_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_97_0_HCLK clkbuf_7_48_0_HCLK/X VGND VGND VPWR VPWR _24641_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_71_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12623_ _12623_/A _12623_/B VGND VGND VPWR VPWR _12625_/B sky130_fd_sc_hd__or2_4
X_15411_ _15296_/A _15410_/X VGND VGND VPWR VPWR _15411_/Y sky130_fd_sc_hd__nand2_4
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16391_ HWDATA[22] VGND VGND VPWR VPWR _16391_/X sky130_fd_sc_hd__buf_2
X_24609_ _24597_/CLK _16377_/X HRESETn VGND VGND VPWR VPWR _15104_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_43_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15342_ _15301_/X _15320_/D _15137_/Y VGND VGND VPWR VPWR _15342_/X sky130_fd_sc_hd__o21a_4
X_18130_ _18098_/A _18130_/B _18129_/X VGND VGND VPWR VPWR _18131_/C sky130_fd_sc_hd__and3_4
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12554_ _12553_/Y _24867_/Q _12553_/Y _24867_/Q VGND VGND VPWR VPWR _12557_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17353__A1 _17347_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12802__A1_N _12801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15273_ _15273_/A _15273_/B VGND VGND VPWR VPWR _15273_/X sky130_fd_sc_hd__or2_4
X_18061_ _18099_/A _18056_/X _18060_/X VGND VGND VPWR VPWR _18062_/C sky130_fd_sc_hd__or3_4
X_12485_ _12484_/X VGND VGND VPWR VPWR _12485_/Y sky130_fd_sc_hd__inv_2
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15903__A2 _15887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14224_ _25196_/Q VGND VGND VPWR VPWR _14224_/Y sky130_fd_sc_hd__inv_2
X_17012_ _16057_/Y _16957_/A _16067_/Y _17036_/A VGND VGND VPWR VPWR _17013_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21310__B _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14155_ _14111_/X _14087_/X _14087_/D _14154_/X VGND VGND VPWR VPWR _14155_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14205__A _20678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18900__A _18900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13106_ _24030_/Q _13106_/B VGND VGND VPWR VPWR _13124_/C sky130_fd_sc_hd__or2_4
XFILLER_4_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14086_ _14086_/A VGND VGND VPWR VPWR _14095_/A sky130_fd_sc_hd__inv_2
X_18963_ _18962_/Y _18960_/X _18942_/X _18960_/X VGND VGND VPWR VPWR _18963_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_239_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13037_ _13048_/A _13035_/X _13036_/X VGND VGND VPWR VPWR _25356_/D sky130_fd_sc_hd__and3_4
X_17914_ _17914_/A VGND VGND VPWR VPWR _17914_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18894_ _18871_/A _18885_/A _23952_/Q _20982_/B _18888_/A VGND VGND VPWR VPWR _18894_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16420__A HWDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16616__B1 _16435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17845_ _17818_/A _17843_/X _17845_/C VGND VGND VPWR VPWR _17845_/X sky130_fd_sc_hd__and3_4
XFILLER_94_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24667__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17776_ _17768_/C _17775_/X _16952_/X _17769_/Y VGND VGND VPWR VPWR _17776_/X sky130_fd_sc_hd__a211o_4
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14988_ _25036_/Q VGND VGND VPWR VPWR _14989_/A sky130_fd_sc_hd__inv_2
XFILLER_208_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22165__A1 _16605_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19515_ _19502_/Y VGND VGND VPWR VPWR _19515_/X sky130_fd_sc_hd__buf_2
X_16727_ _16723_/Y _16726_/X _15545_/X _16726_/X VGND VGND VPWR VPWR _16727_/X sky130_fd_sc_hd__a2bb2o_4
X_13939_ _13929_/Y _13939_/B _13936_/Y _13938_/X VGND VGND VPWR VPWR _13939_/X sky130_fd_sc_hd__or4_4
XFILLER_62_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17251__A _17179_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19446_ _19446_/A VGND VGND VPWR VPWR _19446_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16658_ _16657_/Y _16655_/X _16386_/X _16655_/X VGND VGND VPWR VPWR _24503_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15609_ _22566_/A _15608_/X _13818_/X _15608_/X VGND VGND VPWR VPWR _15609_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_5_0_HCLK clkbuf_5_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19377_ _18965_/A VGND VGND VPWR VPWR _19377_/X sky130_fd_sc_hd__buf_2
X_16589_ _16589_/A VGND VGND VPWR VPWR _16589_/Y sky130_fd_sc_hd__inv_2
X_18328_ _18328_/A VGND VGND VPWR VPWR _18328_/X sky130_fd_sc_hd__buf_2
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21501__A _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18259_ _11841_/Y _18252_/X _16849_/X _18236_/A VGND VGND VPWR VPWR _18259_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21270_ _21250_/A _20083_/Y VGND VGND VPWR VPWR _21270_/X sky130_fd_sc_hd__or2_4
XFILLER_116_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20221_ _20220_/X VGND VGND VPWR VPWR _20227_/A sky130_fd_sc_hd__inv_2
XANTENNA__21443__A3 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20152_ _23484_/Q VGND VGND VPWR VPWR _21401_/B sky130_fd_sc_hd__inv_2
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24960_ _24959_/CLK _15454_/X HRESETn VGND VGND VPWR VPWR _13902_/A sky130_fd_sc_hd__dfrtp_4
X_20083_ _20083_/A VGND VGND VPWR VPWR _20083_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16607__B1 _16522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21600__B1 _21596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23911_ _23452_/CLK _18943_/X VGND VGND VPWR VPWR _23911_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24891_ _24907_/CLK _15656_/X HRESETn VGND VGND VPWR VPWR _20822_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23842_ _24089_/CLK _23842_/D VGND VGND VPWR VPWR _19140_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23773_ _23889_/CLK _23773_/D VGND VGND VPWR VPWR _23773_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_250_0_HCLK clkbuf_8_251_0_HCLK/A VGND VGND VPWR VPWR _24340_/CLK sky130_fd_sc_hd__clkbuf_1
X_20985_ _20984_/A _20984_/B _24123_/Q _20984_/X VGND VGND VPWR VPWR _20985_/X sky130_fd_sc_hd__o22a_4
XPHY_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18257__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22724_ _22437_/A _22720_/X _23094_/A _22723_/Y VGND VGND VPWR VPWR _22724_/X sky130_fd_sc_hd__o22a_4
X_25512_ _24679_/CLK _25512_/D HRESETn VGND VGND VPWR VPWR _11848_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25443_ _25453_/CLK _12467_/Y HRESETn VGND VGND VPWR VPWR _25443_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22655_ _16539_/A _22654_/X _22138_/C _24833_/Q _22684_/B VGND VGND VPWR VPWR _22656_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15594__B1 _11726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21606_ _22225_/A VGND VGND VPWR VPWR _21756_/A sky130_fd_sc_hd__buf_2
X_25374_ _24795_/CLK _12952_/X HRESETn VGND VGND VPWR VPWR _25374_/Q sky130_fd_sc_hd__dfrtp_4
X_22586_ _20877_/Y _21597_/X _20738_/Y _22992_/A VGND VGND VPWR VPWR _22586_/X sky130_fd_sc_hd__o22a_4
XFILLER_138_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21131__A2 _21119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24325_ _24325_/CLK _17441_/X HRESETn VGND VGND VPWR VPWR _21012_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21411__A _22197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21537_ _22840_/A VGND VGND VPWR VPWR _21537_/X sky130_fd_sc_hd__buf_2
XFILLER_166_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12270_ _12208_/A _12191_/A _12267_/Y _12270_/D VGND VGND VPWR VPWR _12270_/X sky130_fd_sc_hd__or4_4
X_24256_ _24257_/CLK _24256_/D HRESETn VGND VGND VPWR VPWR _17893_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21468_ _21472_/A _21468_/B _21467_/X VGND VGND VPWR VPWR _21468_/X sky130_fd_sc_hd__and3_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23207_ _24574_/Q _23172_/X _23133_/X VGND VGND VPWR VPWR _23207_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25125__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20419_ _20419_/A VGND VGND VPWR VPWR _21762_/B sky130_fd_sc_hd__inv_2
X_24187_ _24675_/CLK _24187_/D HRESETn VGND VGND VPWR VPWR _24187_/Q sky130_fd_sc_hd__dfrtp_4
X_21399_ _21395_/X _21398_/X _14705_/A VGND VGND VPWR VPWR _21399_/X sky130_fd_sc_hd__o21a_4
XFILLER_135_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16846__B1 _16778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23138_ _23138_/A VGND VGND VPWR VPWR _23138_/X sky130_fd_sc_hd__buf_2
XFILLER_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15960_ _15955_/X _15958_/X _16229_/A _24762_/Q _15956_/X VGND VGND VPWR VPWR _24762_/D
+ sky130_fd_sc_hd__a32o_4
X_23069_ _24469_/Q _23002_/X _22891_/X VGND VGND VPWR VPWR _23069_/X sky130_fd_sc_hd__o21a_4
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16240__A _16240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14911_ _24422_/Q VGND VGND VPWR VPWR _14911_/Y sky130_fd_sc_hd__inv_2
X_15891_ _12773_/Y _15889_/X _15752_/X _15889_/X VGND VGND VPWR VPWR _15891_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_60_0_HCLK clkbuf_5_30_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_60_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_237_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17630_ _17543_/Y _17629_/X VGND VGND VPWR VPWR _17630_/X sky130_fd_sc_hd__or2_4
XFILLER_36_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14842_ _14842_/A VGND VGND VPWR VPWR _14842_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24760__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14624__A2 _14611_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17561_ _17561_/A VGND VGND VPWR VPWR _17561_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24078__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11985_ _11977_/A _11977_/B _11984_/Y VGND VGND VPWR VPWR _11985_/X sky130_fd_sc_hd__o21a_4
X_14773_ _14772_/X VGND VGND VPWR VPWR _14773_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22698__A2 _21596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19300_ _19299_/Y VGND VGND VPWR VPWR _19300_/X sky130_fd_sc_hd__buf_2
XFILLER_204_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16512_ _16512_/A VGND VGND VPWR VPWR _16512_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13724_ _13736_/A VGND VGND VPWR VPWR _13724_/X sky130_fd_sc_hd__buf_2
XFILLER_232_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24007__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17492_ _17590_/A _24114_/Q _17590_/A _24114_/Q VGND VGND VPWR VPWR _17497_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_232_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21305__B _21305_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19231_ _13723_/A _20157_/D _13743_/X _13745_/X VGND VGND VPWR VPWR _19232_/A sky130_fd_sc_hd__or4_4
XFILLER_220_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16443_ _22995_/A VGND VGND VPWR VPWR _21845_/A sky130_fd_sc_hd__buf_2
XFILLER_31_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13655_ _13655_/A _13655_/B VGND VGND VPWR VPWR _20823_/B sky130_fd_sc_hd__or2_4
XANTENNA__15585__B1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _12558_/Y _12553_/Y _12681_/B VGND VGND VPWR VPWR _12606_/X sky130_fd_sc_hd__or3_4
X_19162_ _19162_/A VGND VGND VPWR VPWR _19162_/Y sky130_fd_sc_hd__inv_2
X_13586_ _13586_/A VGND VGND VPWR VPWR _14648_/A sky130_fd_sc_hd__buf_2
X_16374_ _16372_/Y _16370_/X _16373_/X _16370_/X VGND VGND VPWR VPWR _24610_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18113_ _18113_/A _19444_/A VGND VGND VPWR VPWR _18113_/X sky130_fd_sc_hd__or2_4
X_12537_ _24864_/Q VGND VGND VPWR VPWR _12537_/Y sky130_fd_sc_hd__inv_2
X_15325_ _25003_/Q _15324_/Y VGND VGND VPWR VPWR _15327_/B sky130_fd_sc_hd__or2_4
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19093_ _23858_/Q VGND VGND VPWR VPWR _19093_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20330__B1 _19600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22136__B _22136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18044_ _18044_/A VGND VGND VPWR VPWR _18124_/A sky130_fd_sc_hd__buf_2
X_12468_ _12191_/X _12459_/X VGND VGND VPWR VPWR _12468_/X sky130_fd_sc_hd__or2_4
X_15256_ _25017_/Q _15256_/B VGND VGND VPWR VPWR _15256_/X sky130_fd_sc_hd__or2_4
X_14207_ _25201_/Q VGND VGND VPWR VPWR _14207_/Y sky130_fd_sc_hd__inv_2
X_15187_ _14995_/X _15064_/X _15242_/B VGND VGND VPWR VPWR _15187_/X sky130_fd_sc_hd__or3_4
X_12399_ _12277_/X _12378_/X _12278_/A VGND VGND VPWR VPWR _12399_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22622__A2 _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14138_ _14135_/X _14137_/Y _14417_/A _14135_/X VGND VGND VPWR VPWR _25219_/D sky130_fd_sc_hd__a2bb2o_4
X_19995_ _23544_/Q VGND VGND VPWR VPWR _22020_/B sky130_fd_sc_hd__inv_2
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22152__A _21439_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_235_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14069_ _23999_/Q _14058_/X _14062_/X _13979_/C _14065_/X VGND VGND VPWR VPWR _25235_/D
+ sky130_fd_sc_hd__a32o_4
X_18946_ _23909_/Q VGND VGND VPWR VPWR _18946_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16150__A _16124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24848__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18877_ _18877_/A _18876_/X VGND VGND VPWR VPWR _18877_/X sky130_fd_sc_hd__or2_4
XANTENNA__20397__B1 _15762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17828_ _17828_/A VGND VGND VPWR VPWR _17829_/B sky130_fd_sc_hd__inv_2
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24430__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17759_ _17757_/Y _17758_/Y _17817_/A _16938_/Y VGND VGND VPWR VPWR _17762_/C sky130_fd_sc_hd__or4_4
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13823__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18077__A _18054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20770_ _20753_/X _20769_/X _15588_/A _20757_/X VGND VGND VPWR VPWR _20770_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21215__B _21346_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19429_ _19428_/Y _19426_/X _19360_/X _19426_/X VGND VGND VPWR VPWR _19429_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_80_0_HCLK clkbuf_7_40_0_HCLK/X VGND VGND VPWR VPWR _25453_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_149_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13014__A _13028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22440_ _12757_/Y _21863_/X _22280_/X _12524_/Y _22294_/X VGND VGND VPWR VPWR _22440_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_222_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22310__A1 _24453_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22371_ _22367_/A _19251_/Y VGND VGND VPWR VPWR _22371_/X sky130_fd_sc_hd__or2_4
XFILLER_136_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20321__B1 _20061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24110_ _25538_/CLK _18908_/X HRESETn VGND VGND VPWR VPWR _24110_/Q sky130_fd_sc_hd__dfrtp_4
X_21322_ _16719_/A VGND VGND VPWR VPWR _23176_/A sky130_fd_sc_hd__buf_2
XFILLER_136_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_HCLK clkbuf_1_0_1_HCLK/X VGND VGND VPWR VPWR clkbuf_3_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_25090_ _24172_/CLK _25090_/D HRESETn VGND VGND VPWR VPWR _14548_/A sky130_fd_sc_hd__dfrtp_4
X_24041_ _24486_/CLK _24041_/D HRESETn VGND VGND VPWR VPWR _24041_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22074__B1 _14666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21253_ _21622_/A _21253_/B VGND VGND VPWR VPWR _21253_/X sky130_fd_sc_hd__or2_4
XFILLER_190_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20204_ _20203_/Y _20201_/X _19743_/X _20201_/X VGND VGND VPWR VPWR _23465_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16828__B1 _15741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21821__B1 _21501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21184_ _21205_/A _21184_/B VGND VGND VPWR VPWR _21184_/X sky130_fd_sc_hd__or2_4
XFILLER_116_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20135_ _23490_/Q VGND VGND VPWR VPWR _20135_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15500__B1 HADDR[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24589__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20066_ _20066_/A VGND VGND VPWR VPWR _20067_/A sky130_fd_sc_hd__inv_2
X_24943_ _25510_/CLK _15497_/X HRESETn VGND VGND VPWR VPWR _15496_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24518__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_4_0_HCLK_A clkbuf_3_5_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24874_ _24874_/CLK _24874_/D HRESETn VGND VGND VPWR VPWR _12521_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_57_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21406__A _22196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24171__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23825_ _23831_/CLK _23825_/D VGND VGND VPWR VPWR _18018_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__13814__B1 _11739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17005__B1 _24736_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24100__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _13829_/A VGND VGND VPWR VPWR _11770_/X sky130_fd_sc_hd__buf_2
X_23756_ _23767_/CLK _23756_/D VGND VGND VPWR VPWR _18168_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ _20968_/A _13506_/A VGND VGND VPWR VPWR _24096_/D sky130_fd_sc_hd__and2_4
XFILLER_198_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21352__A2 _21351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _24529_/Q _22416_/B _21730_/A _22706_/X VGND VGND VPWR VPWR _22708_/C sky130_fd_sc_hd__a211o_4
XFILLER_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23687_ _23706_/CLK _23687_/D VGND VGND VPWR VPWR _21969_/D sky130_fd_sc_hd__dfxtp_4
XPHY_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20899_ _24051_/Q _20921_/C VGND VGND VPWR VPWR _20899_/X sky130_fd_sc_hd__or2_4
XPHY_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13231_/X _13438_/X _13439_/X VGND VGND VPWR VPWR _13441_/C sky130_fd_sc_hd__and3_4
XANTENNA__25377__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22638_ _22638_/A _22638_/B VGND VGND VPWR VPWR _22638_/X sky130_fd_sc_hd__or2_4
X_25426_ _24872_/CLK _12643_/X HRESETn VGND VGND VPWR VPWR _25426_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_108_0_HCLK clkbuf_7_54_0_HCLK/X VGND VGND VPWR VPWR _24626_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_186_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22301__B2 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25306__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13371_ _13264_/X _13371_/B VGND VGND VPWR VPWR _13371_/X sky130_fd_sc_hd__or2_4
X_25357_ _25387_/CLK _25357_/D HRESETn VGND VGND VPWR VPWR _25357_/Q sky130_fd_sc_hd__dfrtp_4
X_22569_ _22758_/A _22569_/B VGND VGND VPWR VPWR _22569_/Y sky130_fd_sc_hd__nor2_4
XFILLER_155_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22852__A2 _22850_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12322_ _24822_/Q VGND VGND VPWR VPWR _12322_/Y sky130_fd_sc_hd__inv_2
X_15110_ _15110_/A VGND VGND VPWR VPWR _15110_/Y sky130_fd_sc_hd__inv_2
X_16090_ _24710_/Q VGND VGND VPWR VPWR _16090_/Y sky130_fd_sc_hd__inv_2
X_24308_ _25533_/CLK _17647_/X HRESETn VGND VGND VPWR VPWR _24308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25288_ _25292_/CLK _25288_/D HRESETn VGND VGND VPWR VPWR _11814_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20980__A scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15041_ _14898_/X _15020_/Y _14886_/A _15010_/Y VGND VGND VPWR VPWR _15041_/X sky130_fd_sc_hd__a2bb2o_4
X_12253_ _12252_/X _24751_/Q _12268_/A _12219_/Y VGND VGND VPWR VPWR _12253_/X sky130_fd_sc_hd__a2bb2o_4
X_24239_ _24341_/CLK _24239_/D HRESETn VGND VGND VPWR VPWR _11844_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22065__B1 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16819__B1 HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23068__A _24603_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12184_ _21078_/A VGND VGND VPWR VPWR _12184_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18800_ _18789_/A _18798_/A VGND VGND VPWR VPWR _18801_/C sky130_fd_sc_hd__or2_4
XANTENNA__15098__A2 _24604_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19780_ _23619_/Q VGND VGND VPWR VPWR _21243_/B sky130_fd_sc_hd__inv_2
XANTENNA__24941__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16992_ _24717_/Q _17041_/C _24721_/Q _16991_/Y VGND VGND VPWR VPWR _16995_/B sky130_fd_sc_hd__a2bb2o_4
X_18731_ _18733_/B VGND VGND VPWR VPWR _18732_/B sky130_fd_sc_hd__inv_2
XFILLER_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15943_ _12247_/Y _15935_/X _15942_/X _15935_/X VGND VGND VPWR VPWR _24770_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24259__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18662_ _18655_/X _18662_/B _18662_/C _18661_/X VGND VGND VPWR VPWR _18669_/C sky130_fd_sc_hd__or4_4
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15874_ _12810_/Y _15872_/X _11711_/X _15872_/X VGND VGND VPWR VPWR _24805_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23317__B1 _24114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17613_ _17613_/A VGND VGND VPWR VPWR _17613_/Y sky130_fd_sc_hd__inv_2
X_14825_ _14820_/X _14824_/X _25055_/Q _14820_/X VGND VGND VPWR VPWR _14825_/X sky130_fd_sc_hd__a2bb2o_4
X_18593_ _18593_/A _18592_/Y _18593_/C VGND VGND VPWR VPWR _18593_/X sky130_fd_sc_hd__and3_4
XFILLER_221_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17544_ _17585_/A _25546_/Q _11710_/A _17543_/Y VGND VGND VPWR VPWR _17544_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_233_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14756_ _14756_/A VGND VGND VPWR VPWR _14758_/B sky130_fd_sc_hd__inv_2
X_11968_ _11932_/C _11967_/X _11965_/X VGND VGND VPWR VPWR _11968_/X sky130_fd_sc_hd__o21a_4
XFILLER_72_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13707_ _11810_/Y _13673_/B VGND VGND VPWR VPWR _13707_/Y sky130_fd_sc_hd__nand2_4
XFILLER_204_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15558__B1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17475_ _17480_/A VGND VGND VPWR VPWR _17476_/A sky130_fd_sc_hd__inv_2
XFILLER_189_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11899_ _11895_/Y _11898_/X RsRx_S1 _11898_/X VGND VGND VPWR VPWR _25510_/D sky130_fd_sc_hd__a2bb2o_4
X_14687_ _22196_/A VGND VGND VPWR VPWR _14688_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_67_0_HCLK clkbuf_7_67_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_19214_ _19213_/Y _19211_/X _19122_/X _19211_/X VGND VGND VPWR VPWR _19214_/X sky130_fd_sc_hd__a2bb2o_4
X_16426_ _16418_/A VGND VGND VPWR VPWR _16426_/X sky130_fd_sc_hd__buf_2
XFILLER_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13638_ _13638_/A VGND VGND VPWR VPWR _13640_/A sky130_fd_sc_hd__inv_2
XANTENNA__14230__B1 _13798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23096__A2 _22559_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22147__A _15704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21051__A _21051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25047__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19145_ _19140_/Y _19143_/X _19144_/X _19143_/X VGND VGND VPWR VPWR _23842_/D sky130_fd_sc_hd__a2bb2o_4
X_16357_ _24613_/Q VGND VGND VPWR VPWR _16357_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13569_ _13569_/A VGND VGND VPWR VPWR _14552_/A sky130_fd_sc_hd__inv_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22843__A2 _22838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16145__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15308_ _15070_/Y _15308_/B VGND VGND VPWR VPWR _15308_/X sky130_fd_sc_hd__or2_4
XFILLER_185_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19076_ _19076_/A VGND VGND VPWR VPWR _22215_/B sky130_fd_sc_hd__inv_2
XANTENNA__16996__A1_N _16040_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16288_ _16287_/Y _16285_/X _16001_/X _16285_/X VGND VGND VPWR VPWR _24640_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18027_ _18027_/A _23768_/Q VGND VGND VPWR VPWR _18030_/B sky130_fd_sc_hd__or2_4
X_15239_ _15204_/B _15233_/X _15194_/X _15236_/B VGND VGND VPWR VPWR _15240_/A sky130_fd_sc_hd__a211o_4
XANTENNA__15730__B1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19978_ _19976_/Y _19971_/X _19977_/X _19971_/X VGND VGND VPWR VPWR _23550_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24682__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18929_ _23915_/Q VGND VGND VPWR VPWR _18929_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24611__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_HCLK HCLK VGND VGND VPWR VPWR clkbuf_0_HCLK/X sky130_fd_sc_hd__clkbuf_16
X_21940_ _21463_/A _21940_/B VGND VGND VPWR VPWR _21940_/X sky130_fd_sc_hd__or2_4
XFILLER_82_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21226__A _22829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21871_ _23171_/A VGND VGND VPWR VPWR _21871_/X sky130_fd_sc_hd__buf_2
XFILLER_242_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15797__B1 _15564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23610_ _23610_/CLK _23610_/D VGND VGND VPWR VPWR _23610_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11752__A _25529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20822_ _20822_/A VGND VGND VPWR VPWR _20823_/A sky130_fd_sc_hd__inv_2
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24590_ _24597_/CLK _24590_/D HRESETn VGND VGND VPWR VPWR _24590_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23541_ _23411_/CLK _20004_/X VGND VGND VPWR VPWR _23541_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20753_ _20780_/A VGND VGND VPWR VPWR _20753_/X sky130_fd_sc_hd__buf_2
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15013__A2 _24476_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23472_ _23490_/CLK _20186_/X VGND VGND VPWR VPWR _20184_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20684_ _20684_/A VGND VGND VPWR VPWR _20685_/A sky130_fd_sc_hd__inv_2
XANTENNA__14221__B1 _13785_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25211_ _25211_/CLK _14169_/Y HRESETn VGND VGND VPWR VPWR _14162_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22423_ _22423_/A VGND VGND VPWR VPWR _22423_/X sky130_fd_sc_hd__buf_2
XFILLER_210_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16055__A _14400_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25142_ _23958_/CLK _14411_/X HRESETn VGND VGND VPWR VPWR _25142_/Q sky130_fd_sc_hd__dfstp_4
X_22354_ _22020_/A _19596_/Y VGND VGND VPWR VPWR _22354_/X sky130_fd_sc_hd__or2_4
XANTENNA__21896__A _22069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21305_ _24480_/Q _21305_/B VGND VGND VPWR VPWR _21305_/X sky130_fd_sc_hd__or2_4
XFILLER_136_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25073_ _25073_/CLK _14657_/X HRESETn VGND VGND VPWR VPWR _25073_/Q sky130_fd_sc_hd__dfrtp_4
X_22285_ _22725_/A _22284_/Y VGND VGND VPWR VPWR _22285_/Y sky130_fd_sc_hd__nor2_4
X_24024_ _24060_/CLK _20785_/X HRESETn VGND VGND VPWR VPWR _20781_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22598__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21236_ _21225_/Y _21119_/X _21227_/X _21235_/X VGND VGND VPWR VPWR _21286_/C sky130_fd_sc_hd__a211o_4
XFILLER_116_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11927__A _19620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21167_ _16536_/Y _21583_/A _11701_/X _21166_/X VGND VGND VPWR VPWR _21168_/C sky130_fd_sc_hd__a211o_4
X_20118_ _20118_/A VGND VGND VPWR VPWR _20118_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24352__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21098_ _21098_/A VGND VGND VPWR VPWR _21098_/X sky130_fd_sc_hd__buf_2
XFILLER_93_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22520__A _22520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12940_ _12756_/X _12931_/X VGND VGND VPWR VPWR _12941_/A sky130_fd_sc_hd__or2_4
X_20049_ _20048_/Y _20046_/X _19827_/X _20046_/X VGND VGND VPWR VPWR _23524_/D sky130_fd_sc_hd__a2bb2o_4
X_24926_ _23378_/CLK _15536_/X HRESETn VGND VGND VPWR VPWR _13581_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_86_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12871_ _12842_/B _12851_/B _12744_/Y VGND VGND VPWR VPWR _12871_/X sky130_fd_sc_hd__o21a_4
X_24857_ _25403_/CLK _15766_/X HRESETn VGND VGND VPWR VPWR _24857_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14610_/A _14610_/B VGND VGND VPWR VPWR _14610_/X sky130_fd_sc_hd__or2_4
XFILLER_215_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11822_ _11815_/X _11817_/X _11822_/C _11822_/D VGND VGND VPWR VPWR _11847_/B sky130_fd_sc_hd__or4_4
X_23808_ _23808_/CLK _19239_/X VGND VGND VPWR VPWR _23808_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _22878_/A _15584_/X _11718_/X _15589_/X VGND VGND VPWR VPWR _24911_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13580__C _11659_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24788_ _24886_/CLK _15899_/X HRESETn VGND VGND VPWR VPWR _24788_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14460__B1 _14389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ HWDATA[9] VGND VGND VPWR VPWR _11753_/X sky130_fd_sc_hd__buf_2
X_14541_ _14540_/X VGND VGND VPWR VPWR _23339_/A sky130_fd_sc_hd__buf_2
XFILLER_121_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23739_ _25073_/CLK _23739_/D VGND VGND VPWR VPWR _18207_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_198_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21876__A3 _22816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17261_/A _17260_/B VGND VGND VPWR VPWR _17263_/B sky130_fd_sc_hd__or2_4
XFILLER_42_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11683_/X VGND VGND VPWR VPWR _11684_/X sky130_fd_sc_hd__buf_2
X_14472_ _25117_/Q VGND VGND VPWR VPWR _21715_/A sky130_fd_sc_hd__inv_2
XFILLER_186_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _16209_/Y _16210_/X _16020_/X _16210_/X VGND VGND VPWR VPWR _16211_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _13391_/A _23811_/Q VGND VGND VPWR VPWR _13425_/B sky130_fd_sc_hd__or2_4
X_25409_ _25409_/CLK _25409_/D HRESETn VGND VGND VPWR VPWR _25409_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17191_ _17273_/A VGND VGND VPWR VPWR _17191_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15960__B1 _24762_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13354_ _11951_/X _13338_/X _13353_/X _25330_/Q _13243_/X VGND VGND VPWR VPWR _13354_/X
+ sky130_fd_sc_hd__o32a_4
X_16142_ _16124_/A VGND VGND VPWR VPWR _16142_/X sky130_fd_sc_hd__buf_2
XFILLER_167_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12305_ _12305_/A VGND VGND VPWR VPWR _13073_/A sky130_fd_sc_hd__inv_2
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13285_ _13285_/A _23871_/Q VGND VGND VPWR VPWR _13285_/X sky130_fd_sc_hd__or2_4
X_16073_ _24716_/Q VGND VGND VPWR VPWR _16073_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18180__A _18052_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12236_ _12236_/A VGND VGND VPWR VPWR _12273_/A sky130_fd_sc_hd__inv_2
X_15024_ _25012_/Q _15022_/Y _25014_/Q _15023_/Y VGND VGND VPWR VPWR _15024_/X sky130_fd_sc_hd__a2bb2o_4
X_19901_ _22386_/B _19900_/X _19807_/X _19900_/X VGND VGND VPWR VPWR _23578_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_4_9_0_HCLK clkbuf_3_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__23250__A2 _22282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19832_ _25280_/Q VGND VGND VPWR VPWR _20136_/A sky130_fd_sc_hd__buf_2
XFILLER_111_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12167_ _12167_/A VGND VGND VPWR VPWR _12376_/A sky130_fd_sc_hd__inv_2
XFILLER_123_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19763_ _19763_/A VGND VGND VPWR VPWR _19764_/A sky130_fd_sc_hd__inv_2
XANTENNA__24093__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12098_ _12097_/Y _12095_/X _11765_/X _12095_/X VGND VGND VPWR VPWR _12098_/X sky130_fd_sc_hd__a2bb2o_4
X_16975_ _24380_/Q VGND VGND VPWR VPWR _16975_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22430__A _22429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18714_ _24155_/Q _18714_/B VGND VGND VPWR VPWR _18714_/X sky130_fd_sc_hd__or2_4
X_15926_ _15925_/X VGND VGND VPWR VPWR _15926_/X sky130_fd_sc_hd__buf_2
XFILLER_232_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24022__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19694_ _19694_/A VGND VGND VPWR VPWR _19694_/X sky130_fd_sc_hd__buf_2
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_30_0_HCLK clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_30_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18645_ _16589_/Y _24138_/Q _16589_/Y _24138_/Q VGND VGND VPWR VPWR _18645_/X sky130_fd_sc_hd__a2bb2o_4
X_15857_ _15857_/A VGND VGND VPWR VPWR _15857_/X sky130_fd_sc_hd__buf_2
XFILLER_92_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14808_ _23994_/Q _14808_/B _14808_/C VGND VGND VPWR VPWR _14809_/B sky130_fd_sc_hd__or3_4
XANTENNA__25299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18576_ _18572_/A _18567_/B _18575_/Y VGND VGND VPWR VPWR _24166_/D sky130_fd_sc_hd__and3_4
X_15788_ _15777_/X _15784_/X _15702_/X _24851_/Q _15787_/X VGND VGND VPWR VPWR _24851_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_224_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14451__B1 _14380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22513__A1 _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17527_ _24308_/Q VGND VGND VPWR VPWR _17646_/A sky130_fd_sc_hd__inv_2
XANTENNA__25228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14739_ _21787_/A _14697_/A _14699_/B VGND VGND VPWR VPWR _14739_/X sky130_fd_sc_hd__o21a_4
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19390__B1 _19301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17458_ _18326_/C _13157_/X _18326_/C _13157_/X VGND VGND VPWR VPWR _17487_/A sky130_fd_sc_hd__a2bb2o_4
X_16409_ _16408_/Y _16406_/X _16226_/X _16406_/X VGND VGND VPWR VPWR _24595_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22277__B1 _24826_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17389_ _23980_/Q _17389_/B VGND VGND VPWR VPWR _20640_/A sky130_fd_sc_hd__or2_4
XFILLER_146_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19128_ _19128_/A VGND VGND VPWR VPWR _19128_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_154_0_HCLK clkbuf_7_77_0_HCLK/X VGND VGND VPWR VPWR _25479_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__22605__A _16689_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19059_ _23870_/Q VGND VGND VPWR VPWR _19059_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24863__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18090__A _18090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16603__A _24522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22070_ _22367_/A _22070_/B VGND VGND VPWR VPWR _22070_/X sky130_fd_sc_hd__or2_4
XFILLER_160_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21021_ _21021_/A VGND VGND VPWR VPWR _21022_/A sky130_fd_sc_hd__buf_2
XANTENNA__11747__A HWDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22972_ _22972_/A _22901_/B VGND VGND VPWR VPWR _22972_/X sky130_fd_sc_hd__or2_4
XFILLER_101_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18956__B1 _17415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24711_ _24681_/CLK _16089_/X HRESETn VGND VGND VPWR VPWR _24711_/Q sky130_fd_sc_hd__dfrtp_4
X_21923_ _21207_/A VGND VGND VPWR VPWR _21933_/A sky130_fd_sc_hd__buf_2
XFILLER_243_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21854_ _21575_/X _21852_/X _21569_/X _21853_/X VGND VGND VPWR VPWR _21854_/X sky130_fd_sc_hd__o22a_4
X_24642_ _24641_/CLK _16282_/X HRESETn VGND VGND VPWR VPWR _24642_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_222_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20805_ _20805_/A VGND VGND VPWR VPWR _20810_/B sky130_fd_sc_hd__inv_2
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23171__A _23171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21785_ _21643_/X _21784_/X _25274_/Q _18263_/X VGND VGND VPWR VPWR _21785_/X sky130_fd_sc_hd__o22a_4
X_24573_ _24573_/CLK _16471_/X HRESETn VGND VGND VPWR VPWR _16469_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19381__B1 _19357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20736_ _20735_/X VGND VGND VPWR VPWR _20736_/X sky130_fd_sc_hd__buf_2
X_23524_ _23525_/CLK _23524_/D VGND VGND VPWR VPWR _23524_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_50_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23455_ _23456_/CLK _23455_/D VGND VGND VPWR VPWR _23455_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20667_ _20667_/A _20664_/X _20666_/X VGND VGND VPWR VPWR _20667_/X sky130_fd_sc_hd__and3_4
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22406_ _22821_/B _22405_/X _22296_/X VGND VGND VPWR VPWR _22406_/X sky130_fd_sc_hd__and3_4
X_23386_ _23916_/CLK _23386_/D VGND VGND VPWR VPWR _13395_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_109_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20598_ _20598_/A VGND VGND VPWR VPWR _20598_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22283__A3 _21306_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22337_ _21466_/A _22337_/B VGND VGND VPWR VPWR _22337_/X sky130_fd_sc_hd__or2_4
X_25125_ _23927_/CLK _14453_/X HRESETn VGND VGND VPWR VPWR _25125_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13070_ _12330_/Y _13089_/A VGND VGND VPWR VPWR _13091_/A sky130_fd_sc_hd__or2_4
X_25056_ _25056_/CLK _25056_/D HRESETn VGND VGND VPWR VPWR _25056_/Q sky130_fd_sc_hd__dfrtp_4
X_22268_ _22268_/A VGND VGND VPWR VPWR _22268_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24533__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12021_ _12019_/Y _12015_/X _12022_/A _12020_/X VGND VGND VPWR VPWR _25493_/D sky130_fd_sc_hd__a2bb2o_4
X_24007_ _24037_/CLK _24007_/D HRESETn VGND VGND VPWR VPWR _13114_/A sky130_fd_sc_hd__dfrtp_4
X_21219_ _13804_/Y _21218_/Y _24226_/Q _13804_/Y VGND VGND VPWR VPWR _21219_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22440__B1 _12524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22199_ _22199_/A _20036_/Y VGND VGND VPWR VPWR _22200_/C sky130_fd_sc_hd__or2_4
XANTENNA__23991__D sda_i_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22888__C _22887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15467__A1_N _15465_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16760_ _16766_/A VGND VGND VPWR VPWR _16760_/X sky130_fd_sc_hd__buf_2
X_13972_ _13991_/B VGND VGND VPWR VPWR _14007_/D sky130_fd_sc_hd__buf_2
XFILLER_59_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15711_ _15540_/X _15709_/X _15710_/X _24885_/Q _15707_/X VGND VGND VPWR VPWR _15711_/X
+ sky130_fd_sc_hd__a32o_4
X_12923_ _22667_/A _12920_/X VGND VGND VPWR VPWR _12924_/C sky130_fd_sc_hd__or2_4
X_24909_ _24910_/CLK _15594_/X HRESETn VGND VGND VPWR VPWR _15593_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_206_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16691_ _24489_/Q VGND VGND VPWR VPWR _16691_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18430_ _21335_/A _18561_/C _22097_/A _18563_/A VGND VGND VPWR VPWR _18433_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25392__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15642_ _21296_/A VGND VGND VPWR VPWR _15642_/X sky130_fd_sc_hd__buf_2
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12854_ _12887_/A VGND VGND VPWR VPWR _12854_/X sky130_fd_sc_hd__buf_2
XPHY_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25321__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11803_/Y _24230_/Q _13678_/A _24237_/Q VGND VGND VPWR VPWR _11805_/X sky130_fd_sc_hd__a2bb2o_4
X_18361_ _18361_/A VGND VGND VPWR VPWR _21983_/A sky130_fd_sc_hd__inv_2
XPHY_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15572_/Y _15570_/X _11688_/X _15570_/X VGND VGND VPWR VPWR _24917_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _25369_/Q _12783_/Y _25373_/Q _12784_/Y VGND VGND VPWR VPWR _12792_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17249_/D _17307_/B _17276_/X _17309_/B VGND VGND VPWR VPWR _17313_/A sky130_fd_sc_hd__a211o_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14523_/A VGND VGND VPWR VPWR _14524_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11736_ _11732_/Y _11733_/X _11735_/X _11733_/X VGND VGND VPWR VPWR _11736_/X sky130_fd_sc_hd__a2bb2o_4
X_18292_ _21822_/A _18283_/X _17703_/X VGND VGND VPWR VPWR _18292_/X sky130_fd_sc_hd__a21o_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16186__B1 _15991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _17193_/Y _17243_/B _17171_/Y _17344_/A VGND VGND VPWR VPWR _17243_/X sky130_fd_sc_hd__or4_4
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _14455_/A VGND VGND VPWR VPWR _14455_/X sky130_fd_sc_hd__buf_2
XANTENNA__15933__B1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15311__B _15311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11667_ _11667_/A _11667_/B VGND VGND VPWR VPWR _11668_/B sky130_fd_sc_hd__or2_4
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14208__A _14208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _13438_/A _23788_/Q VGND VGND VPWR VPWR _13406_/X sky130_fd_sc_hd__or2_4
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17174_ _17174_/A VGND VGND VPWR VPWR _17249_/C sky130_fd_sc_hd__inv_2
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14386_ _25148_/Q VGND VGND VPWR VPWR _14386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17416__A2_N _17414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_227_0_HCLK clkbuf_8_227_0_HCLK/A VGND VGND VPWR VPWR _25204_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_127_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16125_ _16122_/Y _16124_/X _11726_/X _16124_/X VGND VGND VPWR VPWR _24697_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13337_ _13369_/A _13333_/X _13336_/X VGND VGND VPWR VPWR _13337_/X sky130_fd_sc_hd__or3_4
XFILLER_227_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16056_ _16054_/Y _16050_/X _16055_/X _16050_/X VGND VGND VPWR VPWR _24723_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24274__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13268_ _13397_/A VGND VGND VPWR VPWR _13268_/X sky130_fd_sc_hd__buf_2
X_15007_ _14999_/X _15007_/B _15007_/C _15007_/D VGND VGND VPWR VPWR _15017_/C sky130_fd_sc_hd__or4_4
XFILLER_170_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12219_ _21442_/A VGND VGND VPWR VPWR _12219_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24203__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13199_ _13199_/A VGND VGND VPWR VPWR _13200_/A sky130_fd_sc_hd__buf_2
XFILLER_243_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19815_ _19812_/Y _19806_/X _19813_/X _19814_/X VGND VGND VPWR VPWR _23608_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_243_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17254__A _17234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16958_ _24722_/Q _16957_/Y _16003_/Y _16965_/A VGND VGND VPWR VPWR _16960_/C sky130_fd_sc_hd__a2bb2o_4
X_19746_ HWDATA[5] VGND VGND VPWR VPWR _19746_/X sky130_fd_sc_hd__buf_2
XFILLER_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15909_ _15681_/X _14764_/A _15688_/A _15904_/B VGND VGND VPWR VPWR _15910_/A sky130_fd_sc_hd__a211o_4
XANTENNA__25409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19677_ _13266_/B VGND VGND VPWR VPWR _19677_/Y sky130_fd_sc_hd__inv_2
X_16889_ _22190_/A VGND VGND VPWR VPWR _16889_/Y sky130_fd_sc_hd__inv_2
X_18628_ _24145_/Q VGND VGND VPWR VPWR _18693_/C sky130_fd_sc_hd__inv_2
XFILLER_225_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25062__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18559_ _18559_/A VGND VGND VPWR VPWR _18559_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25467__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19363__B1 _19295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21570_ _21570_/A VGND VGND VPWR VPWR _21570_/X sky130_fd_sc_hd__buf_2
XANTENNA__21223__B _21213_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_37_0_HCLK clkbuf_6_37_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_75_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20521_ _20465_/B _20520_/X _20505_/X VGND VGND VPWR VPWR _20521_/X sky130_fd_sc_hd__o21a_4
XFILLER_192_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23240_ _16550_/A _23171_/X _22839_/X _23239_/X VGND VGND VPWR VPWR _23240_/X sky130_fd_sc_hd__a211o_4
X_20452_ _20464_/C VGND VGND VPWR VPWR _20453_/D sky130_fd_sc_hd__inv_2
XFILLER_134_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23171_ _23171_/A VGND VGND VPWR VPWR _23171_/X sky130_fd_sc_hd__buf_2
XFILLER_106_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20383_ _14084_/Y _23935_/Q VGND VGND VPWR VPWR _20384_/A sky130_fd_sc_hd__or2_4
XFILLER_134_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22122_ _14251_/Y _21721_/B _17420_/Y _21722_/B VGND VGND VPWR VPWR _22122_/X sky130_fd_sc_hd__o22a_4
XANTENNA__15152__B2 _24584_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22053_ _19530_/Y _22001_/Y _22395_/A _22052_/X VGND VGND VPWR VPWR _22053_/X sky130_fd_sc_hd__a211o_4
XFILLER_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21004_ _23972_/Q VGND VGND VPWR VPWR _21006_/A sky130_fd_sc_hd__inv_2
XFILLER_153_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12910__B1 _12862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23997__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23926__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22955_ _14964_/A _22838_/X _22098_/X _22954_/X VGND VGND VPWR VPWR _22956_/C sky130_fd_sc_hd__a211o_4
XFILLER_46_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21906_ _21913_/A _21906_/B VGND VGND VPWR VPWR _21906_/X sky130_fd_sc_hd__or2_4
XFILLER_216_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22886_ _24565_/Q _22885_/X _22802_/X VGND VGND VPWR VPWR _22886_/X sky130_fd_sc_hd__o21a_4
XFILLER_70_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_119_0_HCLK clkbuf_6_59_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_239_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24625_ _24618_/CLK _16328_/X HRESETn VGND VGND VPWR VPWR _24625_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21837_ _14220_/Y _14212_/A _15465_/Y _15457_/A VGND VGND VPWR VPWR _21839_/B sky130_fd_sc_hd__o22a_4
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23332__C _23331_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19354__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12570_ _24883_/Q VGND VGND VPWR VPWR _12570_/Y sky130_fd_sc_hd__inv_2
X_21768_ _22379_/A _19909_/Y VGND VGND VPWR VPWR _21769_/C sky130_fd_sc_hd__or2_4
X_24556_ _24555_/CLK _16514_/X HRESETn VGND VGND VPWR VPWR _16512_/A sky130_fd_sc_hd__dfrtp_4
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20719_ _13117_/A _13117_/B _20718_/Y VGND VGND VPWR VPWR _20719_/Y sky130_fd_sc_hd__a21oi_4
X_23507_ _23525_/CLK _20084_/X VGND VGND VPWR VPWR _20083_/A sky130_fd_sc_hd__dfxtp_4
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24785__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21699_ _16637_/A _21698_/X _21436_/X _25523_/Q _22522_/B VGND VGND VPWR VPWR _21700_/B
+ sky130_fd_sc_hd__a32o_4
X_24487_ _24487_/CLK _16698_/X HRESETn VGND VGND VPWR VPWR _16696_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_169_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240_ _23997_/Q _14236_/X _14239_/X VGND VGND VPWR VPWR _14240_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_109_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23438_ _23437_/CLK _23438_/D VGND VGND VPWR VPWR _23438_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24714__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14171_ _25130_/Q VGND VGND VPWR VPWR _14171_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23369_ _21016_/X VGND VGND VPWR VPWR IRQ[25] sky130_fd_sc_hd__buf_2
X_13122_ _20789_/A _13122_/B _20754_/A VGND VGND VPWR VPWR _13122_/X sky130_fd_sc_hd__or3_4
X_25108_ _25109_/CLK _25108_/D HRESETn VGND VGND VPWR VPWR _25108_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16340__B1 _16145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_57_0_HCLK clkbuf_7_28_0_HCLK/X VGND VGND VPWR VPWR _24233_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13053_ _13041_/B VGND VGND VPWR VPWR _13054_/B sky130_fd_sc_hd__inv_2
X_17930_ _24250_/Q _17917_/Y _17926_/X VGND VGND VPWR VPWR _24250_/D sky130_fd_sc_hd__o21a_4
XFILLER_124_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25039_ _25015_/CLK _25039_/D HRESETn VGND VGND VPWR VPWR _14883_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16891__B2 _24283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22413__B1 _24723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12004_ _12000_/Y _20968_/A _12000_/Y _20968_/A VGND VGND VPWR VPWR _12004_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12901__B1 _12854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17861_ _17860_/X VGND VGND VPWR VPWR _24268_/D sky130_fd_sc_hd__inv_2
XANTENNA__24957__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16812_ _14966_/Y _16808_/X HWDATA[22] _16808_/X VGND VGND VPWR VPWR _16812_/X sky130_fd_sc_hd__a2bb2o_4
X_19600_ _19600_/A VGND VGND VPWR VPWR _19600_/X sky130_fd_sc_hd__buf_2
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17792_ _17764_/X _17773_/X _17743_/Y VGND VGND VPWR VPWR _17792_/X sky130_fd_sc_hd__o21a_4
X_19531_ _19526_/A VGND VGND VPWR VPWR _19531_/X sky130_fd_sc_hd__buf_2
XFILLER_219_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16743_ _16743_/A VGND VGND VPWR VPWR _16743_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25502__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13955_ _13956_/A _13955_/B VGND VGND VPWR VPWR _13955_/X sky130_fd_sc_hd__and2_4
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19593__B1 _19543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12906_ _12889_/X _12906_/B _12905_/Y VGND VGND VPWR VPWR _25386_/D sky130_fd_sc_hd__and3_4
X_19462_ _19462_/A VGND VGND VPWR VPWR _22026_/B sky130_fd_sc_hd__inv_2
X_16674_ _16672_/Y _16668_/X _16400_/X _16673_/X VGND VGND VPWR VPWR _16674_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13886_ _13903_/B VGND VGND VPWR VPWR _13907_/B sky130_fd_sc_hd__buf_2
XANTENNA__15749__A3 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18413_ _24165_/Q VGND VGND VPWR VPWR _18577_/A sky130_fd_sc_hd__inv_2
XFILLER_62_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15625_ _15625_/A VGND VGND VPWR VPWR _15625_/Y sky130_fd_sc_hd__inv_2
X_12837_ _12800_/Y _12837_/B _12836_/Y _12813_/Y VGND VGND VPWR VPWR _12837_/X sky130_fd_sc_hd__or4_4
X_19393_ _19391_/Y _19389_/X _19392_/X _19389_/X VGND VGND VPWR VPWR _23753_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18344_ _17450_/X _18341_/A VGND VGND VPWR VPWR _18344_/X sky130_fd_sc_hd__and2_4
XFILLER_188_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15556_ _15556_/A VGND VGND VPWR VPWR _15556_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12768_ _12766_/A _22901_/A _12766_/Y _12767_/Y VGND VGND VPWR VPWR _12768_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21152__B1 _21574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14507_ _14491_/X _14505_/X _25121_/Q _14506_/X VGND VGND VPWR VPWR _25109_/D sky130_fd_sc_hd__o22a_4
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11719_ _11717_/Y _11714_/X _11718_/X _11714_/X VGND VGND VPWR VPWR _25538_/D sky130_fd_sc_hd__a2bb2o_4
X_18275_ _13772_/D _18240_/A _13459_/A _13682_/A _18274_/X VGND VGND VPWR VPWR _24220_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_175_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15487_ _11651_/Y _15486_/X HWRITE _15486_/X VGND VGND VPWR VPWR _24949_/D sky130_fd_sc_hd__a2bb2o_4
X_12699_ _12498_/Y _12701_/B _12698_/Y VGND VGND VPWR VPWR _25412_/D sky130_fd_sc_hd__o21a_4
XFILLER_147_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17226_ _17226_/A _17223_/X _17224_/X _17226_/D VGND VGND VPWR VPWR _17227_/D sky130_fd_sc_hd__or4_4
X_14438_ _14158_/Y _14437_/X _14384_/X _14437_/X VGND VGND VPWR VPWR _14438_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24455__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17157_ _17153_/B _17157_/B _17148_/C VGND VGND VPWR VPWR _17157_/X sky130_fd_sc_hd__and3_4
XFILLER_116_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14369_ _13965_/X _14369_/B VGND VGND VPWR VPWR _14369_/X sky130_fd_sc_hd__or2_4
XANTENNA__12681__A _12681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16108_ _24703_/Q VGND VGND VPWR VPWR _16108_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17088_ _17020_/Y _17088_/B VGND VGND VPWR VPWR _17097_/B sky130_fd_sc_hd__or2_4
XFILLER_170_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16039_ _16037_/Y _16033_/X _11735_/X _16038_/X VGND VGND VPWR VPWR _16039_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19729_ _19727_/Y _19723_/X _19728_/X _19723_/X VGND VGND VPWR VPWR _23638_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19584__B1 _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22740_ _22740_/A VGND VGND VPWR VPWR _22740_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21391__B1 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22671_ _15014_/Y _21047_/X VGND VGND VPWR VPWR _22671_/X sky130_fd_sc_hd__and2_4
XFILLER_41_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11760__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21622_ _21622_/A VGND VGND VPWR VPWR _22381_/A sky130_fd_sc_hd__buf_2
X_24410_ _23808_/CLK _24410_/D HRESETn VGND VGND VPWR VPWR _20099_/A sky130_fd_sc_hd__dfrtp_4
X_25390_ _25390_/CLK _25390_/D HRESETn VGND VGND VPWR VPWR _25390_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21143__B1 _21343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21553_ _14382_/Y _14183_/X _14454_/Y _17412_/X VGND VGND VPWR VPWR _21553_/X sky130_fd_sc_hd__o22a_4
X_24341_ _24341_/CLK _24341_/D HRESETn VGND VGND VPWR VPWR _17239_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_139_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20504_ _20504_/A _20503_/X VGND VGND VPWR VPWR _24081_/D sky130_fd_sc_hd__or2_4
XANTENNA__24076__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24272_ _24278_/CLK _24272_/D HRESETn VGND VGND VPWR VPWR _24272_/Q sky130_fd_sc_hd__dfrtp_4
X_21484_ _21462_/A VGND VGND VPWR VPWR _21484_/X sky130_fd_sc_hd__buf_2
XANTENNA__24196__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16570__B1 _16395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23223_ _23044_/X _23222_/X _23046_/X _24744_/Q _23152_/X VGND VGND VPWR VPWR _23223_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_165_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20435_ _20437_/A _20435_/B VGND VGND VPWR VPWR _20435_/X sky130_fd_sc_hd__and2_4
XANTENNA__17495__A1_N _25526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12591__A _12680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24125__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_210_0_HCLK clkbuf_8_211_0_HCLK/A VGND VGND VPWR VPWR _24487_/CLK sky130_fd_sc_hd__clkbuf_1
X_23154_ _23153_/X VGND VGND VPWR VPWR _23154_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20366_ _23402_/Q VGND VGND VPWR VPWR _21179_/B sky130_fd_sc_hd__inv_2
X_22105_ _23924_/Q VGND VGND VPWR VPWR _22105_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23085_ _16657_/Y _22829_/X _15572_/Y _22832_/X VGND VGND VPWR VPWR _23085_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20297_ _20297_/A VGND VGND VPWR VPWR _21807_/B sky130_fd_sc_hd__inv_2
XFILLER_121_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22036_ _21670_/X _19883_/Y _21674_/X VGND VGND VPWR VPWR _22036_/X sky130_fd_sc_hd__o21a_4
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21409__A _22202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17822__B1 _16952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23987_ _25050_/CLK _20670_/Y HRESETn VGND VGND VPWR VPWR _17396_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13740_ _13739_/Y VGND VGND VPWR VPWR _13741_/D sky130_fd_sc_hd__buf_2
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20951__A1_N _20828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22938_ _22913_/X _22920_/X _22924_/Y _22937_/X VGND VGND VPWR VPWR HRDATA[19] sky130_fd_sc_hd__a211o_4
XFILLER_44_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13671_ _11803_/Y _13670_/X VGND VGND VPWR VPWR _13672_/B sky130_fd_sc_hd__or2_4
XFILLER_44_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22869_ _22145_/B VGND VGND VPWR VPWR _22909_/B sky130_fd_sc_hd__buf_2
XANTENNA__12766__A _12766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24966__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15410_ _15296_/B _15418_/A VGND VGND VPWR VPWR _15410_/X sky130_fd_sc_hd__or2_4
XFILLER_232_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15142__A _24600_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12622_ _12624_/B VGND VGND VPWR VPWR _12623_/B sky130_fd_sc_hd__inv_2
X_24608_ _24591_/CLK _16378_/X HRESETn VGND VGND VPWR VPWR _23242_/A sky130_fd_sc_hd__dfrtp_4
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16390_ _16389_/Y _16387_/X _16301_/X _16387_/X VGND VGND VPWR VPWR _16390_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16074__A1_N _16073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15341_ _15338_/A _15333_/B _15341_/C VGND VGND VPWR VPWR _15341_/X sky130_fd_sc_hd__and3_4
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12553_ _12553_/A VGND VGND VPWR VPWR _12553_/Y sky130_fd_sc_hd__inv_2
X_24539_ _24539_/CLK _16561_/X HRESETn VGND VGND VPWR VPWR _24539_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19549__A _19548_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18060_ _18060_/A _18060_/B _18059_/X VGND VGND VPWR VPWR _18060_/X sky130_fd_sc_hd__and3_4
Xclkbuf_6_20_0_HCLK clkbuf_5_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15272_ _15272_/A _15243_/B VGND VGND VPWR VPWR _15273_/B sky130_fd_sc_hd__or2_4
XFILLER_8_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ _12266_/C _12458_/B _12398_/X _12482_/B VGND VGND VPWR VPWR _12484_/X sky130_fd_sc_hd__a211o_4
XANTENNA__16561__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17011_ _24744_/Q _17022_/A _16064_/Y _17039_/A VGND VGND VPWR VPWR _17011_/X sky130_fd_sc_hd__a2bb2o_4
X_14223_ _14222_/Y _14218_/X _13788_/X _14218_/X VGND VGND VPWR VPWR _14223_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22406__C _22296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22634__B1 _24832_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14154_ _14154_/A _14162_/A _14160_/A _14111_/X VGND VGND VPWR VPWR _14154_/X sky130_fd_sc_hd__or4_4
XFILLER_125_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13105_ _13105_/A VGND VGND VPWR VPWR _13105_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14085_ scl_oen_o_S4 _14084_/Y _23935_/Q VGND VGND VPWR VPWR _14096_/B sky130_fd_sc_hd__and3_4
X_18962_ _18078_/B VGND VGND VPWR VPWR _18962_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13036_ _12975_/Y _13033_/X VGND VGND VPWR VPWR _13036_/X sky130_fd_sc_hd__or2_4
X_17913_ _17912_/Y _17908_/Y _21993_/A _17908_/A VGND VGND VPWR VPWR _24254_/D sky130_fd_sc_hd__o22a_4
XANTENNA__11689__B1 _11688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21319__A _21111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18893_ _18871_/X _18885_/X _20982_/B _24120_/Q _18888_/X VGND VGND VPWR VPWR _24120_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12350__B2 _12293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17844_ _17755_/Y _17842_/A VGND VGND VPWR VPWR _17845_/C sky130_fd_sc_hd__or2_4
XFILLER_67_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18653__A2_N _18769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17775_ _16913_/Y _16945_/X _17775_/C VGND VGND VPWR VPWR _17775_/X sky130_fd_sc_hd__or3_4
X_14987_ _15272_/A _16786_/A _25013_/Q _14986_/Y VGND VGND VPWR VPWR _14987_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22165__A2 _21325_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16726_ _16726_/A VGND VGND VPWR VPWR _16726_/X sky130_fd_sc_hd__buf_2
X_19514_ _23709_/Q VGND VGND VPWR VPWR _21681_/B sky130_fd_sc_hd__inv_2
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13938_ _13927_/A _13938_/B _13913_/X _13937_/Y VGND VGND VPWR VPWR _13938_/X sky130_fd_sc_hd__and4_4
XFILLER_47_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23253__B _22817_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20176__B2 _20158_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14875__B _14817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19445_ _19444_/Y _19440_/X _19377_/X _19440_/X VGND VGND VPWR VPWR _23734_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21054__A _11664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16657_ _24503_/Q VGND VGND VPWR VPWR _16657_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13869_ _25245_/Q _13849_/X _25244_/Q _13844_/X VGND VGND VPWR VPWR _13869_/X sky130_fd_sc_hd__o22a_4
XFILLER_222_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19318__B1 _19295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_102_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_205_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15608_ _15608_/A VGND VGND VPWR VPWR _15608_/X sky130_fd_sc_hd__buf_2
XFILLER_223_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19376_ _19376_/A VGND VGND VPWR VPWR _19376_/Y sky130_fd_sc_hd__inv_2
X_16588_ _16587_/Y _16585_/X _16233_/X _16585_/X VGND VGND VPWR VPWR _24528_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24636__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18327_ _20054_/B VGND VGND VPWR VPWR _18328_/A sky130_fd_sc_hd__buf_2
XFILLER_188_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15539_ _11706_/X VGND VGND VPWR VPWR _15724_/A sky130_fd_sc_hd__buf_2
XFILLER_203_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18258_ _13807_/D _18256_/X _18257_/X _24229_/Q _18241_/A VGND VGND VPWR VPWR _24229_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_163_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17209_ _16327_/Y _17336_/A _16327_/Y _17336_/A VGND VGND VPWR VPWR _17213_/A sky130_fd_sc_hd__a2bb2o_4
X_18189_ _18125_/A _23844_/Q VGND VGND VPWR VPWR _18191_/B sky130_fd_sc_hd__or2_4
XFILLER_162_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20220_ _20220_/A _20220_/B _20387_/A _20220_/D VGND VGND VPWR VPWR _20220_/X sky130_fd_sc_hd__or4_4
XANTENNA__13300__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16304__B1 _15942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20151_ _21623_/B _20150_/X _20106_/X _20150_/X VGND VGND VPWR VPWR _20151_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25495__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_40_0_HCLK clkbuf_7_20_0_HCLK/X VGND VGND VPWR VPWR _24679_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__25424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20082_ _21412_/B _20079_/X _19827_/X _20079_/X VGND VGND VPWR VPWR _23508_/D sky130_fd_sc_hd__a2bb2o_4
X_23910_ _23452_/CLK _23910_/D VGND VGND VPWR VPWR _18944_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21600__A1 _21119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12341__B2 _24833_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24890_ _24907_/CLK _15672_/X HRESETn VGND VGND VPWR VPWR _13658_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_245_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23841_ _23831_/CLK _23841_/D VGND VGND VPWR VPWR _23841_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20984_ _20984_/A _20984_/B VGND VGND VPWR VPWR _20984_/X sky130_fd_sc_hd__and2_4
X_23772_ _23889_/CLK _19337_/X VGND VGND VPWR VPWR _23772_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25511_ _24679_/CLK _11893_/X HRESETn VGND VGND VPWR VPWR _11848_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_225_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22723_ _22723_/A VGND VGND VPWR VPWR _22723_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16058__A _16038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19309__B1 _19194_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25442_ _25444_/CLK _12472_/X HRESETn VGND VGND VPWR VPWR _12207_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22654_ _24761_/Q _22654_/B VGND VGND VPWR VPWR _22654_/X sky130_fd_sc_hd__or2_4
XFILLER_230_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24377__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21605_ _21775_/A _21605_/B VGND VGND VPWR VPWR _21605_/X sky130_fd_sc_hd__or2_4
XFILLER_185_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22585_ _22515_/X _22583_/X _21956_/X _22584_/X VGND VGND VPWR VPWR _22585_/X sky130_fd_sc_hd__o22a_4
X_25373_ _25373_/CLK _25373_/D HRESETn VGND VGND VPWR VPWR _25373_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24306__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24324_ _25081_/CLK _24324_/D HRESETn VGND VGND VPWR VPWR _24324_/Q sky130_fd_sc_hd__dfstp_4
X_21536_ _21535_/X VGND VGND VPWR VPWR _21536_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16543__B1 _15545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21467_ _21662_/A _21467_/B VGND VGND VPWR VPWR _21467_/X sky130_fd_sc_hd__or2_4
X_24255_ _24257_/CLK _24255_/D HRESETn VGND VGND VPWR VPWR _21991_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13210__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20418_ _21897_/B _20415_/X _16867_/X _20415_/X VGND VGND VPWR VPWR _23381_/D sky130_fd_sc_hd__a2bb2o_4
X_23206_ _23206_/A _23063_/X VGND VGND VPWR VPWR _23206_/X sky130_fd_sc_hd__or2_4
XFILLER_135_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21398_ _14681_/A _21396_/X _21397_/X VGND VGND VPWR VPWR _21398_/X sky130_fd_sc_hd__and3_4
X_24186_ _24159_/CLK _24186_/D HRESETn VGND VGND VPWR VPWR _24186_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22631__A3 _22296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20349_ _20348_/X VGND VGND VPWR VPWR _20349_/Y sky130_fd_sc_hd__inv_2
X_23137_ _24605_/Q _23177_/B VGND VGND VPWR VPWR _23141_/B sky130_fd_sc_hd__or2_4
XFILLER_134_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23941__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23068_ _24603_/Q _23177_/B VGND VGND VPWR VPWR _23071_/B sky130_fd_sc_hd__or2_4
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14910_ _25016_/Q VGND VGND VPWR VPWR _15002_/A sky130_fd_sc_hd__inv_2
X_22019_ _22014_/A _20333_/Y VGND VGND VPWR VPWR _22019_/X sky130_fd_sc_hd__or2_4
XFILLER_248_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15890_ _12743_/Y _15889_/X _13818_/X _15889_/X VGND VGND VPWR VPWR _15890_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14841_ _14811_/A _14811_/B _14811_/A _14811_/B VGND VGND VPWR VPWR _14842_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17560_ _17559_/Y VGND VGND VPWR VPWR _17614_/A sky130_fd_sc_hd__buf_2
XANTENNA__12096__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17352__A _17358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14772_ _25059_/Q _14769_/B _14758_/A _14758_/B VGND VGND VPWR VPWR _14772_/X sky130_fd_sc_hd__a211o_4
XFILLER_91_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11984_ _11977_/X VGND VGND VPWR VPWR _11984_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12635__A2 _12626_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16511_ _16510_/Y _16508_/X _16420_/X _16508_/X VGND VGND VPWR VPWR _16511_/X sky130_fd_sc_hd__a2bb2o_4
X_13723_ _13723_/A VGND VGND VPWR VPWR _19072_/C sky130_fd_sc_hd__buf_2
X_17491_ _17491_/A VGND VGND VPWR VPWR _17590_/A sky130_fd_sc_hd__inv_2
XANTENNA__12496__A _21078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19230_ _19230_/A VGND VGND VPWR VPWR _22365_/B sky130_fd_sc_hd__inv_2
XFILLER_232_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16442_ _16180_/A VGND VGND VPWR VPWR _22995_/A sky130_fd_sc_hd__inv_2
X_13654_ _20953_/A _20953_/B _24065_/Q _13653_/X VGND VGND VPWR VPWR _13655_/B sky130_fd_sc_hd__or4_4
XFILLER_231_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12605_ _12600_/X _12605_/B _12605_/C VGND VGND VPWR VPWR _12681_/B sky130_fd_sc_hd__or3_4
X_19161_ _19160_/Y _19156_/X _19138_/X _19149_/A VGND VGND VPWR VPWR _23835_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21602__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16373_ HWDATA[30] VGND VGND VPWR VPWR _16373_/X sky130_fd_sc_hd__buf_2
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19279__A _18981_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24047__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13585_ _14364_/A _21283_/A _25057_/Q _13584_/X VGND VGND VPWR VPWR _13586_/A sky130_fd_sc_hd__or4_4
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18112_ _14636_/A _18110_/X _18111_/X VGND VGND VPWR VPWR _18112_/X sky130_fd_sc_hd__and3_4
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22417__B _22417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15324_ _15324_/A VGND VGND VPWR VPWR _15324_/Y sky130_fd_sc_hd__inv_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12536_ _25410_/Q VGND VGND VPWR VPWR _12696_/A sky130_fd_sc_hd__inv_2
X_19092_ _21250_/B _19086_/X _19091_/X _19074_/A VGND VGND VPWR VPWR _23859_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18043_ _17947_/A _18043_/B _18042_/X VGND VGND VPWR VPWR _18043_/X sky130_fd_sc_hd__and3_4
XFILLER_184_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15888__A2 _15887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15255_ _15254_/X VGND VGND VPWR VPWR _15256_/B sky130_fd_sc_hd__inv_2
XFILLER_145_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12467_ _12466_/X VGND VGND VPWR VPWR _12467_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14206_ _14205_/Y _14190_/A _13788_/X _14190_/A VGND VGND VPWR VPWR _14206_/X sky130_fd_sc_hd__a2bb2o_4
X_15186_ _15185_/X VGND VGND VPWR VPWR _25034_/D sky130_fd_sc_hd__inv_2
X_12398_ _12415_/A VGND VGND VPWR VPWR _12398_/X sky130_fd_sc_hd__buf_2
XFILLER_126_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14137_ _14137_/A VGND VGND VPWR VPWR _14137_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19994_ _19993_/Y _19991_/X _19967_/X _19991_/X VGND VGND VPWR VPWR _19994_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_152_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16581__A1_N _16578_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_27_0_HCLK clkbuf_7_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24070__D _24070_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14068_ _13979_/C _14054_/X _14067_/X _13987_/X _14065_/X VGND VGND VPWR VPWR _14068_/X
+ sky130_fd_sc_hd__a32o_4
X_18945_ _18944_/Y _18939_/X _16783_/X _18939_/X VGND VGND VPWR VPWR _23910_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19787__B1 _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13019_ _13028_/A VGND VGND VPWR VPWR _13019_/X sky130_fd_sc_hd__buf_2
X_18876_ _18876_/A _18875_/X VGND VGND VPWR VPWR _18876_/X sky130_fd_sc_hd__or2_4
XFILLER_121_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21594__B1 _22290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17827_ _17818_/A _17827_/B _17826_/Y VGND VGND VPWR VPWR _24276_/D sky130_fd_sc_hd__and3_4
XANTENNA__24888__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23335__A1 _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15812__A2 _15789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17262__A _17261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17758_ _24272_/Q VGND VGND VPWR VPWR _17758_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24817__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16709_ _16692_/A VGND VGND VPWR VPWR _16709_/X sky130_fd_sc_hd__buf_2
X_17689_ _17578_/Y _17666_/B _17687_/B _17604_/X VGND VGND VPWR VPWR _17690_/A sky130_fd_sc_hd__a211o_4
X_19428_ _18175_/B VGND VGND VPWR VPWR _19428_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16773__B1 _16518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24470__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21512__A _18900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19359_ _23764_/Q VGND VGND VPWR VPWR _19359_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22310__A2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22327__B _22327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22370_ _22366_/X _22369_/X _21773_/X VGND VGND VPWR VPWR _22370_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_175_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20128__A _20116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21321_ _21289_/X _21301_/X _21306_/X _21314_/X _21320_/X VGND VGND VPWR VPWR _21321_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_163_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21252_ _21252_/A VGND VGND VPWR VPWR _22223_/A sky130_fd_sc_hd__buf_2
X_24040_ _24486_/CLK _24040_/D HRESETn VGND VGND VPWR VPWR _13644_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_117_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20203_ _17980_/B VGND VGND VPWR VPWR _20203_/Y sky130_fd_sc_hd__inv_2
X_21183_ _24212_/Q VGND VGND VPWR VPWR _21205_/A sky130_fd_sc_hd__buf_2
XANTENNA__16341__A _24619_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20134_ _21269_/B _20128_/X _20133_/X _20116_/A VGND VGND VPWR VPWR _20134_/X sky130_fd_sc_hd__a2bb2o_4
X_20065_ _23514_/Q VGND VGND VPWR VPWR _20065_/Y sky130_fd_sc_hd__inv_2
X_24942_ _25510_/CLK _15500_/X HRESETn VGND VGND VPWR VPWR _24942_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_219_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19652__A _19006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21585__B1 _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24873_ _25409_/CLK _15733_/X HRESETn VGND VGND VPWR VPWR _24873_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_245_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23824_ _23831_/CLK _19192_/X VGND VGND VPWR VPWR _19190_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24558__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ _23774_/CLK _19385_/X VGND VGND VPWR VPWR _18200_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _11983_/B _13506_/A VGND VGND VPWR VPWR _24095_/D sky130_fd_sc_hd__and2_4
XPHY_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18753__A1 _18658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22706_ _24561_/Q _21843_/B _21864_/C VGND VGND VPWR VPWR _22706_/X sky130_fd_sc_hd__and3_4
XFILLER_198_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13205__A _13289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23686_ _24208_/CLK _23686_/D VGND VGND VPWR VPWR _23686_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_110_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16764__B1 _15746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _24051_/Q VGND VGND VPWR VPWR _20898_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25425_ _24872_/CLK _25425_/D HRESETn VGND VGND VPWR VPWR _12526_/A sky130_fd_sc_hd__dfrtp_4
X_22637_ _21077_/A _22634_/X _21114_/X _22636_/X VGND VGND VPWR VPWR _22637_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__24140__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13370_ _13434_/A _13370_/B _13370_/C VGND VGND VPWR VPWR _13370_/X sky130_fd_sc_hd__and3_4
X_25356_ _25346_/CLK _25356_/D HRESETn VGND VGND VPWR VPWR _25356_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16516__B1 _16145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22568_ _21121_/A _22566_/X _22111_/X _22567_/X VGND VGND VPWR VPWR _22569_/B sky130_fd_sc_hd__o22a_4
XFILLER_221_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12321_ _12321_/A VGND VGND VPWR VPWR _12321_/Y sky130_fd_sc_hd__inv_2
X_24307_ _25533_/CLK _17649_/X HRESETn VGND VGND VPWR VPWR _24307_/Q sky130_fd_sc_hd__dfrtp_4
X_21519_ _21519_/A VGND VGND VPWR VPWR _21843_/B sky130_fd_sc_hd__buf_2
X_25287_ _25292_/CLK _25287_/D HRESETn VGND VGND VPWR VPWR _11810_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_108_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22499_ _21531_/X VGND VGND VPWR VPWR _22499_/X sky130_fd_sc_hd__buf_2
XFILLER_6_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15040_ _15039_/X _24460_/Q _15039_/X _24460_/Q VGND VGND VPWR VPWR _15040_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18269__B1 _16849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12252_ _12269_/A VGND VGND VPWR VPWR _12252_/X sky130_fd_sc_hd__buf_2
X_24238_ _24341_/CLK _18244_/X HRESETn VGND VGND VPWR VPWR _22620_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_170_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25346__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12183_ _25454_/Q _12181_/Y _12170_/A _12182_/Y VGND VGND VPWR VPWR _12186_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17347__A _17358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24169_ _24325_/CLK _24169_/D HRESETn VGND VGND VPWR VPWR _18473_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16991_ _16991_/A VGND VGND VPWR VPWR _16991_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17492__B2 _24114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15942_ HWDATA[22] VGND VGND VPWR VPWR _15942_/X sky130_fd_sc_hd__buf_2
X_18730_ _18730_/A _18730_/B VGND VGND VPWR VPWR _18733_/B sky130_fd_sc_hd__or2_4
XFILLER_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18661_ _16564_/A _18728_/A _16569_/Y _24146_/Q VGND VGND VPWR VPWR _18661_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_236_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15873_ _12746_/Y _15872_/X _15581_/X _15872_/X VGND VGND VPWR VPWR _15873_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24981__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23317__A1 _22552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23317__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14824_ _14826_/A _14822_/X _14215_/Y _14823_/X VGND VGND VPWR VPWR _14824_/X sky130_fd_sc_hd__o22a_4
X_17612_ _17625_/A _17607_/Y _17612_/C VGND VGND VPWR VPWR _17613_/A sky130_fd_sc_hd__or3_4
X_18592_ _18420_/Y _18592_/B VGND VGND VPWR VPWR _18592_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24299__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24910__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17543_ _17543_/A VGND VGND VPWR VPWR _17543_/Y sky130_fd_sc_hd__inv_2
X_14755_ _14755_/A VGND VGND VPWR VPWR _14756_/A sky130_fd_sc_hd__buf_2
XANTENNA__24228__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11967_ _11967_/A _11932_/B _11962_/X VGND VGND VPWR VPWR _11967_/X sky130_fd_sc_hd__and3_4
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13706_ _13675_/B _13694_/X _13705_/Y _13701_/X _11814_/A VGND VGND VPWR VPWR _25288_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_205_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17474_ _17473_/Y _17448_/A VGND VGND VPWR VPWR _17480_/A sky130_fd_sc_hd__or2_4
X_14686_ _21252_/A VGND VGND VPWR VPWR _22196_/A sky130_fd_sc_hd__inv_2
X_11898_ _11897_/X VGND VGND VPWR VPWR _11898_/X sky130_fd_sc_hd__buf_2
X_16425_ _15100_/Y _16422_/X _16055_/X _16422_/X VGND VGND VPWR VPWR _16425_/X sky130_fd_sc_hd__a2bb2o_4
X_19213_ _23817_/Q VGND VGND VPWR VPWR _19213_/Y sky130_fd_sc_hd__inv_2
X_13637_ _24056_/Q _24055_/Q _24057_/Q _13637_/D VGND VGND VPWR VPWR _13637_/X sky130_fd_sc_hd__or4_4
XFILLER_220_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23096__A3 _22849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19144_ _19006_/A VGND VGND VPWR VPWR _19144_/X sky130_fd_sc_hd__buf_2
X_16356_ _16355_/Y _16350_/X _15976_/X _16350_/X VGND VGND VPWR VPWR _16356_/X sky130_fd_sc_hd__a2bb2o_4
X_13568_ _13820_/A _14557_/A _22540_/A _25093_/Q VGND VGND VPWR VPWR _13568_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_185_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15307_ _15070_/A _15307_/B VGND VGND VPWR VPWR _15307_/X sky130_fd_sc_hd__or2_4
XFILLER_158_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12519_ _12519_/A _12513_/X _12516_/X _12519_/D VGND VGND VPWR VPWR _12519_/X sky130_fd_sc_hd__or4_4
X_19075_ _19071_/Y _19074_/X _16860_/X _19074_/X VGND VGND VPWR VPWR _23866_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16287_ _24640_/Q VGND VGND VPWR VPWR _16287_/Y sky130_fd_sc_hd__inv_2
X_13499_ _13499_/A VGND VGND VPWR VPWR _13499_/X sky130_fd_sc_hd__buf_2
XFILLER_246_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18026_ _18026_/A VGND VGND VPWR VPWR _18030_/A sky130_fd_sc_hd__buf_2
XFILLER_8_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15238_ _15203_/X _15236_/X _15237_/X VGND VGND VPWR VPWR _25021_/D sky130_fd_sc_hd__and3_4
XANTENNA__25087__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17257__A _17333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13785__A _14380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25016__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15169_ _14982_/A VGND VGND VPWR VPWR _15169_/X sky130_fd_sc_hd__buf_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18275__A3 _13459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16161__A _21435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19977_ _19977_/A VGND VGND VPWR VPWR _19977_/X sky130_fd_sc_hd__buf_2
XANTENNA__14297__A1 MSO_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18928_ _18927_/Y _18925_/X _16787_/X _18925_/X VGND VGND VPWR VPWR _18928_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_28_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18859_ _16500_/Y _24140_/Q _16500_/Y _24140_/Q VGND VGND VPWR VPWR _18859_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_114_0_HCLK clkbuf_7_57_0_HCLK/X VGND VGND VPWR VPWR _24800_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23308__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23308__B2 _22838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_177_0_HCLK clkbuf_7_88_0_HCLK/X VGND VGND VPWR VPWR _25140_/CLK sky130_fd_sc_hd__clkbuf_1
X_21870_ _21745_/B VGND VGND VPWR VPWR _23171_/A sky130_fd_sc_hd__buf_2
XFILLER_131_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24651__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16994__B1 _16037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20821_ _20684_/A _13126_/A _13125_/X _23324_/A _20735_/X VGND VGND VPWR VPWR _24034_/D
+ sky130_fd_sc_hd__a32o_4
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23540_ _23411_/CLK _20006_/X VGND VGND VPWR VPWR _23540_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_211_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20752_ _20731_/X _20751_/X _24907_/Q _20736_/X VGND VGND VPWR VPWR _24017_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_211_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16746__B1 _16483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21242__A _22196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18535__B _18467_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20683_ _20613_/B _20514_/B VGND VGND VPWR VPWR _23998_/D sky130_fd_sc_hd__and2_4
X_23471_ _23487_/CLK _20188_/X VGND VGND VPWR VPWR _23471_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25210_ _23932_/CLK _25210_/D HRESETn VGND VGND VPWR VPWR _14160_/A sky130_fd_sc_hd__dfrtp_4
X_22422_ _22298_/A _22422_/B VGND VGND VPWR VPWR _22422_/X sky130_fd_sc_hd__and2_4
XFILLER_148_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25141_ _23958_/CLK _14413_/X HRESETn VGND VGND VPWR VPWR _25141_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_148_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22353_ _21935_/A _22353_/B VGND VGND VPWR VPWR _22353_/X sky130_fd_sc_hd__or2_4
XFILLER_148_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21304_ _21124_/B VGND VGND VPWR VPWR _21305_/B sky130_fd_sc_hd__buf_2
XFILLER_108_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22284_ _21077_/X _22277_/X _22946_/A _22283_/X VGND VGND VPWR VPWR _22284_/Y sky130_fd_sc_hd__a22oi_4
X_25072_ _23735_/CLK _25072_/D HRESETn VGND VGND VPWR VPWR _19116_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_191_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21235_ _21235_/A _21235_/B _21235_/C VGND VGND VPWR VPWR _21235_/X sky130_fd_sc_hd__and3_4
X_24023_ _24501_/CLK _24023_/D HRESETn VGND VGND VPWR VPWR _13108_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_151_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16071__A _24717_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21166_ _18560_/A _15845_/A _21327_/B VGND VGND VPWR VPWR _21166_/X sky130_fd_sc_hd__and3_4
XFILLER_132_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20117_ _20113_/Y _20116_/X _20089_/X _20116_/X VGND VGND VPWR VPWR _23498_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_219_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_10_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21097_ _24820_/Q _21082_/X _21034_/X _21096_/X VGND VGND VPWR VPWR _21097_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24739__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_73_0_HCLK clkbuf_7_73_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_73_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20048_ _23524_/Q VGND VGND VPWR VPWR _20048_/Y sky130_fd_sc_hd__inv_2
X_24925_ _23378_/CLK _24925_/D HRESETn VGND VGND VPWR VPWR _13581_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__20230__B1 _15762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12870_ _12887_/A VGND VGND VPWR VPWR _12872_/A sky130_fd_sc_hd__buf_2
X_24856_ _24866_/CLK _15767_/X HRESETn VGND VGND VPWR VPWR _12550_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24392__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23973__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11820_/Y _22696_/A _11820_/Y _22696_/A VGND VGND VPWR VPWR _11822_/D sky130_fd_sc_hd__a2bb2o_4
X_23807_ _23808_/CLK _23807_/D VGND VGND VPWR VPWR _23807_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13799__B1 _13798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24321__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ _25375_/CLK _24787_/D HRESETn VGND VGND VPWR VPWR _24787_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21999_ _13772_/D _23346_/B VGND VGND VPWR VPWR _21999_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__14460__B2 _14455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23989__D scl_i_S5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ HSEL VGND VGND VPWR VPWR _14540_/X sky130_fd_sc_hd__buf_2
XFILLER_199_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _25529_/Q VGND VGND VPWR VPWR _11752_/Y sky130_fd_sc_hd__inv_2
X_23738_ _23785_/CLK _23738_/D VGND VGND VPWR VPWR _17958_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _21846_/A _14468_/X _14380_/X _14468_/X VGND VGND VPWR VPWR _25118_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11682_/Y VGND VGND VPWR VPWR _11683_/X sky130_fd_sc_hd__buf_2
X_23669_ _25326_/CLK _19642_/X VGND VGND VPWR VPWR _13375_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16190_/X VGND VGND VPWR VPWR _16210_/X sky130_fd_sc_hd__buf_2
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _13422_/A _13422_/B _13422_/C VGND VGND VPWR VPWR _13426_/B sky130_fd_sc_hd__and3_4
X_25408_ _25403_/CLK _25408_/D HRESETn VGND VGND VPWR VPWR _25408_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17190_ _24631_/Q _24360_/Q _16310_/Y _17251_/C VGND VGND VPWR VPWR _17190_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25527__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12774__A1 _12772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16141_ HWDATA[9] VGND VGND VPWR VPWR _16141_/X sky130_fd_sc_hd__buf_2
X_13353_ _13353_/A _13345_/X _13352_/X VGND VGND VPWR VPWR _13353_/X sky130_fd_sc_hd__and3_4
X_25339_ _25341_/CLK _25339_/D HRESETn VGND VGND VPWR VPWR _12351_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12304_ _25354_/Q _24839_/Q _12302_/Y _12303_/Y VGND VGND VPWR VPWR _12304_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16072_ _16071_/Y _15990_/A _15901_/X _15990_/A VGND VGND VPWR VPWR _16072_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13284_ _13284_/A VGND VGND VPWR VPWR _13434_/A sky130_fd_sc_hd__buf_2
XFILLER_182_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15023_ _24452_/Q VGND VGND VPWR VPWR _15023_/Y sky130_fd_sc_hd__inv_2
X_19900_ _19900_/A VGND VGND VPWR VPWR _19900_/X sky130_fd_sc_hd__buf_2
X_12235_ _12428_/B _24765_/Q _25454_/Q _12181_/Y VGND VGND VPWR VPWR _12239_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21797__B1 _17725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19831_ _23602_/Q VGND VGND VPWR VPWR _19831_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20064__A3 _13459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12166_ _12266_/A _22597_/A _12266_/A _22597_/A VGND VGND VPWR VPWR _12166_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15476__B1 _15475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19762_ _13723_/A _20157_/D _13743_/X _14683_/X VGND VGND VPWR VPWR _19763_/A sky130_fd_sc_hd__or4_4
XANTENNA__17805__A _17744_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12097_ _12097_/A VGND VGND VPWR VPWR _12097_/Y sky130_fd_sc_hd__inv_2
X_16974_ _24740_/Q _24397_/Q _16011_/Y _16973_/Y VGND VGND VPWR VPWR _16977_/C sky130_fd_sc_hd__o22a_4
XFILLER_111_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25139__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18713_ _18713_/A VGND VGND VPWR VPWR _18714_/B sky130_fd_sc_hd__inv_2
X_15925_ _15924_/X VGND VGND VPWR VPWR _15925_/X sky130_fd_sc_hd__buf_2
XFILLER_83_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19693_ _19693_/A VGND VGND VPWR VPWR _19694_/A sky130_fd_sc_hd__inv_2
XANTENNA__24409__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15856_ _15881_/A VGND VGND VPWR VPWR _15857_/A sky130_fd_sc_hd__buf_2
X_18644_ _24516_/Q _18815_/A _24520_/Q _18804_/A VGND VGND VPWR VPWR _18647_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14807_ _14798_/C VGND VGND VPWR VPWR _14814_/A sky130_fd_sc_hd__inv_2
XFILLER_52_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24062__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15787_ _15786_/X VGND VGND VPWR VPWR _15787_/X sky130_fd_sc_hd__buf_2
X_18575_ _18409_/Y _18566_/B VGND VGND VPWR VPWR _18575_/Y sky130_fd_sc_hd__nand2_4
X_12999_ _12999_/A VGND VGND VPWR VPWR _12999_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22513__A2 _22511_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14738_ _14737_/Y _14718_/Y _22044_/A _14718_/A VGND VGND VPWR VPWR _25065_/D sky130_fd_sc_hd__o22a_4
X_17526_ _17497_/X _17506_/X _17526_/C _17526_/D VGND VGND VPWR VPWR _17555_/A sky130_fd_sc_hd__or4_4
XFILLER_233_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16728__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22158__A _22041_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21062__A _22525_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17457_ _19208_/B VGND VGND VPWR VPWR _18326_/C sky130_fd_sc_hd__buf_2
XFILLER_32_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14669_ _14668_/X VGND VGND VPWR VPWR _21622_/A sky130_fd_sc_hd__buf_2
X_16408_ _24595_/Q VGND VGND VPWR VPWR _16408_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17388_ _17388_/A _17388_/B VGND VGND VPWR VPWR _17389_/B sky130_fd_sc_hd__or2_4
XFILLER_119_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22277__B2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16339_ _24620_/Q VGND VGND VPWR VPWR _16339_/Y sky130_fd_sc_hd__inv_2
X_19127_ _19124_/Y _19119_/X _19125_/X _19126_/X VGND VGND VPWR VPWR _19127_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15995__A _24745_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19058_ _19056_/Y _19054_/X _19057_/X _19054_/X VGND VGND VPWR VPWR _23871_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18009_ _18009_/A _18009_/B _18009_/C VGND VGND VPWR VPWR _18021_/B sky130_fd_sc_hd__or3_4
XANTENNA__18248__A3 _16597_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21020_ _21019_/X VGND VGND VPWR VPWR _21021_/A sky130_fd_sc_hd__inv_2
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18653__B1 _16582_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14214__A1_N _14207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15467__B1 _15466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24832__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12554__A2_N _24867_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22971_ _22451_/A VGND VGND VPWR VPWR _22971_/X sky130_fd_sc_hd__buf_2
XFILLER_68_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24710_ _24704_/CLK _24710_/D HRESETn VGND VGND VPWR VPWR _24710_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11763__A _25526_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21922_ _21937_/A _21919_/X _21922_/C VGND VGND VPWR VPWR _21922_/X sky130_fd_sc_hd__and3_4
XFILLER_82_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16967__B1 _16073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24641_ _24641_/CLK _24641_/D HRESETn VGND VGND VPWR VPWR _23253_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21853_ _11986_/Y _12086_/X _12022_/Y _12057_/X VGND VGND VPWR VPWR _21853_/X sky130_fd_sc_hd__o22a_4
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22504__A2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20804_ _20780_/X _20803_/X _15566_/A _20784_/X VGND VGND VPWR VPWR _20804_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24572_ _24419_/CLK _16473_/X HRESETn VGND VGND VPWR VPWR _16472_/A sky130_fd_sc_hd__dfrtp_4
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21784_ _23686_/Q _21959_/B _23702_/Q _22397_/B VGND VGND VPWR VPWR _21784_/X sky130_fd_sc_hd__o22a_4
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23523_ _23525_/CLK _20051_/X VGND VGND VPWR VPWR _23523_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_223_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20735_ _20784_/A VGND VGND VPWR VPWR _20735_/X sky130_fd_sc_hd__buf_2
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23454_ _23456_/CLK _20232_/X VGND VGND VPWR VPWR _20231_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_149_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20666_ _23986_/Q _17394_/X _20665_/Y _20615_/A VGND VGND VPWR VPWR _20666_/X sky130_fd_sc_hd__a211o_4
XFILLER_183_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22405_ _22405_/A _21064_/B VGND VGND VPWR VPWR _22405_/X sky130_fd_sc_hd__or2_4
X_20597_ _14117_/Y _20543_/A _20556_/X _20596_/Y VGND VGND VPWR VPWR _20598_/A sky130_fd_sc_hd__a211o_4
X_23385_ _23388_/CLK _23385_/D VGND VGND VPWR VPWR _13427_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_176_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25124_ _23927_/CLK _25124_/D HRESETn VGND VGND VPWR VPWR _25124_/Q sky130_fd_sc_hd__dfrtp_4
X_22336_ _17720_/A _22336_/B VGND VGND VPWR VPWR _22336_/X sky130_fd_sc_hd__or2_4
XFILLER_164_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25055_ _25052_/CLK _14825_/X HRESETn VGND VGND VPWR VPWR _25055_/Q sky130_fd_sc_hd__dfrtp_4
X_22267_ _23400_/Q _22001_/Y _22051_/X _22266_/X VGND VGND VPWR VPWR _22268_/A sky130_fd_sc_hd__a211o_4
XFILLER_105_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _12014_/Y VGND VGND VPWR VPWR _12020_/X sky130_fd_sc_hd__buf_2
X_24006_ _24037_/CLK _24006_/D HRESETn VGND VGND VPWR VPWR _13113_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21218_ _21217_/X VGND VGND VPWR VPWR _21218_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18644__B1 _24520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22198_ _22209_/A _22198_/B VGND VGND VPWR VPWR _22200_/B sky130_fd_sc_hd__or2_4
XANTENNA__22440__B2 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17625__A _17625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21149_ _13503_/Y _21151_/A _21568_/B _21148_/Y VGND VGND VPWR VPWR _21149_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24573__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13971_ _14008_/A VGND VGND VPWR VPWR _14007_/C sky130_fd_sc_hd__inv_2
XFILLER_47_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24502__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15710_ HWDATA[30] VGND VGND VPWR VPWR _15710_/X sky130_fd_sc_hd__buf_2
XFILLER_58_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22743__A2 _21098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12922_ _12793_/A _12921_/Y VGND VGND VPWR VPWR _12924_/B sky130_fd_sc_hd__or2_4
X_24908_ _24907_/CLK _15597_/X HRESETn VGND VGND VPWR VPWR _24908_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19840__A _19835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16690_ _16689_/Y _16685_/X _15748_/X _16685_/X VGND VGND VPWR VPWR _16690_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15641_ _15644_/A VGND VGND VPWR VPWR _21296_/A sky130_fd_sc_hd__inv_2
XANTENNA__23362__A _23349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12853_ _12825_/X VGND VGND VPWR VPWR _12887_/A sky130_fd_sc_hd__inv_2
X_24839_ _24809_/CLK _24839_/D HRESETn VGND VGND VPWR VPWR _24839_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_160_0_HCLK clkbuf_7_80_0_HCLK/X VGND VGND VPWR VPWR _23747_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_3_0_HCLK clkbuf_7_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _11804_/A VGND VGND VPWR VPWR _13678_/A sky130_fd_sc_hd__inv_2
X_18360_ _18359_/X VGND VGND VPWR VPWR _18360_/Y sky130_fd_sc_hd__inv_2
XPHY_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15572_/A VGND VGND VPWR VPWR _15572_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_17_0_HCLK clkbuf_7_8_0_HCLK/X VGND VGND VPWR VPWR _23691_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _22130_/A VGND VGND VPWR VPWR _12784_/Y sky130_fd_sc_hd__inv_2
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17338_/A _17311_/B _17311_/C VGND VGND VPWR VPWR _24362_/D sky130_fd_sc_hd__and3_4
XPHY_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14523_/A _14060_/X VGND VGND VPWR VPWR _14523_/X sky130_fd_sc_hd__and2_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _16229_/A VGND VGND VPWR VPWR _11735_/X sky130_fd_sc_hd__buf_2
X_18291_ _18280_/C _17706_/X _18289_/X VGND VGND VPWR VPWR _24216_/D sky130_fd_sc_hd__o21a_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17241_/Y _17242_/B _17203_/A VGND VGND VPWR VPWR _17344_/A sky130_fd_sc_hd__or3_4
XFILLER_202_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14197__B1 _13785_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _25124_/Q VGND VGND VPWR VPWR _14454_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25361__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _12050_/A VGND VGND VPWR VPWR _11667_/B sky130_fd_sc_hd__inv_2
XFILLER_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13300_/A _13403_/X _13404_/X VGND VGND VPWR VPWR _13405_/X sky130_fd_sc_hd__and3_4
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17173_ _24622_/Q _17347_/C _16291_/Y _24367_/Q VGND VGND VPWR VPWR _17173_/X sky130_fd_sc_hd__a2bb2o_4
X_14385_ _14382_/Y _14383_/X _14384_/X _14373_/X VGND VGND VPWR VPWR _25149_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16933__A1_N _16126_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16124_ _16124_/A VGND VGND VPWR VPWR _16124_/X sky130_fd_sc_hd__buf_2
X_13336_ _13193_/A _13334_/X _13335_/X VGND VGND VPWR VPWR _13336_/X sky130_fd_sc_hd__and3_4
XANTENNA__23208__B1 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16055_ _14400_/A VGND VGND VPWR VPWR _16055_/X sky130_fd_sc_hd__buf_2
X_13267_ _13219_/X _13267_/B _13266_/X VGND VGND VPWR VPWR _13267_/X sky130_fd_sc_hd__and3_4
XFILLER_108_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15006_ _25010_/Q _24448_/Q _15273_/A _15005_/Y VGND VGND VPWR VPWR _15007_/D sky130_fd_sc_hd__o22a_4
X_12218_ _12234_/A _12216_/Y _12217_/Y _22150_/A VGND VGND VPWR VPWR _12228_/A sky130_fd_sc_hd__a2bb2o_4
X_13198_ _13249_/A VGND VGND VPWR VPWR _13199_/A sky130_fd_sc_hd__buf_2
X_19814_ _19805_/Y VGND VGND VPWR VPWR _19814_/X sky130_fd_sc_hd__buf_2
XFILLER_151_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12149_ _25166_/Q _12149_/B VGND VGND VPWR VPWR _12149_/X sky130_fd_sc_hd__or2_4
XFILLER_97_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20993__A1 sda_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21057__A _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19745_ _19745_/A VGND VGND VPWR VPWR _19745_/Y sky130_fd_sc_hd__inv_2
X_16957_ _16957_/A VGND VGND VPWR VPWR _16957_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24243__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15908_ _15908_/A _15907_/Y VGND VGND VPWR VPWR _15908_/X sky130_fd_sc_hd__and2_4
XFILLER_65_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19060__B1 _18965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19676_ _19675_/Y _19673_/X _19630_/X _19673_/X VGND VGND VPWR VPWR _23657_/D sky130_fd_sc_hd__a2bb2o_4
X_16888_ _16081_/Y _23320_/A _16081_/Y _23320_/A VGND VGND VPWR VPWR _16892_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18627_ _18627_/A _18622_/X _18627_/C _18626_/X VGND VGND VPWR VPWR _18627_/X sky130_fd_sc_hd__or4_4
X_15839_ _15773_/B _15836_/B VGND VGND VPWR VPWR _15839_/X sky130_fd_sc_hd__or2_4
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18558_ _18479_/B _18553_/B _18555_/B _18489_/X VGND VGND VPWR VPWR _18559_/A sky130_fd_sc_hd__a211o_4
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19363__B2 _19343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17509_ _17509_/A VGND VGND VPWR VPWR _17670_/A sky130_fd_sc_hd__inv_2
XFILLER_178_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18489_ _18823_/B VGND VGND VPWR VPWR _18489_/X sky130_fd_sc_hd__buf_2
XFILLER_220_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20520_ _20603_/A _20453_/D VGND VGND VPWR VPWR _20520_/X sky130_fd_sc_hd__and2_4
X_20451_ _25111_/Q _14490_/B _25112_/Q VGND VGND VPWR VPWR _20464_/C sky130_fd_sc_hd__or3_4
XANTENNA__21520__A _21843_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25031__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20382_ _20372_/X _19523_/Y _13459_/A _21216_/A _20369_/X VGND VGND VPWR VPWR _23394_/D
+ sky130_fd_sc_hd__a32o_4
X_23170_ _23170_/A _23063_/X VGND VGND VPWR VPWR _23170_/X sky130_fd_sc_hd__or2_4
XFILLER_173_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22121_ _22121_/A VGND VGND VPWR VPWR _22121_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22052_ _19580_/Y _22229_/B VGND VGND VPWR VPWR _22052_/X sky130_fd_sc_hd__and2_4
XFILLER_88_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14783__A1_N _18020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21003_ _21002_/A _21002_/B _24339_/Q _21002_/X VGND VGND VPWR VPWR _23972_/D sky130_fd_sc_hd__o22a_4
XFILLER_114_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12910__A1 _12741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12589__A _12588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22186__B1 _23968_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22954_ _15047_/A _23263_/B _23263_/C VGND VGND VPWR VPWR _22954_/X sky130_fd_sc_hd__and3_4
X_21905_ _21902_/A _19842_/Y VGND VGND VPWR VPWR _21905_/X sky130_fd_sc_hd__or2_4
XFILLER_16_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22885_ _23172_/A VGND VGND VPWR VPWR _22885_/X sky130_fd_sc_hd__buf_2
XFILLER_204_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23966__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_233_0_HCLK clkbuf_7_116_0_HCLK/X VGND VGND VPWR VPWR _24958_/CLK sky130_fd_sc_hd__clkbuf_1
X_24624_ _24618_/CLK _24624_/D HRESETn VGND VGND VPWR VPWR _24624_/Q sky130_fd_sc_hd__dfrtp_4
X_21836_ _21835_/Y _21159_/X _17424_/Y _17412_/X VGND VGND VPWR VPWR _21836_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12426__B1 _12390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25119__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24555_ _24555_/CLK _16516_/X HRESETn VGND VGND VPWR VPWR _24555_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16168__A1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21767_ _22381_/A _20147_/Y VGND VGND VPWR VPWR _21767_/X sky130_fd_sc_hd__or2_4
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21161__A1 _14229_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21133__C _13807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21161__B2 _21368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23506_ _23497_/CLK _23506_/D VGND VGND VPWR VPWR _23506_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13213__A _13199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20718_ _20718_/A VGND VGND VPWR VPWR _20718_/Y sky130_fd_sc_hd__inv_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24486_ _24486_/CLK _24486_/D HRESETn VGND VGND VPWR VPWR _24486_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_178_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21698_ _21698_/A _23002_/A VGND VGND VPWR VPWR _21698_/X sky130_fd_sc_hd__or2_4
XFILLER_184_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23437_ _23437_/CLK _23437_/D VGND VGND VPWR VPWR _20276_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20649_ _17392_/B _20648_/Y _20661_/C VGND VGND VPWR VPWR _20649_/X sky130_fd_sc_hd__and3_4
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16524__A _24552_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14170_ _14160_/A _14111_/X VGND VGND VPWR VPWR _14170_/Y sky130_fd_sc_hd__nand2_4
XFILLER_171_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23368_ _23368_/A VGND VGND VPWR VPWR IRQ[24] sky130_fd_sc_hd__buf_2
XFILLER_109_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18865__B1 _16485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20046__A _20034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13121_ _13121_/A _13121_/B _13121_/C _13121_/D VGND VGND VPWR VPWR _20754_/A sky130_fd_sc_hd__or4_4
X_25107_ _25117_/CLK _25107_/D HRESETn VGND VGND VPWR VPWR _25107_/Q sky130_fd_sc_hd__dfrtp_4
X_22319_ _22319_/A VGND VGND VPWR VPWR _22320_/D sky130_fd_sc_hd__inv_2
XANTENNA__19835__A _19835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23299_ _24545_/Q _23171_/X _22839_/X _23298_/X VGND VGND VPWR VPWR _23299_/X sky130_fd_sc_hd__a211o_4
XFILLER_106_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24754__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13052_ _13048_/A _13046_/B _13051_/Y VGND VGND VPWR VPWR _13052_/X sky130_fd_sc_hd__and3_4
X_25038_ _25015_/CLK _15171_/Y HRESETn VGND VGND VPWR VPWR _25038_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18617__B1 _16619_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22413__A1 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22413__B2 _22282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24324__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12003_ _12001_/A _11981_/A _12002_/Y VGND VGND VPWR VPWR _20968_/A sky130_fd_sc_hd__o21a_4
XFILLER_239_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12901__A1 _12766_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17355__A _17352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17860_ _16895_/X _17859_/X _17793_/A _17856_/B VGND VGND VPWR VPWR _17860_/X sky130_fd_sc_hd__a211o_4
XFILLER_120_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16811_ _16810_/Y _16808_/X _15725_/X _16808_/X VGND VGND VPWR VPWR _16811_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17791_ _17791_/A VGND VGND VPWR VPWR _17793_/A sky130_fd_sc_hd__buf_2
XFILLER_143_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19530_ _23704_/Q VGND VGND VPWR VPWR _19530_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13954_ _13954_/A _13907_/X _14234_/A VGND VGND VPWR VPWR _13955_/B sky130_fd_sc_hd__or3_4
X_16742_ _16741_/Y _16739_/X _15725_/X _16739_/X VGND VGND VPWR VPWR _16742_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_6_43_0_HCLK clkbuf_6_43_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_87_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12665__B1 _12641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12905_ _12838_/A _12904_/X VGND VGND VPWR VPWR _12905_/Y sky130_fd_sc_hd__nand2_4
X_16673_ _16668_/A VGND VGND VPWR VPWR _16673_/X sky130_fd_sc_hd__buf_2
X_19461_ _22235_/B _19458_/X _11906_/X _19458_/X VGND VGND VPWR VPWR _19461_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13885_ _13903_/A VGND VGND VPWR VPWR _13907_/A sky130_fd_sc_hd__inv_2
XANTENNA__18186__A _18014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18412_ _23074_/A _18411_/A _16202_/Y _18462_/B VGND VGND VPWR VPWR _18412_/X sky130_fd_sc_hd__o22a_4
X_12836_ _12895_/A VGND VGND VPWR VPWR _12836_/Y sky130_fd_sc_hd__inv_2
X_15624_ _15621_/Y _15622_/X _15623_/X _15622_/X VGND VGND VPWR VPWR _15624_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25542__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19392_ _18981_/A VGND VGND VPWR VPWR _19392_/X sky130_fd_sc_hd__buf_2
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15555_ _15549_/Y _15553_/X _15554_/X _15553_/X VGND VGND VPWR VPWR _15555_/X sky130_fd_sc_hd__a2bb2o_4
X_18343_ _13263_/A _18342_/X _13263_/A _18342_/X VGND VGND VPWR VPWR _18343_/X sky130_fd_sc_hd__a2bb2o_4
X_12767_ _22901_/A VGND VGND VPWR VPWR _12767_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21152__A1 _12111_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14495_/Y VGND VGND VPWR VPWR _14506_/X sky130_fd_sc_hd__buf_2
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ HWDATA[18] VGND VGND VPWR VPWR _11718_/X sky130_fd_sc_hd__buf_2
X_18274_ _18274_/A _20369_/A VGND VGND VPWR VPWR _18274_/X sky130_fd_sc_hd__or2_4
XFILLER_187_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15486_ _15489_/A VGND VGND VPWR VPWR _15486_/X sky130_fd_sc_hd__buf_2
XFILLER_147_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15906__A1 _14764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12698_ _12498_/Y _12701_/B _12641_/X VGND VGND VPWR VPWR _12698_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__12571__A1_N _12569_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14437_ _14431_/A VGND VGND VPWR VPWR _14437_/X sky130_fd_sc_hd__buf_2
X_17225_ _16343_/Y _24347_/Q _16352_/Y _17241_/A VGND VGND VPWR VPWR _17226_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16434__A HWDATA[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17156_ _16982_/Y _17151_/X VGND VGND VPWR VPWR _17157_/B sky130_fd_sc_hd__nand2_4
X_14368_ _14183_/X _14425_/B VGND VGND VPWR VPWR _14370_/B sky130_fd_sc_hd__or2_4
XANTENNA__22652__A1 _16539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16107_ _16106_/Y _16104_/X _11691_/X _16104_/X VGND VGND VPWR VPWR _16107_/X sky130_fd_sc_hd__a2bb2o_4
X_13319_ _13310_/X _13313_/X _13319_/C VGND VGND VPWR VPWR _13319_/X sky130_fd_sc_hd__or3_4
XFILLER_183_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17087_ _17087_/A VGND VGND VPWR VPWR _17105_/A sky130_fd_sc_hd__buf_2
X_14299_ _25177_/Q _14291_/X _25176_/Q _14296_/X VGND VGND VPWR VPWR _14299_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24495__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16038_ _16038_/A VGND VGND VPWR VPWR _16038_/X sky130_fd_sc_hd__buf_2
XANTENNA__18608__B1 _16578_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24424__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_125_0_HCLK clkbuf_6_62_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_251_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22955__A2 _22838_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16095__B1 _16001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17989_ _17984_/X _17986_/X _17988_/X VGND VGND VPWR VPWR _17989_/X sky130_fd_sc_hd__and3_4
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22707__A2 _22416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19728_ _11780_/A VGND VGND VPWR VPWR _19728_/X sky130_fd_sc_hd__buf_2
XFILLER_238_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21915__B1 _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19659_ _13303_/B VGND VGND VPWR VPWR _19659_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22670_ _22670_/A VGND VGND VPWR VPWR _22670_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21621_ _21901_/A _21613_/X _21620_/X VGND VGND VPWR VPWR _21621_/X sky130_fd_sc_hd__or3_4
XANTENNA__25212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24340_ _24340_/CLK _17402_/X HRESETn VGND VGND VPWR VPWR _21002_/A sky130_fd_sc_hd__dfstp_4
Xclkbuf_8_63_0_HCLK clkbuf_8_63_0_HCLK/A VGND VGND VPWR VPWR _24172_/CLK sky130_fd_sc_hd__clkbuf_1
X_21552_ _14414_/Y _14212_/A _14158_/Y _15457_/A VGND VGND VPWR VPWR _21554_/C sky130_fd_sc_hd__o22a_4
XFILLER_166_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22346__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20503_ _20503_/A _15451_/X _20503_/C VGND VGND VPWR VPWR _20503_/X sky130_fd_sc_hd__and3_4
X_24271_ _24686_/CLK _17845_/X HRESETn VGND VGND VPWR VPWR _17755_/A sky130_fd_sc_hd__dfrtp_4
X_21483_ _21656_/A _21483_/B _21483_/C VGND VGND VPWR VPWR _21483_/X sky130_fd_sc_hd__and3_4
XFILLER_119_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23222_ _24640_/Q _21528_/B VGND VGND VPWR VPWR _23222_/X sky130_fd_sc_hd__or2_4
XFILLER_153_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20434_ _20466_/B VGND VGND VPWR VPWR _20435_/B sky130_fd_sc_hd__inv_2
XANTENNA__18847__B1 _16510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23153_ _23044_/X _23151_/X _23046_/X _16006_/A _23152_/X VGND VGND VPWR VPWR _23153_/X
+ sky130_fd_sc_hd__a32o_4
X_20365_ _21480_/B _20362_/X _19620_/A _20362_/X VGND VGND VPWR VPWR _23403_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22104_ _22104_/A VGND VGND VPWR VPWR _22109_/B sky130_fd_sc_hd__inv_2
X_20296_ _21941_/B _20293_/X _19974_/X _20293_/X VGND VGND VPWR VPWR _23430_/D sky130_fd_sc_hd__a2bb2o_4
X_23084_ _24059_/Q _21303_/A _20793_/A _21598_/X VGND VGND VPWR VPWR _23084_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__24165__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20406__B1 _15643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14884__B2 _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22035_ _22016_/A _19969_/Y VGND VGND VPWR VPWR _22035_/X sky130_fd_sc_hd__or2_4
XFILLER_102_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15833__B1 _15472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23986_ _23986_/CLK _20667_/X HRESETn VGND VGND VPWR VPWR _23986_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_229_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22937_ _23072_/A _22926_/Y _22931_/X _22937_/D VGND VGND VPWR VPWR _22937_/X sky130_fd_sc_hd__or4_4
XFILLER_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13670_ _13670_/A _13669_/X VGND VGND VPWR VPWR _13670_/X sky130_fd_sc_hd__or2_4
X_22868_ _22194_/A VGND VGND VPWR VPWR _22868_/X sky130_fd_sc_hd__buf_2
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12621_ _12594_/Y _12503_/Y _12681_/A _12630_/B VGND VGND VPWR VPWR _12624_/B sky130_fd_sc_hd__or4_4
X_24607_ _24591_/CLK _24607_/D HRESETn VGND VGND VPWR VPWR _15085_/A sky130_fd_sc_hd__dfrtp_4
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21819_ _21815_/X _21818_/X _21686_/X VGND VGND VPWR VPWR _21819_/X sky130_fd_sc_hd__o21a_4
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22799_ _23128_/A VGND VGND VPWR VPWR _23072_/A sky130_fd_sc_hd__buf_2
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15340_ _24999_/Q _15340_/B VGND VGND VPWR VPWR _15341_/C sky130_fd_sc_hd__or2_4
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12552_ _12724_/A _12550_/Y _25406_/Q _12551_/Y VGND VGND VPWR VPWR _12557_/B sky130_fd_sc_hd__a2bb2o_4
X_24538_ _24539_/CLK _16563_/X HRESETn VGND VGND VPWR VPWR _24538_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16010__B1 _11685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15271_ _15271_/A VGND VGND VPWR VPWR _25012_/D sky130_fd_sc_hd__inv_2
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _12480_/A _12476_/B _12483_/C VGND VGND VPWR VPWR _12483_/X sky130_fd_sc_hd__and3_4
X_24469_ _25021_/CLK _16742_/X HRESETn VGND VGND VPWR VPWR _24469_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24935__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ _15993_/Y _24403_/Q _15993_/Y _24403_/Q VGND VGND VPWR VPWR _17010_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ _25197_/Q VGND VGND VPWR VPWR _14222_/Y sky130_fd_sc_hd__inv_2
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18838__B1 _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22634__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14153_ _14113_/X _14152_/Y _14102_/C _14113_/X VGND VGND VPWR VPWR _25214_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_5_27_0_HCLK_A clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17510__B1 _11755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13104_ _12983_/D _13005_/D _12998_/A _13101_/Y VGND VGND VPWR VPWR _13105_/A sky130_fd_sc_hd__a211o_4
XFILLER_3_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14084_ _20987_/B VGND VGND VPWR VPWR _14084_/Y sky130_fd_sc_hd__inv_2
X_18961_ _18959_/Y _18960_/X _17421_/X _18960_/X VGND VGND VPWR VPWR _23904_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13035_ _25356_/Q _13035_/B VGND VGND VPWR VPWR _13035_/X sky130_fd_sc_hd__or2_4
X_17912_ _21993_/A VGND VGND VPWR VPWR _17912_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17085__A _17381_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18892_ _18871_/X _18885_/X _24120_/Q _24121_/Q _18888_/X VGND VGND VPWR VPWR _18892_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12886__B1 _12804_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17843_ _17755_/A _17843_/B VGND VGND VPWR VPWR _17843_/X sky130_fd_sc_hd__or2_4
XANTENNA__14859__D _14817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14627__A1 _13525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17540__A1_N _11694_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15824__B1 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17774_ _17766_/X _17773_/X VGND VGND VPWR VPWR _17775_/C sky130_fd_sc_hd__or2_4
X_14986_ _14986_/A VGND VGND VPWR VPWR _14986_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19513_ _21814_/B _19508_/X _11920_/X _19508_/X VGND VGND VPWR VPWR _19513_/X sky130_fd_sc_hd__a2bb2o_4
X_16725_ _16725_/A VGND VGND VPWR VPWR _16726_/A sky130_fd_sc_hd__buf_2
X_13937_ _13937_/A VGND VGND VPWR VPWR _13937_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24082__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23253__C _22817_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22570__B1 _21832_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16429__A _24584_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12338__A2_N _24834_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19444_ _19444_/A VGND VGND VPWR VPWR _19444_/Y sky130_fd_sc_hd__inv_2
X_13868_ _13860_/X _13867_/X _25187_/Q _13845_/Y VGND VGND VPWR VPWR _13868_/X sky130_fd_sc_hd__o22a_4
X_16656_ _16654_/Y _16655_/X _16295_/X _16655_/X VGND VGND VPWR VPWR _16656_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17251__C _17251_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12819_ _12845_/C _24815_/Q _12845_/C _24815_/Q VGND VGND VPWR VPWR _12823_/B sky130_fd_sc_hd__a2bb2o_4
X_15607_ _15607_/A VGND VGND VPWR VPWR _22566_/A sky130_fd_sc_hd__inv_2
XFILLER_50_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19375_ _19374_/Y _19372_/X _19351_/X _19372_/X VGND VGND VPWR VPWR _19375_/X sky130_fd_sc_hd__a2bb2o_4
X_13799_ _13796_/Y _13792_/X _13798_/X _13792_/X VGND VGND VPWR VPWR _25271_/D sky130_fd_sc_hd__a2bb2o_4
X_16587_ _24528_/Q VGND VGND VPWR VPWR _16587_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18326_ _20220_/A _18326_/B _18326_/C _20220_/D VGND VGND VPWR VPWR _20054_/B sky130_fd_sc_hd__and4_4
X_15538_ _15537_/Y _15533_/X HADDR[0] _15533_/X VGND VGND VPWR VPWR _24925_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15987__B _15986_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13788__A _14392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15469_ _14392_/A VGND VGND VPWR VPWR _15469_/X sky130_fd_sc_hd__buf_2
X_18257_ _11780_/A VGND VGND VPWR VPWR _18257_/X sky130_fd_sc_hd__buf_2
XFILLER_129_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24676__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17208_ _17201_/X _17208_/B _17208_/C _17208_/D VGND VGND VPWR VPWR _17227_/A sky130_fd_sc_hd__or4_4
XFILLER_175_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18188_ _18124_/A _18184_/X _18187_/X VGND VGND VPWR VPWR _18196_/B sky130_fd_sc_hd__or3_4
XANTENNA__24605__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17139_ _16971_/Y _17129_/X VGND VGND VPWR VPWR _17140_/C sky130_fd_sc_hd__nand2_4
X_20150_ _20137_/Y VGND VGND VPWR VPWR _20150_/X sky130_fd_sc_hd__buf_2
XFILLER_170_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20081_ _20081_/A VGND VGND VPWR VPWR _21412_/B sky130_fd_sc_hd__inv_2
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16068__B1 _15469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23338__C1 _23337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15815__B1 _24834_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23840_ _23846_/CLK _23840_/D VGND VGND VPWR VPWR _19148_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__13028__A _13028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16134__A1_N _16133_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23771_ _23889_/CLK _23771_/D VGND VGND VPWR VPWR _23771_/Q sky130_fd_sc_hd__dfxtp_4
X_20983_ _24121_/Q _20982_/B _24120_/Q _20982_/X VGND VGND VPWR VPWR _20983_/X sky130_fd_sc_hd__o22a_4
XANTENNA__12867__A _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25510_ _25510_/CLK _25510_/D HRESETn VGND VGND VPWR VPWR _19964_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22722_ _24762_/Q _22274_/X _15958_/A _24834_/Q _21833_/X VGND VGND VPWR VPWR _22723_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_214_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25441_ _25444_/CLK _12474_/Y HRESETn VGND VGND VPWR VPWR _25441_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22653_ _22141_/X _22652_/X VGND VGND VPWR VPWR _22665_/B sky130_fd_sc_hd__and2_4
XFILLER_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21116__A1 _21077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21604_ _22221_/A VGND VGND VPWR VPWR _21775_/A sky130_fd_sc_hd__buf_2
X_25372_ _25369_/CLK _12957_/Y HRESETn VGND VGND VPWR VPWR _12806_/A sky130_fd_sc_hd__dfrtp_4
X_22584_ _22584_/A _22735_/B VGND VGND VPWR VPWR _22584_/X sky130_fd_sc_hd__and2_4
XFILLER_159_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24323_ _23425_/CLK _17489_/Y HRESETn VGND VGND VPWR VPWR _21220_/A sky130_fd_sc_hd__dfrtp_4
X_21535_ _16637_/A _21534_/X _21436_/X _24822_/Q _21336_/X VGND VGND VPWR VPWR _21535_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_166_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24254_ _24257_/CLK _24254_/D HRESETn VGND VGND VPWR VPWR _21993_/A sky130_fd_sc_hd__dfrtp_4
X_21466_ _21466_/A VGND VGND VPWR VPWR _21662_/A sky130_fd_sc_hd__buf_2
XANTENNA__24346__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_7_0_HCLK clkbuf_6_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23205_ _23169_/A _23204_/Y VGND VGND VPWR VPWR _23205_/Y sky130_fd_sc_hd__nor2_4
X_20417_ _23381_/Q VGND VGND VPWR VPWR _21897_/B sky130_fd_sc_hd__inv_2
X_24185_ _24675_/CLK _18506_/X HRESETn VGND VGND VPWR VPWR _24185_/Q sky130_fd_sc_hd__dfrtp_4
X_21397_ _22202_/A _21397_/B VGND VGND VPWR VPWR _21397_/X sky130_fd_sc_hd__or2_4
XFILLER_175_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22523__B _22523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23136_ _23209_/A _23132_/X _23135_/X VGND VGND VPWR VPWR _23142_/C sky130_fd_sc_hd__and3_4
XFILLER_1_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20348_ _18276_/X _19960_/X _19479_/X VGND VGND VPWR VPWR _20348_/X sky130_fd_sc_hd__or3_4
XFILLER_162_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23067_ _23209_/A _23064_/X _23066_/X VGND VGND VPWR VPWR _23072_/C sky130_fd_sc_hd__and3_4
X_20279_ _20266_/Y VGND VGND VPWR VPWR _20279_/X sky130_fd_sc_hd__buf_2
XANTENNA__21052__B1 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22018_ _22013_/X _22017_/X _21489_/X VGND VGND VPWR VPWR _22018_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_88_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13583__D _13765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23981__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14840_ _14826_/A VGND VGND VPWR VPWR _14840_/X sky130_fd_sc_hd__buf_2
XFILLER_208_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14771_ _14769_/B _14769_/C VGND VGND VPWR VPWR _14771_/X sky130_fd_sc_hd__and2_4
XFILLER_17_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17352__B _17352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11983_ _11976_/Y _11983_/B VGND VGND VPWR VPWR _11983_/Y sky130_fd_sc_hd__nor2_4
X_23969_ _25243_/CLK _21005_/X HRESETn VGND VGND VPWR VPWR _23969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13722_ _13721_/Y VGND VGND VPWR VPWR _13723_/A sky130_fd_sc_hd__buf_2
X_16510_ _16510_/A VGND VGND VPWR VPWR _16510_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17490_ _11746_/Y _24302_/Q _11746_/Y _24302_/Q VGND VGND VPWR VPWR _17490_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16231__B1 _16229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12496__B _13028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23370__A _21017_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13653_ _24060_/Q _24059_/Q _13635_/X _20932_/B VGND VGND VPWR VPWR _13653_/X sky130_fd_sc_hd__or4_4
X_16441_ _18560_/A VGND VGND VPWR VPWR _16441_/X sky130_fd_sc_hd__buf_2
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12604_ _12692_/A _12569_/Y _12716_/A _12689_/A VGND VGND VPWR VPWR _12605_/C sky130_fd_sc_hd__or4_4
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _24610_/Q VGND VGND VPWR VPWR _16372_/Y sky130_fd_sc_hd__inv_2
X_19160_ _23835_/Q VGND VGND VPWR VPWR _19160_/Y sky130_fd_sc_hd__inv_2
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ _19570_/A _14422_/A VGND VGND VPWR VPWR _13584_/X sky130_fd_sc_hd__or2_4
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15323_ _15323_/A _15303_/X VGND VGND VPWR VPWR _15324_/A sky130_fd_sc_hd__or2_4
X_18111_ _17972_/A _18111_/B VGND VGND VPWR VPWR _18111_/X sky130_fd_sc_hd__or2_4
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ _12623_/A _24884_/Q _12624_/A _12534_/Y VGND VGND VPWR VPWR _12535_/X sky130_fd_sc_hd__o22a_4
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19091_ _19852_/A VGND VGND VPWR VPWR _19091_/X sky130_fd_sc_hd__buf_2
XFILLER_173_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13401__A _13433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15254_ _15254_/A _15254_/B VGND VGND VPWR VPWR _15254_/X sky130_fd_sc_hd__or2_4
X_18042_ _18227_/A _18038_/X _18042_/C VGND VGND VPWR VPWR _18042_/X sky130_fd_sc_hd__or3_4
XFILLER_157_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12466_ _12267_/Y _12465_/X _12398_/X _12461_/Y VGND VGND VPWR VPWR _12466_/X sky130_fd_sc_hd__a211o_4
XFILLER_144_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15888__A3 _16240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24087__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22714__A _22714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14205_ _20678_/A VGND VGND VPWR VPWR _14205_/Y sky130_fd_sc_hd__inv_2
X_15185_ _15185_/A _15180_/Y _15184_/X VGND VGND VPWR VPWR _15185_/X sky130_fd_sc_hd__or3_4
XFILLER_172_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24016__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12397_ _12413_/A _12395_/X _12396_/X VGND VGND VPWR VPWR _25460_/D sky130_fd_sc_hd__and3_4
X_14136_ _14105_/A _14105_/B _14105_/A _14105_/B VGND VGND VPWR VPWR _14137_/A sky130_fd_sc_hd__a2bb2o_4
X_19993_ _23545_/Q VGND VGND VPWR VPWR _19993_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14067_ _14067_/A VGND VGND VPWR VPWR _14067_/X sky130_fd_sc_hd__buf_2
X_18944_ _18944_/A VGND VGND VPWR VPWR _18944_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13018_ _12308_/Y _13017_/X VGND VGND VPWR VPWR _13018_/X sky130_fd_sc_hd__or2_4
XFILLER_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12323__A2 _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18875_ _18875_/A _18874_/X VGND VGND VPWR VPWR _18875_/X sky130_fd_sc_hd__or2_4
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21594__A1 _21597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18639__A _24143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17826_ _17761_/A _17826_/B VGND VGND VPWR VPWR _17826_/Y sky130_fd_sc_hd__nand2_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23335__A2 _22282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15812__A3 _15735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21065__A _15661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17757_ _17757_/A VGND VGND VPWR VPWR _17757_/Y sky130_fd_sc_hd__inv_2
X_14969_ _14960_/X _14969_/B _14969_/C _14968_/X VGND VGND VPWR VPWR _14969_/X sky130_fd_sc_hd__or4_4
XFILLER_82_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_13_0_HCLK clkbuf_4_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__16159__A _21521_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16708_ _16708_/A VGND VGND VPWR VPWR _16708_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17688_ _17668_/B _17688_/B _17688_/C VGND VGND VPWR VPWR _24296_/D sky130_fd_sc_hd__and3_4
XFILLER_222_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19427_ _19425_/Y _19426_/X _19357_/X _19426_/X VGND VGND VPWR VPWR _23741_/D sky130_fd_sc_hd__a2bb2o_4
X_16639_ _16639_/A VGND VGND VPWR VPWR _16639_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12837__D _12813_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24857__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19358_ _19355_/Y _19356_/X _19357_/X _19356_/X VGND VGND VPWR VPWR _19358_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18309_ _21189_/A VGND VGND VPWR VPWR _21920_/A sky130_fd_sc_hd__buf_2
X_19289_ _23789_/Q VGND VGND VPWR VPWR _19289_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14407__A _14407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21320_ _24036_/Q _21315_/X _21318_/X _21319_/X VGND VGND VPWR VPWR _21320_/X sky130_fd_sc_hd__a211o_4
XFILLER_163_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_137_0_HCLK clkbuf_7_68_0_HCLK/X VGND VGND VPWR VPWR _23754_/CLK sky130_fd_sc_hd__clkbuf_1
X_21251_ _21627_/A _21249_/X _21251_/C VGND VGND VPWR VPWR _21251_/X sky130_fd_sc_hd__and3_4
XFILLER_209_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20202_ _20198_/Y _20201_/X _18250_/X _20201_/X VGND VGND VPWR VPWR _20202_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21282__B1 _21178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21182_ _24213_/Q VGND VGND VPWR VPWR _21204_/A sky130_fd_sc_hd__inv_2
XFILLER_104_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20133_ _19852_/A VGND VGND VPWR VPWR _20133_/X sky130_fd_sc_hd__buf_2
XANTENNA__19227__B1 _19203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20064_ _20054_/A _18328_/A _13459_/A _13431_/B _20055_/A VGND VGND VPWR VPWR _20064_/X
+ sky130_fd_sc_hd__a32o_4
X_24941_ _25510_/CLK _24941_/D HRESETn VGND VGND VPWR VPWR _24941_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_225_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22782__B1 _24274_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24872_ _24872_/CLK _15734_/X HRESETn VGND VGND VPWR VPWR _24872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23823_ _23831_/CLK _19195_/X VGND VGND VPWR VPWR _23823_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16069__A _24718_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23754_ _23754_/CLK _19390_/X VGND VGND VPWR VPWR _17955_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ _11995_/X _13506_/A VGND VGND VPWR VPWR _24094_/D sky130_fd_sc_hd__and2_4
XPHY_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16213__B1 _15946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _22705_/A _22701_/B VGND VGND VPWR VPWR _22705_/X sky130_fd_sc_hd__or2_4
XPHY_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21703__A _22716_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23685_ _23425_/CLK _23685_/D VGND VGND VPWR VPWR _23685_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _20892_/X _20895_/Y _16679_/A _20896_/X VGND VGND VPWR VPWR _24050_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_198_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24598__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25424_ _24872_/CLK _12648_/X HRESETn VGND VGND VPWR VPWR _12560_/A sky130_fd_sc_hd__dfrtp_4
X_22636_ _21305_/B _22635_/X _21312_/X _16042_/A _21708_/X VGND VGND VPWR VPWR _22636_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24527__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25355_ _25346_/CLK _25355_/D HRESETn VGND VGND VPWR VPWR _25355_/Q sky130_fd_sc_hd__dfrtp_4
X_22567_ _16691_/Y _22641_/B VGND VGND VPWR VPWR _22567_/X sky130_fd_sc_hd__and2_4
XFILLER_10_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_33_0_HCLK clkbuf_7_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_67_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12320_ _25344_/Q _24829_/Q _13074_/A _12319_/Y VGND VGND VPWR VPWR _12327_/B sky130_fd_sc_hd__o22a_4
X_24306_ _24310_/CLK _17652_/X HRESETn VGND VGND VPWR VPWR _24306_/Q sky130_fd_sc_hd__dfrtp_4
X_21518_ _21321_/X _21419_/X _21518_/C _21518_/D VGND VGND VPWR VPWR HRDATA[1] sky130_fd_sc_hd__or4_4
XFILLER_139_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_96_0_HCLK clkbuf_7_97_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_96_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_25286_ _25292_/CLK _25286_/D HRESETn VGND VGND VPWR VPWR _11823_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_155_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24180__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22498_ _22781_/A _22480_/X _22498_/C _22497_/X VGND VGND VPWR VPWR _22498_/X sky130_fd_sc_hd__or4_4
X_12251_ _12251_/A VGND VGND VPWR VPWR _12269_/A sky130_fd_sc_hd__inv_2
X_24237_ _24341_/CLK _18246_/X HRESETn VGND VGND VPWR VPWR _24237_/Q sky130_fd_sc_hd__dfrtp_4
X_21449_ _17880_/A _21447_/X _12492_/A _21448_/X VGND VGND VPWR VPWR _21449_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17628__A _17559_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23933__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16656__A1_N _16654_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12182_ _23184_/A VGND VGND VPWR VPWR _12182_/Y sky130_fd_sc_hd__inv_2
X_24168_ _24650_/CLK _18572_/X HRESETn VGND VGND VPWR VPWR _18400_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17347__B _17352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23119_ _22686_/A VGND VGND VPWR VPWR _23235_/A sky130_fd_sc_hd__buf_2
XANTENNA__23014__A1 _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25386__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_16990_ _16990_/A VGND VGND VPWR VPWR _17041_/C sky130_fd_sc_hd__inv_2
X_24099_ _23951_/CLK MSI_S2 HRESETn VGND VGND VPWR VPWR _24099_/Q sky130_fd_sc_hd__dfrtp_4
X_15941_ _15923_/X _15928_/X HWDATA[23] _23036_/A _15926_/X VGND VGND VPWR VPWR _24771_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23365__A _21012_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20181__A2_N _20180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17363__A _17366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18660_ _24148_/Q VGND VGND VPWR VPWR _18728_/A sky130_fd_sc_hd__inv_2
X_15872_ _15861_/X VGND VGND VPWR VPWR _15872_/X sky130_fd_sc_hd__buf_2
X_17611_ _17584_/X _17602_/X _17585_/A VGND VGND VPWR VPWR _17612_/C sky130_fd_sc_hd__o21a_4
X_14823_ _14805_/A VGND VGND VPWR VPWR _14823_/X sky130_fd_sc_hd__buf_2
X_18591_ _18591_/A _18591_/B _18593_/C VGND VGND VPWR VPWR _18591_/X sky130_fd_sc_hd__and3_4
XFILLER_76_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17542_ _11772_/Y _24295_/Q _17561_/A _17541_/Y VGND VGND VPWR VPWR _17542_/X sky130_fd_sc_hd__a2bb2o_4
X_11966_ _11934_/A _11932_/X _11963_/X _11931_/A _11965_/X VGND VGND VPWR VPWR _25499_/D
+ sky130_fd_sc_hd__a32o_4
X_14754_ _14753_/X _14740_/Y _14747_/X VGND VGND VPWR VPWR _25061_/D sky130_fd_sc_hd__a21oi_4
XFILLER_91_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16204__B1 _15939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13705_ _11814_/Y _13673_/X VGND VGND VPWR VPWR _13705_/Y sky130_fd_sc_hd__nand2_4
XFILLER_60_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14685_ _14684_/X VGND VGND VPWR VPWR _14685_/Y sky130_fd_sc_hd__inv_2
X_17473_ _17443_/X VGND VGND VPWR VPWR _17473_/Y sky130_fd_sc_hd__inv_2
X_11897_ _11897_/A VGND VGND VPWR VPWR _11897_/X sky130_fd_sc_hd__buf_2
XFILLER_204_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24950__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19212_ _19207_/Y _19211_/X _19144_/X _19211_/X VGND VGND VPWR VPWR _23818_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_220_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13636_ _24052_/Q _24053_/Q _24051_/Q _13636_/D VGND VGND VPWR VPWR _13637_/D sky130_fd_sc_hd__or4_4
X_16424_ _15094_/Y _16422_/X _16145_/X _16422_/X VGND VGND VPWR VPWR _16424_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24268__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19143_ _19149_/A VGND VGND VPWR VPWR _19143_/X sky130_fd_sc_hd__buf_2
XFILLER_9_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22147__C _22146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13567_ _13567_/A VGND VGND VPWR VPWR _22540_/A sky130_fd_sc_hd__inv_2
X_16355_ _24614_/Q VGND VGND VPWR VPWR _16355_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12241__B2 _12178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12518_ _12689_/A _24855_/Q _12689_/A _24855_/Q VGND VGND VPWR VPWR _12519_/D sky130_fd_sc_hd__a2bb2o_4
X_15306_ _15308_/B VGND VGND VPWR VPWR _15307_/B sky130_fd_sc_hd__inv_2
X_16286_ _16283_/Y _16279_/X _15996_/X _16285_/X VGND VGND VPWR VPWR _24641_/D sky130_fd_sc_hd__a2bb2o_4
X_19074_ _19074_/A VGND VGND VPWR VPWR _19074_/X sky130_fd_sc_hd__buf_2
X_13498_ _13498_/A VGND VGND VPWR VPWR _13498_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17180__B2 _17179_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18025_ _17966_/X _18023_/X _24248_/Q _18024_/X VGND VGND VPWR VPWR _18025_/X sky130_fd_sc_hd__o22a_4
X_12449_ _12448_/X VGND VGND VPWR VPWR _12450_/B sky130_fd_sc_hd__inv_2
X_15237_ _15204_/A _15234_/X VGND VGND VPWR VPWR _15237_/X sky130_fd_sc_hd__or2_4
XFILLER_161_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16442__A _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15168_ _15168_/A _15168_/B _15168_/C VGND VGND VPWR VPWR _15168_/X sky130_fd_sc_hd__or3_4
X_14119_ _14115_/X _14116_/X _14117_/Y _14118_/X VGND VGND VPWR VPWR _14119_/X sky130_fd_sc_hd__o22a_4
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15099_ _24983_/Q VGND VGND VPWR VPWR _15294_/C sky130_fd_sc_hd__inv_2
X_19976_ _19976_/A VGND VGND VPWR VPWR _19976_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18927_ _18927_/A VGND VGND VPWR VPWR _18927_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25056__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18858_ _24571_/Q _18730_/A _24571_/Q _18730_/A VGND VGND VPWR VPWR _18861_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17704__C _17704_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17809_ _17808_/X VGND VGND VPWR VPWR _17809_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18789_ _18789_/A _18797_/A _18789_/C _18797_/B VGND VGND VPWR VPWR _18789_/X sky130_fd_sc_hd__or4_4
X_20820_ _20690_/X _20819_/X _24923_/Q _20735_/X VGND VGND VPWR VPWR _20820_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21523__A _21232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20751_ _20748_/Y _20749_/Y _20750_/X VGND VGND VPWR VPWR _20751_/X sky130_fd_sc_hd__o21a_4
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24691__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16617__A _24516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23470_ _23487_/CLK _20190_/X VGND VGND VPWR VPWR _20189_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20682_ _20485_/X _20503_/C _20613_/B VGND VGND VPWR VPWR _23995_/D sky130_fd_sc_hd__o21a_4
XANTENNA__14444__A1_N _20600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24620__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22421_ _22294_/X _22420_/X _22296_/X _24862_/Q _22282_/A VGND VGND VPWR VPWR _22422_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_148_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25140_ _25140_/CLK _14416_/X HRESETn VGND VGND VPWR VPWR _14414_/A sky130_fd_sc_hd__dfstp_4
X_22352_ _21933_/A _22350_/X _22351_/X VGND VGND VPWR VPWR _22352_/X sky130_fd_sc_hd__and3_4
X_21303_ _21303_/A VGND VGND VPWR VPWR _21303_/X sky130_fd_sc_hd__buf_2
X_25071_ _23735_/CLK _14662_/X HRESETn VGND VGND VPWR VPWR _13600_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17448__A _17448_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22283_ _22279_/X _22281_/X _21306_/C _24722_/Q _22282_/X VGND VGND VPWR VPWR _22283_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19448__B1 _19357_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16352__A _24615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24022_ _24051_/CLK _20775_/Y HRESETn VGND VGND VPWR VPWR _24022_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21234_ _21128_/B _21231_/X _21232_/X _21233_/Y VGND VGND VPWR VPWR _21235_/C sky130_fd_sc_hd__a211o_4
X_21165_ _16619_/Y _11700_/A VGND VGND VPWR VPWR _21168_/B sky130_fd_sc_hd__or2_4
XFILLER_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20116_ _20116_/A VGND VGND VPWR VPWR _20116_/X sky130_fd_sc_hd__buf_2
XFILLER_132_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21096_ _21085_/X _21096_/B _21096_/C VGND VGND VPWR VPWR _21096_/X sky130_fd_sc_hd__and3_4
XANTENNA__20602__A _14391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18423__A1 _22883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20047_ _21634_/B _20046_/X _19824_/X _20046_/X VGND VGND VPWR VPWR _23525_/D sky130_fd_sc_hd__a2bb2o_4
X_24924_ _24910_/CLK _15548_/X HRESETn VGND VGND VPWR VPWR _23324_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24855_ _24855_/CLK _24855_/D HRESETn VGND VGND VPWR VPWR _24855_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15788__A2 _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16985__A1 _24734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24779__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11820_/A VGND VGND VPWR VPWR _11820_/Y sky130_fd_sc_hd__inv_2
XPHY_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23806_ _23806_/CLK _23806_/D VGND VGND VPWR VPWR _19242_/A sky130_fd_sc_hd__dfxtp_4
X_24786_ _24795_/CLK _15902_/X HRESETn VGND VGND VPWR VPWR _21425_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _21995_/Y _21996_/X _21984_/X _21997_/X VGND VGND VPWR VPWR _23346_/B sky130_fd_sc_hd__a211o_4
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24708__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21433__A _15851_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11699_/X _11707_/X _15965_/A _25530_/Q _11708_/X VGND VGND VPWR VPWR _25530_/D
+ sky130_fd_sc_hd__a32o_4
X_23737_ _23735_/CLK _19438_/X VGND VGND VPWR VPWR _17992_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_242_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20949_ _20948_/Y _20949_/B VGND VGND VPWR VPWR _20949_/X sky130_fd_sc_hd__and2_4
XPHY_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16527__A _16527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _25118_/Q VGND VGND VPWR VPWR _21846_/A sky130_fd_sc_hd__inv_2
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11681_/X VGND VGND VPWR VPWR _11682_/Y sky130_fd_sc_hd__inv_2
X_23668_ _25326_/CLK _19644_/X VGND VGND VPWR VPWR _13407_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_81_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24361__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13421_/A _19113_/A VGND VGND VPWR VPWR _13422_/C sky130_fd_sc_hd__or2_4
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22619_ _13533_/Y _22619_/B VGND VGND VPWR VPWR _22619_/X sky130_fd_sc_hd__and2_4
X_25407_ _25403_/CLK _25407_/D HRESETn VGND VGND VPWR VPWR _25407_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23599_ _23575_/CLK _19843_/X VGND VGND VPWR VPWR _19842_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16140_ _22494_/A VGND VGND VPWR VPWR _16140_/Y sky130_fd_sc_hd__inv_2
X_13352_ _13310_/X _13348_/X _13352_/C VGND VGND VPWR VPWR _13352_/X sky130_fd_sc_hd__or3_4
X_25338_ _25341_/CLK _25338_/D HRESETn VGND VGND VPWR VPWR _25338_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12303_ _24839_/Q VGND VGND VPWR VPWR _12303_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16071_ _24717_/Q VGND VGND VPWR VPWR _16071_/Y sky130_fd_sc_hd__inv_2
X_13283_ _13186_/X _13282_/X _25331_/Q _13245_/X VGND VGND VPWR VPWR _13283_/X sky130_fd_sc_hd__o22a_4
X_25269_ _24172_/CLK _25269_/D HRESETn VGND VGND VPWR VPWR _13549_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_127_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17358__A _17358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23079__B _22817_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15022_ _15022_/A VGND VGND VPWR VPWR _15022_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_120_0_HCLK clkbuf_7_60_0_HCLK/X VGND VGND VPWR VPWR _24819_/CLK sky130_fd_sc_hd__clkbuf_1
X_12234_ _12234_/A VGND VGND VPWR VPWR _12428_/B sky130_fd_sc_hd__inv_2
XFILLER_154_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_183_0_HCLK clkbuf_7_91_0_HCLK/X VGND VGND VPWR VPWR _23926_/CLK sky130_fd_sc_hd__clkbuf_1
X_19830_ _21238_/B _19823_/X _19091_/X _19805_/Y VGND VGND VPWR VPWR _19830_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12165_ _25444_/Q VGND VGND VPWR VPWR _12266_/A sky130_fd_sc_hd__inv_2
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19761_ _19761_/A VGND VGND VPWR VPWR _19761_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12096_ _12119_/A _12090_/X _11761_/X _12095_/X VGND VGND VPWR VPWR _12096_/X sky130_fd_sc_hd__a2bb2o_4
X_16973_ _24397_/Q VGND VGND VPWR VPWR _16973_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13487__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22746__B1 _24870_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18712_ _18707_/B _18699_/X VGND VGND VPWR VPWR _18713_/A sky130_fd_sc_hd__or2_4
X_15924_ _15781_/A _15855_/B VGND VGND VPWR VPWR _15924_/X sky130_fd_sc_hd__or2_4
X_19692_ _20052_/A _18911_/B _20387_/C VGND VGND VPWR VPWR _19693_/A sky130_fd_sc_hd__or3_4
XANTENNA__21327__B _21327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16425__B1 _16055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18643_ _18643_/A VGND VGND VPWR VPWR _18804_/A sky130_fd_sc_hd__buf_2
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15855_ _15698_/A _15855_/B VGND VGND VPWR VPWR _15881_/A sky130_fd_sc_hd__or2_4
XFILLER_225_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16976__A1 _24723_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14806_ _14830_/A VGND VGND VPWR VPWR _14806_/X sky130_fd_sc_hd__buf_2
X_18574_ _18572_/A _18567_/X _18574_/C VGND VGND VPWR VPWR _18574_/X sky130_fd_sc_hd__and3_4
XANTENNA__14987__B1 _25013_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15786_ _15811_/A VGND VGND VPWR VPWR _15786_/X sky130_fd_sc_hd__buf_2
XANTENNA__24449__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12998_ _12998_/A _12998_/B _12997_/X VGND VGND VPWR VPWR _12999_/A sky130_fd_sc_hd__or3_4
X_17525_ _17518_/X _17520_/X _17525_/C _17525_/D VGND VGND VPWR VPWR _17526_/D sky130_fd_sc_hd__or4_4
XANTENNA__21343__A _21343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14737_ _22044_/A VGND VGND VPWR VPWR _14737_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11949_ _11948_/X VGND VGND VPWR VPWR _11950_/A sky130_fd_sc_hd__buf_2
XANTENNA__12965__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24211__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22158__B _22127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17456_ _17451_/X _17453_/X _18342_/A _17455_/Y VGND VGND VPWR VPWR _17459_/A sky130_fd_sc_hd__o22a_4
X_14668_ _25061_/Q VGND VGND VPWR VPWR _14668_/X sky130_fd_sc_hd__buf_2
X_16407_ _16404_/Y _16406_/X _16320_/X _16406_/X VGND VGND VPWR VPWR _24596_/D sky130_fd_sc_hd__a2bb2o_4
X_13619_ _19117_/A _13618_/X _19117_/A _13618_/X VGND VGND VPWR VPWR _13620_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_177_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17387_ _20630_/A _17386_/X VGND VGND VPWR VPWR _17388_/B sky130_fd_sc_hd__or2_4
XANTENNA__24031__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14599_ _25084_/Q _25083_/Q VGND VGND VPWR VPWR _14599_/X sky130_fd_sc_hd__or2_4
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19126_ _19133_/A VGND VGND VPWR VPWR _19126_/X sky130_fd_sc_hd__buf_2
X_16338_ _16336_/Y _16332_/X _16141_/X _16337_/X VGND VGND VPWR VPWR _24621_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19057_ _18942_/A VGND VGND VPWR VPWR _19057_/X sky130_fd_sc_hd__buf_2
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23226__A1 _22552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16269_ _15642_/X _15986_/Y _16267_/X _21013_/A _16268_/X VGND VGND VPWR VPWR _16269_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__23226__B2 _22555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16172__A _13577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16900__B2 _21059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18008_ _18123_/A _18008_/B _18007_/X VGND VGND VPWR VPWR _18009_/C sky130_fd_sc_hd__and3_4
XANTENNA__25237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21788__A1 _21649_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18653__B2 _18769_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16664__B1 _16391_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21518__A _21321_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19959_ _23554_/Q VGND VGND VPWR VPWR _22359_/B sky130_fd_sc_hd__inv_2
XANTENNA__20422__A _20409_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22970_ _23103_/A _22969_/X VGND VGND VPWR VPWR _22970_/X sky130_fd_sc_hd__and2_4
XFILLER_67_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16416__B1 _16236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21921_ _21926_/A _21921_/B VGND VGND VPWR VPWR _21922_/C sky130_fd_sc_hd__or2_4
XFILLER_56_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24872__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24640_ _24639_/CLK _24640_/D HRESETn VGND VGND VPWR VPWR _24640_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21852_ _12101_/Y _12086_/X _18381_/Y _12057_/X VGND VGND VPWR VPWR _21852_/X sky130_fd_sc_hd__o22a_4
XFILLER_70_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22316__A1_N _14096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24801__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23162__B1 _25394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20803_ _20800_/Y _20801_/Y _20802_/X VGND VGND VPWR VPWR _20803_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21253__A _21622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24571_ _24573_/CLK _16476_/X HRESETn VGND VGND VPWR VPWR _24571_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17450__B _13388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21783_ _21766_/X _21782_/X _22393_/A VGND VGND VPWR VPWR _21783_/Y sky130_fd_sc_hd__a21oi_4
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23522_ _23912_/CLK _20056_/X VGND VGND VPWR VPWR _13178_/B sky130_fd_sc_hd__dfxtp_4
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20734_ _20686_/A VGND VGND VPWR VPWR _20784_/A sky130_fd_sc_hd__inv_2
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23453_ _23452_/CLK _23453_/D VGND VGND VPWR VPWR _13360_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20665_ _17396_/B VGND VGND VPWR VPWR _20665_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19669__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22404_ _22132_/B VGND VGND VPWR VPWR _22821_/B sky130_fd_sc_hd__buf_2
X_23384_ _24413_/CLK _20411_/X VGND VGND VPWR VPWR _20407_/A sky130_fd_sc_hd__dfxtp_4
X_20596_ _23949_/Q _20593_/A _18885_/A VGND VGND VPWR VPWR _20596_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_192_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22084__A _22386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25123_ _23927_/CLK _25123_/D HRESETn VGND VGND VPWR VPWR _25123_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22335_ _21345_/Y _22320_/X _22322_/X _22326_/Y _22334_/X VGND VGND VPWR VPWR _22335_/X
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__25145__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16082__A _22816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25054_ _25052_/CLK _14828_/X HRESETn VGND VGND VPWR VPWR _14798_/C sky130_fd_sc_hd__dfrtp_4
X_22266_ _22266_/A _22229_/B VGND VGND VPWR VPWR _22266_/X sky130_fd_sc_hd__and2_4
XFILLER_191_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11716__B1 _11715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24005_ _24037_/CLK _20699_/Y HRESETn VGND VGND VPWR VPWR _13109_/A sky130_fd_sc_hd__dfrtp_4
X_21217_ _13779_/X _21214_/X _21216_/X _23348_/A _13780_/Y VGND VGND VPWR VPWR _21217_/X
+ sky130_fd_sc_hd__a32o_4
X_22197_ _22197_/A VGND VGND VPWR VPWR _22209_/A sky130_fd_sc_hd__buf_2
XFILLER_160_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22440__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21148_ _21151_/A _21147_/X VGND VGND VPWR VPWR _21148_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21428__A _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13970_ _13991_/A VGND VGND VPWR VPWR _14008_/A sky130_fd_sc_hd__buf_2
X_21079_ _11701_/X VGND VGND VPWR VPWR _22756_/B sky130_fd_sc_hd__buf_2
XFILLER_247_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16407__B1 _16320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12921_ _12920_/X VGND VGND VPWR VPWR _12921_/Y sky130_fd_sc_hd__inv_2
X_24907_ _24907_/CLK _15599_/X HRESETn VGND VGND VPWR VPWR _24907_/Q sky130_fd_sc_hd__dfrtp_4
X_15640_ _15640_/A _15640_/B _15640_/C _14422_/A VGND VGND VPWR VPWR _15644_/A sky130_fd_sc_hd__or4_4
XFILLER_246_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12852_ _12769_/Y _12857_/A _12851_/X VGND VGND VPWR VPWR _12852_/X sky130_fd_sc_hd__or3_4
X_24838_ _25344_/CLK _15808_/X HRESETn VGND VGND VPWR VPWR _24838_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24542__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11803_ _11803_/A VGND VGND VPWR VPWR _11803_/Y sky130_fd_sc_hd__inv_2
XPHY_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _21425_/A VGND VGND VPWR VPWR _12783_/Y sky130_fd_sc_hd__inv_2
X_15571_ _15569_/Y _15570_/X _11685_/X _15570_/X VGND VGND VPWR VPWR _15571_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _24766_/CLK _15945_/X HRESETn VGND VGND VPWR VPWR _22968_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_15_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17249_/C _17310_/B VGND VGND VPWR VPWR _17311_/C sky130_fd_sc_hd__or2_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ HWDATA[14] VGND VGND VPWR VPWR _16229_/A sky130_fd_sc_hd__buf_2
X_14522_ _23957_/Q _14521_/X _25114_/Q _14495_/Y VGND VGND VPWR VPWR _14522_/X sky130_fd_sc_hd__o22a_4
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18290_ _18280_/A _18289_/X _18280_/A _18289_/X VGND VGND VPWR VPWR _24217_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16900__A2_N _21059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17241_/A VGND VGND VPWR VPWR _17241_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _14180_/A _12043_/A VGND VGND VPWR VPWR _11668_/A sky130_fd_sc_hd__or2_4
X_14453_ _14452_/Y _14448_/X _14392_/X _14448_/X VGND VGND VPWR VPWR _14453_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22706__B _21843_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _13260_/A _13404_/B VGND VGND VPWR VPWR _13404_/X sky130_fd_sc_hd__or2_4
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _15472_/A VGND VGND VPWR VPWR _14384_/X sky130_fd_sc_hd__buf_2
X_17172_ _17171_/Y VGND VGND VPWR VPWR _17347_/C sky130_fd_sc_hd__buf_2
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13335_ _13431_/A _13335_/B VGND VGND VPWR VPWR _13335_/X sky130_fd_sc_hd__or2_4
X_16123_ _16084_/X VGND VGND VPWR VPWR _16124_/A sky130_fd_sc_hd__buf_2
XFILLER_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17088__A _17020_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13266_ _13443_/A _13266_/B VGND VGND VPWR VPWR _13266_/X sky130_fd_sc_hd__or2_4
X_16054_ _24723_/Q VGND VGND VPWR VPWR _16054_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25330__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12217_ _12217_/A VGND VGND VPWR VPWR _12217_/Y sky130_fd_sc_hd__inv_2
X_15005_ _24448_/Q VGND VGND VPWR VPWR _15005_/Y sky130_fd_sc_hd__inv_2
X_13197_ _13252_/A _23817_/Q VGND VGND VPWR VPWR _13201_/B sky130_fd_sc_hd__or2_4
X_19813_ _16863_/A VGND VGND VPWR VPWR _19813_/X sky130_fd_sc_hd__buf_2
XANTENNA__16646__B1 _16459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12148_ _14326_/A _14338_/A _12148_/C _25165_/Q VGND VGND VPWR VPWR _12149_/B sky130_fd_sc_hd__and4_4
XFILLER_111_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12171__A1_N _25439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19744_ _19742_/Y _19740_/X _19743_/X _19740_/X VGND VGND VPWR VPWR _19744_/X sky130_fd_sc_hd__a2bb2o_4
X_12079_ _12078_/Y _12072_/X _11793_/X _12060_/A VGND VGND VPWR VPWR _25479_/D sky130_fd_sc_hd__a2bb2o_4
X_16956_ _15980_/Y _17050_/A _15980_/Y _17050_/A VGND VGND VPWR VPWR _16956_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15907_ _15905_/X VGND VGND VPWR VPWR _15907_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19675_ _13223_/B VGND VGND VPWR VPWR _19675_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16887_ _16135_/Y _17747_/A _16135_/Y _17747_/A VGND VGND VPWR VPWR _16887_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18626_ _24522_/Q _24133_/Q _16603_/Y _18686_/A VGND VGND VPWR VPWR _18626_/X sky130_fd_sc_hd__o22a_4
X_15838_ _19646_/A VGND VGND VPWR VPWR _15838_/X sky130_fd_sc_hd__buf_2
XANTENNA__24283__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18557_ _18572_/A _18557_/B _18557_/C VGND VGND VPWR VPWR _24171_/D sky130_fd_sc_hd__and3_4
XFILLER_240_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15769_ HWDATA[0] VGND VGND VPWR VPWR _19646_/A sky130_fd_sc_hd__buf_2
XANTENNA__24212__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17508_ _25539_/Q _17507_/A _11713_/Y _17569_/A VGND VGND VPWR VPWR _17508_/X sky130_fd_sc_hd__o22a_4
XFILLER_205_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11789__A3 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18488_ _18580_/A VGND VGND VPWR VPWR _18823_/B sky130_fd_sc_hd__inv_2
XFILLER_33_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14188__A1 _14187_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _13797_/A VGND VGND VPWR VPWR _17440_/A sky130_fd_sc_hd__buf_2
XFILLER_220_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25489__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20450_ _20449_/X VGND VGND VPWR VPWR _20450_/X sky130_fd_sc_hd__buf_2
XANTENNA__25418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19109_ _19101_/A VGND VGND VPWR VPWR _19109_/X sky130_fd_sc_hd__buf_2
X_20381_ _20372_/X _20368_/X _14262_/A _23395_/Q _20370_/X VGND VGND VPWR VPWR _20381_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_118_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14415__A _14408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22120_ _15462_/Y _21365_/X _14217_/Y _14209_/X VGND VGND VPWR VPWR _22121_/A sky130_fd_sc_hd__o22a_4
XANTENNA__25071__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22958__B1 _12354_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22051_ _22582_/A VGND VGND VPWR VPWR _22051_/X sky130_fd_sc_hd__buf_2
XANTENNA__18626__A1 _24522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25000__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21002_ _21002_/A _21002_/B VGND VGND VPWR VPWR _21002_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_23_0_HCLK clkbuf_8_22_0_HCLK/A VGND VGND VPWR VPWR _24390_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_87_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11774__A _11774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_86_0_HCLK clkbuf_8_87_0_HCLK/A VGND VGND VPWR VPWR _25390_/CLK sky130_fd_sc_hd__clkbuf_1
X_22953_ _24600_/Q _23022_/B VGND VGND VPWR VPWR _22956_/B sky130_fd_sc_hd__or2_4
XFILLER_228_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13871__B1 _23442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21904_ _22219_/A _21902_/X _21903_/X VGND VGND VPWR VPWR _21904_/X sky130_fd_sc_hd__and3_4
XFILLER_28_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22884_ _23171_/A VGND VGND VPWR VPWR _22884_/X sky130_fd_sc_hd__buf_2
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21835_ _25248_/Q VGND VGND VPWR VPWR _21835_/Y sky130_fd_sc_hd__inv_2
X_24623_ _24623_/CLK _24623_/D HRESETn VGND VGND VPWR VPWR _24623_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12426__A1 _12248_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24554_ _24555_/CLK _24554_/D HRESETn VGND VGND VPWR VPWR _16517_/A sky130_fd_sc_hd__dfrtp_4
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21766_ _21901_/A _21758_/X _21765_/X VGND VGND VPWR VPWR _21766_/X sky130_fd_sc_hd__or3_4
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21161__A2 _14209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22807__A _22807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20717_ _13117_/A _13117_/B VGND VGND VPWR VPWR _20718_/A sky130_fd_sc_hd__or2_4
X_23505_ _23497_/CLK _23505_/D VGND VGND VPWR VPWR _23505_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24485_ _24486_/CLK _24485_/D HRESETn VGND VGND VPWR VPWR _16701_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21697_ _21548_/X _21601_/X _21697_/C _21697_/D VGND VGND VPWR VPWR HRDATA[2] sky130_fd_sc_hd__or4_4
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23436_ _24317_/CLK _20280_/X VGND VGND VPWR VPWR _20278_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12729__A2 _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20648_ _23982_/Q _20645_/A VGND VGND VPWR VPWR _20648_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__25159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23367_ _21014_/X VGND VGND VPWR VPWR IRQ[23] sky130_fd_sc_hd__buf_2
X_20579_ _20578_/X VGND VGND VPWR VPWR _23944_/D sky130_fd_sc_hd__inv_2
XANTENNA__18865__B2 _18658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13120_ _13120_/A _13120_/B VGND VGND VPWR VPWR _13121_/B sky130_fd_sc_hd__or2_4
X_22318_ _22317_/Y _21349_/A _14394_/Y _21351_/X VGND VGND VPWR VPWR _22319_/A sky130_fd_sc_hd__o22a_4
X_25106_ _25117_/CLK _25106_/D HRESETn VGND VGND VPWR VPWR _21847_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_124_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23298_ _16456_/A _23172_/X _23133_/X VGND VGND VPWR VPWR _23298_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15019__A1_N _25013_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13051_ _12291_/X _13051_/B VGND VGND VPWR VPWR _13051_/Y sky130_fd_sc_hd__nand2_4
X_25037_ _25015_/CLK _15176_/X HRESETn VGND VGND VPWR VPWR _25037_/Q sky130_fd_sc_hd__dfrtp_4
X_22249_ _18296_/A _22245_/X _22249_/C VGND VGND VPWR VPWR _22249_/X sky130_fd_sc_hd__or3_4
XANTENNA__16540__A _16792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12002_ _12002_/A VGND VGND VPWR VPWR _12002_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24794__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16810_ _16810_/A VGND VGND VPWR VPWR _16810_/Y sky130_fd_sc_hd__inv_2
X_17790_ _17790_/A _17790_/B _17790_/C VGND VGND VPWR VPWR _17790_/X sky130_fd_sc_hd__and3_4
XANTENNA__24723__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16741_ _24469_/Q VGND VGND VPWR VPWR _16741_/Y sky130_fd_sc_hd__inv_2
X_13953_ _13953_/A _14236_/D _13939_/X _15424_/C VGND VGND VPWR VPWR _14234_/A sky130_fd_sc_hd__or4_4
XFILLER_247_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19570__B _21159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12904_ _12838_/B _12907_/A VGND VGND VPWR VPWR _12904_/X sky130_fd_sc_hd__or2_4
X_19460_ _19460_/A VGND VGND VPWR VPWR _22235_/B sky130_fd_sc_hd__inv_2
X_16672_ _24497_/Q VGND VGND VPWR VPWR _16672_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13884_ _13916_/C VGND VGND VPWR VPWR _13903_/A sky130_fd_sc_hd__buf_2
XFILLER_62_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18411_ _18411_/A VGND VGND VPWR VPWR _18462_/B sky130_fd_sc_hd__inv_2
XANTENNA__16800__B1 _16459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15623_ _14407_/A VGND VGND VPWR VPWR _15623_/X sky130_fd_sc_hd__buf_2
XFILLER_222_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12835_ _12762_/Y _12948_/A _12835_/C _12834_/X VGND VGND VPWR VPWR _12835_/X sky130_fd_sc_hd__or4_4
X_19391_ _17986_/B VGND VGND VPWR VPWR _19391_/Y sky130_fd_sc_hd__inv_2
X_18342_ _18342_/A _18341_/Y VGND VGND VPWR VPWR _18342_/X sky130_fd_sc_hd__or2_4
X_15554_ HWDATA[30] VGND VGND VPWR VPWR _15554_/X sky130_fd_sc_hd__buf_2
X_12766_ _12766_/A VGND VGND VPWR VPWR _12766_/Y sky130_fd_sc_hd__inv_2
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22717__A _22704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _20601_/A _14500_/X _25108_/Q _14502_/X VGND VGND VPWR VPWR _14505_/X sky130_fd_sc_hd__o22a_4
X_11717_ _11717_/A VGND VGND VPWR VPWR _11717_/Y sky130_fd_sc_hd__inv_2
X_18273_ _21281_/B VGND VGND VPWR VPWR _18274_/A sky130_fd_sc_hd__buf_2
XFILLER_202_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12697_/A _12697_/B VGND VGND VPWR VPWR _12701_/B sky130_fd_sc_hd__or2_4
X_15485_ _15511_/A VGND VGND VPWR VPWR _15489_/A sky130_fd_sc_hd__buf_2
XFILLER_202_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20360__B1 _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17224_ _24640_/Q _17215_/Y _16348_/Y _21856_/A VGND VGND VPWR VPWR _17224_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14436_ _14435_/Y _14431_/X _14392_/X _14431_/X VGND VGND VPWR VPWR _14436_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25511__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17155_ _17153_/Y _17154_/X _17148_/C VGND VGND VPWR VPWR _24376_/D sky130_fd_sc_hd__and3_4
X_14367_ _14366_/X VGND VGND VPWR VPWR _14425_/B sky130_fd_sc_hd__buf_2
XANTENNA__17249__C _17249_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16106_ _23049_/A VGND VGND VPWR VPWR _16106_/Y sky130_fd_sc_hd__inv_2
X_13318_ _13314_/X _13318_/B _13318_/C VGND VGND VPWR VPWR _13319_/C sky130_fd_sc_hd__and3_4
X_14298_ _14295_/X _14297_/Y _25324_/Q _14295_/X VGND VGND VPWR VPWR _25178_/D sky130_fd_sc_hd__a2bb2o_4
X_17086_ _17085_/X VGND VGND VPWR VPWR _17086_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22452__A _23075_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16037_ _24730_/Q VGND VGND VPWR VPWR _16037_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13249_ _13249_/A VGND VGND VPWR VPWR _13389_/A sky130_fd_sc_hd__buf_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18608__B2 _24142_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16450__A _24578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17988_ _17987_/X _19416_/A VGND VGND VPWR VPWR _17988_/X sky130_fd_sc_hd__or2_4
XANTENNA__22168__A1 _14428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24464__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12105__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22168__B2 _21368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19727_ _19727_/A VGND VGND VPWR VPWR _19727_/Y sky130_fd_sc_hd__inv_2
X_16939_ _16098_/Y _24284_/Q _24701_/Q _16938_/Y VGND VGND VPWR VPWR _16942_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19658_ _19656_/Y _19651_/X _19633_/X _19657_/X VGND VGND VPWR VPWR _23664_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23117__B1 _12878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18609_ _24136_/Q VGND VGND VPWR VPWR _18610_/A sky130_fd_sc_hd__inv_2
XFILLER_65_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19589_ _23685_/Q VGND VGND VPWR VPWR _19589_/Y sky130_fd_sc_hd__inv_2
XFILLER_241_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21620_ _21616_/X _21619_/X _14744_/X VGND VGND VPWR VPWR _21620_/X sky130_fd_sc_hd__o21a_4
XANTENNA__13314__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21531__A _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21551_ _25104_/Q _22119_/B VGND VGND VPWR VPWR _21551_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15358__B1 _15334_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20351__B1 _19600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20502_ _14266_/Y _20502_/B _20524_/B VGND VGND VPWR VPWR _20504_/A sky130_fd_sc_hd__and3_4
XFILLER_21_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24270_ _24686_/CLK _17847_/Y HRESETn VGND VGND VPWR VPWR _24270_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21482_ _21677_/A _21482_/B VGND VGND VPWR VPWR _21483_/C sky130_fd_sc_hd__or2_4
XANTENNA__25252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23221_ _23280_/A _23221_/B VGND VGND VPWR VPWR _23228_/C sky130_fd_sc_hd__and2_4
X_20433_ _25152_/Q _23926_/D _20455_/C VGND VGND VPWR VPWR _20466_/B sky130_fd_sc_hd__o21a_4
XFILLER_147_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11769__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23152_ _21232_/X VGND VGND VPWR VPWR _23152_/X sky130_fd_sc_hd__buf_2
XFILLER_162_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16994__A1_N _16037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20364_ _23403_/Q VGND VGND VPWR VPWR _21480_/B sky130_fd_sc_hd__inv_2
X_22103_ _14430_/Y _21365_/A _14447_/Y _17411_/X VGND VGND VPWR VPWR _22104_/A sky130_fd_sc_hd__o22a_4
XFILLER_162_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23083_ _12194_/Y _23268_/A _23082_/X VGND VGND VPWR VPWR _23083_/Y sky130_fd_sc_hd__o21ai_4
X_20295_ _23430_/Q VGND VGND VPWR VPWR _21941_/B sky130_fd_sc_hd__inv_2
XFILLER_88_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22034_ _22020_/A _22034_/B VGND VGND VPWR VPWR _22034_/X sky130_fd_sc_hd__or2_4
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24134__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23985_ _23986_/CLK _20663_/Y HRESETn VGND VGND VPWR VPWR _17394_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15704__A _15704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22936_ _23005_/A _22933_/X _22936_/C VGND VGND VPWR VPWR _22937_/D sky130_fd_sc_hd__and3_4
XANTENNA__21425__B _22420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15597__B1 _11730_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22867_ _22866_/X VGND VGND VPWR VPWR _22867_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21831__A2_N _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12620_ _12620_/A VGND VGND VPWR VPWR _12620_/Y sky130_fd_sc_hd__inv_2
X_24606_ _24520_/CLK _24606_/D HRESETn VGND VGND VPWR VPWR _24606_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21818_ _21803_/A _21816_/X _21818_/C VGND VGND VPWR VPWR _21818_/X sky130_fd_sc_hd__and3_4
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22798_ _22798_/A VGND VGND VPWR VPWR _23128_/A sky130_fd_sc_hd__inv_2
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12551_ _12551_/A VGND VGND VPWR VPWR _12551_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21749_ _20838_/Y _21597_/X _13113_/A _21598_/X VGND VGND VPWR VPWR _21749_/X sky130_fd_sc_hd__a2bb2o_4
X_24537_ _24539_/CLK _24537_/D HRESETn VGND VGND VPWR VPWR _16564_/A sky130_fd_sc_hd__dfrtp_4
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20342__B1 _19617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _12217_/A _12482_/B VGND VGND VPWR VPWR _12483_/C sky130_fd_sc_hd__or2_4
X_15270_ _15244_/A _15244_/B _15185_/A _15268_/B VGND VGND VPWR VPWR _15271_/A sky130_fd_sc_hd__a211o_4
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24468_ _24460_/CLK _16744_/X HRESETn VGND VGND VPWR VPWR _16743_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ _14220_/Y _14218_/X _13785_/X _14218_/X VGND VGND VPWR VPWR _14221_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_200_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23419_ _23425_/CLK _23419_/D VGND VGND VPWR VPWR _23419_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24399_ _24390_/CLK _17073_/Y HRESETn VGND VGND VPWR VPWR _17023_/A sky130_fd_sc_hd__dfrtp_4
X_14152_ _14118_/X _14151_/X _14433_/A _14115_/X VGND VGND VPWR VPWR _14152_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__23368__A _23368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24975__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25201__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13103_ _13095_/B _13102_/X _13091_/C VGND VGND VPWR VPWR _25336_/D sky130_fd_sc_hd__and3_4
X_14083_ _14083_/A VGND VGND VPWR VPWR _14096_/A sky130_fd_sc_hd__inv_2
X_18960_ _14654_/A VGND VGND VPWR VPWR _18960_/X sky130_fd_sc_hd__buf_2
XANTENNA__17366__A _17366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24904__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13034_ _13033_/X VGND VGND VPWR VPWR _13035_/B sky130_fd_sc_hd__inv_2
X_17911_ _17898_/Y _17908_/A _17910_/X _21991_/A _17908_/Y VGND VGND VPWR VPWR _24255_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_98_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18891_ _18871_/X _18885_/X _23954_/Q _20984_/B _18888_/X VGND VGND VPWR VPWR _24122_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_239_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17842_ _17842_/A VGND VGND VPWR VPWR _17843_/B sky130_fd_sc_hd__inv_2
XFILLER_79_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17773_ _16950_/X _17602_/B VGND VGND VPWR VPWR _17773_/X sky130_fd_sc_hd__and2_4
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14985_ _25009_/Q VGND VGND VPWR VPWR _15272_/A sky130_fd_sc_hd__inv_2
X_19512_ _23710_/Q VGND VGND VPWR VPWR _21814_/B sky130_fd_sc_hd__inv_2
X_16724_ _16724_/A _16792_/B VGND VGND VPWR VPWR _16725_/A sky130_fd_sc_hd__nor2_4
X_13936_ _15421_/B _13935_/X VGND VGND VPWR VPWR _13936_/Y sky130_fd_sc_hd__nor2_4
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19443_ _19442_/Y _19440_/X _19351_/X _19440_/X VGND VGND VPWR VPWR _23735_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16655_ _16655_/A VGND VGND VPWR VPWR _16655_/X sky130_fd_sc_hd__buf_2
X_13867_ _21559_/A _13849_/X _25245_/Q _13844_/X VGND VGND VPWR VPWR _13867_/X sky130_fd_sc_hd__o22a_4
XFILLER_223_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17251__D _17314_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15606_ _15605_/Y _15601_/X _11748_/X _15601_/X VGND VGND VPWR VPWR _15606_/X sky130_fd_sc_hd__a2bb2o_4
X_12818_ _12818_/A VGND VGND VPWR VPWR _12845_/C sky130_fd_sc_hd__inv_2
X_19374_ _23759_/Q VGND VGND VPWR VPWR _19374_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16586_ _16584_/Y _16580_/X _16229_/X _16585_/X VGND VGND VPWR VPWR _24529_/D sky130_fd_sc_hd__a2bb2o_4
X_13798_ _16361_/A VGND VGND VPWR VPWR _13798_/X sky130_fd_sc_hd__buf_2
XANTENNA__14260__B1 _13791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18325_ _17460_/A VGND VGND VPWR VPWR _20220_/D sky130_fd_sc_hd__buf_2
XFILLER_231_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21351__A _14209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15537_ _13581_/B VGND VGND VPWR VPWR _15537_/Y sky130_fd_sc_hd__inv_2
X_12749_ _21027_/A VGND VGND VPWR VPWR _12749_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18256_ _18240_/A VGND VGND VPWR VPWR _18256_/X sky130_fd_sc_hd__buf_2
X_15468_ _15468_/A VGND VGND VPWR VPWR _15468_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17207_ _16324_/Y _22709_/A _16324_/Y _22709_/A VGND VGND VPWR VPWR _17208_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14419_ _25138_/Q VGND VGND VPWR VPWR _14419_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22086__B1 _21627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18187_ _18056_/A _18185_/X _18186_/X VGND VGND VPWR VPWR _18187_/X sky130_fd_sc_hd__and3_4
XANTENNA__15760__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15399_ _15294_/C _15386_/X VGND VGND VPWR VPWR _15399_/Y sky130_fd_sc_hd__nand2_4
X_17138_ _17142_/A _17131_/X _17138_/C VGND VGND VPWR VPWR _17138_/X sky130_fd_sc_hd__and3_4
XANTENNA__17501__B2 _25546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17069_ _16965_/Y _17069_/B VGND VGND VPWR VPWR _17070_/C sky130_fd_sc_hd__or2_4
XFILLER_143_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16180__A _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24645__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20080_ _21637_/B _20079_/X _19824_/X _20079_/X VGND VGND VPWR VPWR _23509_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22910__A _23171_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23338__B1 _23326_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15524__A _15530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23770_ _24088_/CLK _19344_/X VGND VGND VPWR VPWR _17948_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_238_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20982_ _24121_/Q _20982_/B VGND VGND VPWR VPWR _20982_/X sky130_fd_sc_hd__and2_4
XFILLER_226_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22721_ _22721_/A VGND VGND VPWR VPWR _23094_/A sky130_fd_sc_hd__buf_2
XANTENNA__15579__B1 _11695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22652_ _16539_/A _22651_/X _22138_/C _16040_/A _15983_/X VGND VGND VPWR VPWR _22652_/X
+ sky130_fd_sc_hd__a32o_4
X_25440_ _24753_/CLK _12478_/X HRESETn VGND VGND VPWR VPWR _12197_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_81_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22357__A _21463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21603_ _22056_/A VGND VGND VPWR VPWR _22221_/A sky130_fd_sc_hd__buf_2
XFILLER_80_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21261__A _22069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22583_ _13531_/Y _22619_/B VGND VGND VPWR VPWR _22583_/X sky130_fd_sc_hd__and2_4
X_25371_ _25375_/CLK _12961_/X HRESETn VGND VGND VPWR VPWR _25371_/Q sky130_fd_sc_hd__dfrtp_4
X_21534_ _21534_/A _23172_/A VGND VGND VPWR VPWR _21534_/X sky130_fd_sc_hd__or2_4
X_24322_ _24317_/CLK _24322_/D HRESETn VGND VGND VPWR VPWR _17491_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24253_ _24252_/CLK _24253_/D HRESETn VGND VGND VPWR VPWR _17914_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21465_ _21920_/A VGND VGND VPWR VPWR _21466_/A sky130_fd_sc_hd__buf_2
XANTENNA__15751__B1 _13818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23204_ _24030_/Q _21292_/X _13635_/A _21315_/X VGND VGND VPWR VPWR _23204_/Y sky130_fd_sc_hd__a22oi_4
X_20416_ _22070_/B _20410_/X _16863_/A _20415_/X VGND VGND VPWR VPWR _23382_/D sky130_fd_sc_hd__a2bb2o_4
X_24184_ _24675_/CLK _18509_/Y HRESETn VGND VGND VPWR VPWR _18459_/A sky130_fd_sc_hd__dfrtp_4
X_21396_ _22197_/A _21396_/B VGND VGND VPWR VPWR _21396_/X sky130_fd_sc_hd__or2_4
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23135_ _16557_/A _22884_/X _22928_/X _23134_/X VGND VGND VPWR VPWR _23135_/X sky130_fd_sc_hd__a211o_4
X_20347_ _23409_/Q VGND VGND VPWR VPWR _22357_/B sky130_fd_sc_hd__inv_2
XANTENNA__23026__C1 _23025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24386__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23066_ _24538_/Q _22884_/X _22928_/X _23065_/X VGND VGND VPWR VPWR _23066_/X sky130_fd_sc_hd__a211o_4
X_20278_ _20278_/A VGND VGND VPWR VPWR _21655_/B sky130_fd_sc_hd__inv_2
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24315__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14322__B _18372_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22017_ _22021_/A _22017_/B _22017_/C VGND VGND VPWR VPWR _22017_/X sky130_fd_sc_hd__and3_4
XANTENNA__21052__A1 _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13219__A _13422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_56_0_HCLK clkbuf_7_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14770_ _16165_/B _14768_/A _25060_/Q _14769_/X VGND VGND VPWR VPWR _14770_/X sky130_fd_sc_hd__o22a_4
X_11982_ _24095_/Q _11979_/X _11981_/Y VGND VGND VPWR VPWR _11983_/B sky130_fd_sc_hd__o21a_4
X_23968_ _25243_/CLK _21009_/X HRESETn VGND VGND VPWR VPWR _23968_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13721_ _25280_/Q VGND VGND VPWR VPWR _13721_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11681__B _11681_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22919_ _21319_/X VGND VGND VPWR VPWR _22919_/X sky130_fd_sc_hd__buf_2
XFILLER_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23899_ _25171_/CLK _23899_/D VGND VGND VPWR VPWR _18210_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__23950__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16440_ _24579_/Q VGND VGND VPWR VPWR _18560_/A sky130_fd_sc_hd__inv_2
XFILLER_44_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13652_ _13651_/X VGND VGND VPWR VPWR _20932_/B sky130_fd_sc_hd__buf_2
XFILLER_71_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12603_ _12724_/A VGND VGND VPWR VPWR _12716_/A sky130_fd_sc_hd__inv_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21171__A _15331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16371_ _16363_/Y _16370_/X _15991_/X _16370_/X VGND VGND VPWR VPWR _16371_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13583_ _12083_/A _13800_/B _11668_/A _13765_/A VGND VGND VPWR VPWR _14422_/A sky130_fd_sc_hd__or4_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18110_ _17985_/X _18110_/B VGND VGND VPWR VPWR _18110_/X sky130_fd_sc_hd__or2_4
X_15322_ _15322_/A VGND VGND VPWR VPWR _25004_/D sky130_fd_sc_hd__inv_2
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _24884_/Q VGND VGND VPWR VPWR _12534_/Y sky130_fd_sc_hd__inv_2
X_19090_ _23859_/Q VGND VGND VPWR VPWR _21250_/B sky130_fd_sc_hd__inv_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18041_ _17990_/X _18039_/X _18041_/C VGND VGND VPWR VPWR _18042_/C sky130_fd_sc_hd__and3_4
XFILLER_157_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15253_ _15253_/A VGND VGND VPWR VPWR _25018_/D sky130_fd_sc_hd__inv_2
X_12465_ _12208_/X _12191_/X _12459_/X VGND VGND VPWR VPWR _12465_/X sky130_fd_sc_hd__or3_4
XANTENNA__15742__B1 _24869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14204_ _14203_/Y _14199_/X _13798_/X _14190_/A VGND VGND VPWR VPWR _25203_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_184_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12396_ _12279_/A _12396_/B VGND VGND VPWR VPWR _12396_/X sky130_fd_sc_hd__or2_4
X_15184_ _15065_/X _15167_/B _15066_/A VGND VGND VPWR VPWR _15184_/X sky130_fd_sc_hd__o21a_4
XFILLER_126_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14135_ _14115_/X VGND VGND VPWR VPWR _14135_/X sky130_fd_sc_hd__buf_2
X_19992_ _22344_/B _19991_/X _19964_/X _19991_/X VGND VGND VPWR VPWR _19992_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14066_ _13987_/X _14054_/X _14046_/X _13986_/X _14065_/X VGND VGND VPWR VPWR _14066_/X
+ sky130_fd_sc_hd__a32o_4
X_18943_ _18941_/Y _18939_/X _18942_/X _18939_/X VGND VGND VPWR VPWR _18943_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22730__A _22730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24056__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13017_ _13017_/A _13016_/X VGND VGND VPWR VPWR _13017_/X sky130_fd_sc_hd__or2_4
X_18874_ _20558_/A _20553_/A VGND VGND VPWR VPWR _18874_/X sky130_fd_sc_hd__or2_4
XANTENNA__12033__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17825_ _16921_/Y _17828_/A VGND VGND VPWR VPWR _17826_/B sky130_fd_sc_hd__or2_4
XFILLER_121_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16839__A1_N _14911_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21346__A _21346_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17756_ _24270_/Q VGND VGND VPWR VPWR _17756_/Y sky130_fd_sc_hd__inv_2
X_14968_ _25030_/Q _14966_/Y _15207_/A _14964_/A VGND VGND VPWR VPWR _14968_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16707_ _16706_/Y _16704_/X _16349_/X _16704_/X VGND VGND VPWR VPWR _24483_/D sky130_fd_sc_hd__a2bb2o_4
X_13919_ _13911_/Y _13912_/X _13915_/X _13923_/D VGND VGND VPWR VPWR _13920_/A sky130_fd_sc_hd__or4_4
X_17687_ _17530_/A _17687_/B VGND VGND VPWR VPWR _17688_/B sky130_fd_sc_hd__or2_4
XANTENNA__20554__B1 _20600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14899_ _24435_/Q VGND VGND VPWR VPWR _14899_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19426_ _19426_/A VGND VGND VPWR VPWR _19426_/X sky130_fd_sc_hd__buf_2
XFILLER_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16638_ _15818_/X _15639_/Y _15702_/X _23323_/A _16640_/A VGND VGND VPWR VPWR _16638_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_223_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21081__A _21080_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19357_ _11785_/A VGND VGND VPWR VPWR _19357_/X sky130_fd_sc_hd__buf_2
X_16569_ _16569_/A VGND VGND VPWR VPWR _16569_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18308_ _24212_/Q VGND VGND VPWR VPWR _21189_/A sky130_fd_sc_hd__inv_2
XANTENNA__12795__B1 _22667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19288_ _19287_/Y _19283_/X _19221_/X _19283_/X VGND VGND VPWR VPWR _23790_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24897__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18239_ _20369_/A VGND VGND VPWR VPWR _18240_/A sky130_fd_sc_hd__inv_2
XFILLER_175_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15733__B1 _11718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24826__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21250_ _21250_/A _21250_/B VGND VGND VPWR VPWR _21251_/C sky130_fd_sc_hd__or2_4
XFILLER_191_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20201_ _20200_/Y VGND VGND VPWR VPWR _20201_/X sky130_fd_sc_hd__buf_2
XANTENNA__17486__B1 _13150_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21181_ _24213_/Q _21181_/B _21181_/C VGND VGND VPWR VPWR _21181_/X sky130_fd_sc_hd__and3_4
XANTENNA__15519__A _15530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14423__A _21365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20132_ _23491_/Q VGND VGND VPWR VPWR _21269_/B sky130_fd_sc_hd__inv_2
XFILLER_171_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20063_ _20054_/A _18328_/A _14262_/A _13399_/B _20055_/A VGND VGND VPWR VPWR _23516_/D
+ sky130_fd_sc_hd__a32o_4
X_24940_ _25510_/CLK _15504_/X HRESETn VGND VGND VPWR VPWR _24940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_225_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21585__A2 _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22782__B2 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21256__A _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24871_ _24866_/CLK _15737_/X HRESETn VGND VGND VPWR VPWR _24871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12878__A _12878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23822_ _23831_/CLK _19197_/X VGND VGND VPWR VPWR _23822_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20965_ _11992_/A _20964_/B VGND VGND VPWR VPWR _20965_/X sky130_fd_sc_hd__and2_4
X_23753_ _23785_/CLK _23753_/D VGND VGND VPWR VPWR _17986_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__20545__B1 _20600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22704_ _23091_/A _22701_/X _22704_/C VGND VGND VPWR VPWR _22704_/X sky130_fd_sc_hd__and3_4
XFILLER_199_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20896_ _20923_/A VGND VGND VPWR VPWR _20896_/X sky130_fd_sc_hd__buf_2
X_23684_ _23706_/CLK _19593_/X VGND VGND VPWR VPWR _19592_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25423_ _24872_/CLK _12651_/Y HRESETn VGND VGND VPWR VPWR _12567_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_201_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22635_ _24624_/Q _21337_/X VGND VGND VPWR VPWR _22635_/X sky130_fd_sc_hd__or2_4
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22566_ _22566_/A _22756_/B VGND VGND VPWR VPWR _22566_/X sky130_fd_sc_hd__and2_4
X_25354_ _25344_/CLK _25354_/D HRESETn VGND VGND VPWR VPWR _25354_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21517_ _21502_/Y _21514_/Y _22041_/A VGND VGND VPWR VPWR _21518_/D sky130_fd_sc_hd__o21a_4
X_24305_ _24305_/CLK _24305_/D HRESETn VGND VGND VPWR VPWR _17568_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23247__C1 _23246_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22497_ _22485_/X _22492_/Y _22493_/X _22496_/X VGND VGND VPWR VPWR _22497_/X sky130_fd_sc_hd__a2bb2o_4
X_25285_ _25285_/CLK _25285_/D HRESETn VGND VGND VPWR VPWR _11803_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24567__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12250_ _12241_/X _12244_/X _12246_/X _12249_/X VGND VGND VPWR VPWR _12250_/X sky130_fd_sc_hd__or4_4
X_21448_ _15780_/B VGND VGND VPWR VPWR _21448_/X sky130_fd_sc_hd__buf_2
X_24236_ _24236_/CLK _24236_/D HRESETn VGND VGND VPWR VPWR _24236_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_182_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12181_ _22968_/A VGND VGND VPWR VPWR _12181_/Y sky130_fd_sc_hd__inv_2
X_24167_ _24650_/CLK _18574_/X HRESETn VGND VGND VPWR VPWR _24167_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21379_ _13794_/Y _21379_/B VGND VGND VPWR VPWR _21379_/X sky130_fd_sc_hd__and2_4
XFILLER_107_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17347__C _17347_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23118_ _23118_/A _23117_/X _22919_/X VGND VGND VPWR VPWR _23118_/X sky130_fd_sc_hd__or3_4
XFILLER_162_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24098_ _25492_/CLK _12012_/C HRESETn VGND VGND VPWR VPWR _24098_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15940_ _12195_/Y _15935_/X _15939_/X _15935_/X VGND VGND VPWR VPWR _15940_/X sky130_fd_sc_hd__a2bb2o_4
X_23049_ _23049_/A _22909_/B VGND VGND VPWR VPWR _23049_/X sky130_fd_sc_hd__or2_4
XFILLER_135_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20379__A3 _18257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21166__A _18560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15871_ _12812_/Y _15865_/X _11695_/X _15865_/X VGND VGND VPWR VPWR _24807_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17610_ _17620_/A _17608_/X _17610_/C VGND VGND VPWR VPWR _24318_/D sky130_fd_sc_hd__and3_4
X_14822_ _25055_/Q _14798_/X _14814_/C _14799_/Y VGND VGND VPWR VPWR _14822_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23317__A3 _22135_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18590_ _18589_/A _18593_/A VGND VGND VPWR VPWR _18591_/B sky130_fd_sc_hd__or2_4
XANTENNA__25355__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17541_ _17541_/A VGND VGND VPWR VPWR _17541_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14753_ _22225_/A VGND VGND VPWR VPWR _14753_/X sky130_fd_sc_hd__buf_2
X_11965_ _11934_/B _11956_/X _11964_/Y VGND VGND VPWR VPWR _11965_/X sky130_fd_sc_hd__a21o_4
XFILLER_245_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13704_ _13676_/B _13694_/X _13703_/Y _13701_/X _11832_/A VGND VGND VPWR VPWR _13704_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_8_143_0_HCLK clkbuf_7_71_0_HCLK/X VGND VGND VPWR VPWR _25171_/CLK sky130_fd_sc_hd__clkbuf_1
X_17472_ _17443_/X _18326_/B _17472_/C _17472_/D VGND VGND VPWR VPWR _17472_/X sky130_fd_sc_hd__or4_4
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14684_ _13745_/X _14683_/X VGND VGND VPWR VPWR _14684_/X sky130_fd_sc_hd__and2_4
X_11896_ _11802_/Y _11896_/B VGND VGND VPWR VPWR _11897_/A sky130_fd_sc_hd__and2_4
XFILLER_72_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19211_ _19224_/A VGND VGND VPWR VPWR _19211_/X sky130_fd_sc_hd__buf_2
X_16423_ _15107_/Y _16418_/X _16141_/X _16422_/X VGND VGND VPWR VPWR _16423_/X sky130_fd_sc_hd__a2bb2o_4
X_13635_ _13635_/A _20941_/A VGND VGND VPWR VPWR _13635_/X sky130_fd_sc_hd__or2_4
XFILLER_44_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15963__B1 _22597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19154__B1 _19106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19142_ _19141_/X VGND VGND VPWR VPWR _19149_/A sky130_fd_sc_hd__inv_2
XANTENNA__13412__A _13254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16354_ _16352_/Y _16350_/X _16353_/X _16350_/X VGND VGND VPWR VPWR _16354_/X sky130_fd_sc_hd__a2bb2o_4
X_13566_ _13566_/A VGND VGND VPWR VPWR _14557_/A sky130_fd_sc_hd__inv_2
XANTENNA__24990__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15305_ _15150_/Y _15323_/A _15304_/X VGND VGND VPWR VPWR _15308_/B sky130_fd_sc_hd__or3_4
XFILLER_8_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12517_ _25401_/Q VGND VGND VPWR VPWR _12689_/A sky130_fd_sc_hd__inv_2
X_19073_ _19073_/A VGND VGND VPWR VPWR _19074_/A sky130_fd_sc_hd__inv_2
X_16285_ _16284_/X VGND VGND VPWR VPWR _16285_/X sky130_fd_sc_hd__buf_2
XANTENNA__15715__B1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13497_ _13496_/Y _13494_/X _11781_/X _13494_/X VGND VGND VPWR VPWR _25310_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16723__A _24477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18024_ _18024_/A VGND VGND VPWR VPWR _18024_/X sky130_fd_sc_hd__buf_2
X_15236_ _25021_/Q _15236_/B VGND VGND VPWR VPWR _15236_/X sky130_fd_sc_hd__or2_4
X_12448_ _12418_/B _12447_/X VGND VGND VPWR VPWR _12448_/X sky130_fd_sc_hd__or2_4
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24237__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_11_0_HCLK_A clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15167_ _15160_/A _15167_/B VGND VGND VPWR VPWR _15168_/C sky130_fd_sc_hd__or2_4
X_12379_ _12379_/A _12378_/X VGND VGND VPWR VPWR _12379_/X sky130_fd_sc_hd__or2_4
XANTENNA__14243__A _14243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14118_ _14099_/A VGND VGND VPWR VPWR _14118_/X sky130_fd_sc_hd__buf_2
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15098_ _25000_/Q _24604_/Q _15333_/A _15097_/Y VGND VGND VPWR VPWR _15102_/C sky130_fd_sc_hd__o22a_4
X_19975_ _21944_/B _19971_/X _19974_/X _19971_/X VGND VGND VPWR VPWR _19975_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14049_ _14049_/A _14049_/B VGND VGND VPWR VPWR _14049_/X sky130_fd_sc_hd__or2_4
X_18926_ _18924_/Y _18925_/X _16849_/X _18925_/X VGND VGND VPWR VPWR _18926_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23275__B _22658_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22764__B2 _22763_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18857_ _16520_/A _18788_/B _16507_/Y _18791_/A VGND VGND VPWR VPWR _18861_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17640__B1 _17593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17808_ _17791_/A _17804_/Y _17807_/X VGND VGND VPWR VPWR _17808_/X sky130_fd_sc_hd__or3_4
X_18788_ _18686_/A _18788_/B _18804_/A _18810_/A VGND VGND VPWR VPWR _18797_/B sky130_fd_sc_hd__or4_4
XANTENNA__25096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17739_ _17703_/X _17706_/X _17737_/Y _17704_/C _17738_/X VGND VGND VPWR VPWR _24290_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25025__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19393__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20750_ _13121_/D _20749_/A VGND VGND VPWR VPWR _20750_/X sky130_fd_sc_hd__or2_4
XFILLER_63_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14206__B1 _13788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19409_ _19407_/Y _19403_/X _19408_/X _19388_/Y VGND VGND VPWR VPWR _19409_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20681_ _20491_/X _20498_/X _20613_/B VGND VGND VPWR VPWR _23996_/D sky130_fd_sc_hd__o21a_4
XFILLER_149_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15954__B1 _15953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19145__B1 _19144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22420_ _22420_/A _22420_/B VGND VGND VPWR VPWR _22420_/X sky130_fd_sc_hd__or2_4
XANTENNA__12768__B1 _12766_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22351_ _22020_/A _22351_/B VGND VGND VPWR VPWR _22351_/X sky130_fd_sc_hd__or2_4
XFILLER_176_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24660__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21302_ _22829_/A VGND VGND VPWR VPWR _21303_/A sky130_fd_sc_hd__inv_2
X_25070_ _25070_/CLK _14703_/Y HRESETn VGND VGND VPWR VPWR _25070_/Q sky130_fd_sc_hd__dfstp_4
X_22282_ _22282_/A VGND VGND VPWR VPWR _22282_/X sky130_fd_sc_hd__buf_2
XFILLER_156_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24021_ _24051_/CLK _20770_/X HRESETn VGND VGND VPWR VPWR _20767_/A sky130_fd_sc_hd__dfrtp_4
X_21233_ _25299_/Q _21128_/B VGND VGND VPWR VPWR _21233_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__11777__A _25523_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15249__A _15249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21164_ _17435_/Y _21132_/Y _14179_/B _21163_/X VGND VGND VPWR VPWR _21175_/A sky130_fd_sc_hd__a211o_4
XFILLER_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20115_ _20115_/A VGND VGND VPWR VPWR _20116_/A sky130_fd_sc_hd__inv_2
XFILLER_104_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21095_ _21040_/X _21092_/X _21864_/C _21094_/X VGND VGND VPWR VPWR _21096_/C sky130_fd_sc_hd__a211o_4
XFILLER_86_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20046_ _20034_/A VGND VGND VPWR VPWR _20046_/X sky130_fd_sc_hd__buf_2
X_24923_ _24508_/CLK _15555_/X HRESETn VGND VGND VPWR VPWR _24923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24854_ _24907_/CLK _15772_/X HRESETn VGND VGND VPWR VPWR _21017_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__18299__A1_N _17731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15788__A3 _15702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_215_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ _23806_/CLK _23805_/D VGND VGND VPWR VPWR _23805_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24785_ _24886_/CLK _24785_/D HRESETn VGND VGND VPWR VPWR _24785_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_199_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _21997_/A _20318_/X VGND VGND VPWR VPWR _21997_/X sky130_fd_sc_hd__and2_4
XFILLER_214_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23180__A1 _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ HWDATA[10] VGND VGND VPWR VPWR _15965_/A sky130_fd_sc_hd__buf_2
X_23736_ _23735_/CLK _19441_/X VGND VGND VPWR VPWR _18039_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_42_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20953_/B VGND VGND VPWR VPWR _20948_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_216_0_HCLK clkbuf_7_108_0_HCLK/X VGND VGND VPWR VPWR _24540_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _16077_/A _11681_/B VGND VGND VPWR VPWR _11681_/X sky130_fd_sc_hd__or2_4
X_23667_ _25326_/CLK _23667_/D VGND VGND VPWR VPWR _13439_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15945__B1 _15581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _20870_/X _20878_/X _16689_/A _20875_/X VGND VGND VPWR VPWR _20879_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19136__B1 _19067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24748__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13388_/A _23867_/Q VGND VGND VPWR VPWR _13422_/B sky130_fd_sc_hd__or2_4
X_25406_ _24032_/CLK _12713_/X HRESETn VGND VGND VPWR VPWR _25406_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13232__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22618_ _22539_/A _22615_/X _22618_/C VGND VGND VPWR VPWR _22618_/X sky130_fd_sc_hd__and3_4
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23598_ _23575_/CLK _23598_/D VGND VGND VPWR VPWR _23598_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15960__A3 _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13351_ _13314_/X _13351_/B _13351_/C VGND VGND VPWR VPWR _13352_/C sky130_fd_sc_hd__and3_4
X_25337_ _25344_/CLK _13100_/X HRESETn VGND VGND VPWR VPWR _12321_/A sky130_fd_sc_hd__dfrtp_4
X_22549_ _16510_/A _22432_/X _22536_/X VGND VGND VPWR VPWR _22549_/X sky130_fd_sc_hd__o21a_4
XFILLER_155_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12302_ _25354_/Q VGND VGND VPWR VPWR _12302_/Y sky130_fd_sc_hd__inv_2
X_16070_ _16069_/Y _16065_/X _15976_/X _16065_/X VGND VGND VPWR VPWR _24718_/D sky130_fd_sc_hd__a2bb2o_4
X_13282_ _11951_/X _13263_/X _13281_/X _25332_/Q _13243_/X VGND VGND VPWR VPWR _13282_/X
+ sky130_fd_sc_hd__o32a_4
X_25268_ _24172_/CLK _13814_/X HRESETn VGND VGND VPWR VPWR _13556_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23079__C _22817_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24330__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15021_ _15214_/B _15025_/A _14898_/X _15020_/Y VGND VGND VPWR VPWR _15021_/X sky130_fd_sc_hd__a2bb2o_4
X_12233_ _12232_/Y _23036_/A _12232_/Y _23036_/A VGND VGND VPWR VPWR _12239_/B sky130_fd_sc_hd__a2bb2o_4
X_24219_ _23555_/CLK _24219_/D HRESETn VGND VGND VPWR VPWR _24219_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15159__A _15242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25199_ _25043_/CLK _14219_/X HRESETn VGND VGND VPWR VPWR _20664_/A sky130_fd_sc_hd__dfstp_4
XFILLER_151_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12164_ _14318_/A _12161_/Y _11793_/X _12161_/Y VGND VGND VPWR VPWR _25465_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22280__A _22130_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17374__A _17242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12095_ _12102_/A VGND VGND VPWR VPWR _12095_/X sky130_fd_sc_hd__buf_2
X_16972_ _16052_/A _24381_/Q _16052_/Y _16971_/Y VGND VGND VPWR VPWR _16972_/X sky130_fd_sc_hd__o22a_4
X_19760_ _19758_/Y _19754_/X _19759_/X _19740_/A VGND VGND VPWR VPWR _23627_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25536__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15923_ _15783_/X VGND VGND VPWR VPWR _15923_/X sky130_fd_sc_hd__buf_2
X_18711_ _18710_/X VGND VGND VPWR VPWR _18711_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19691_ _13152_/B VGND VGND VPWR VPWR _19691_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18642_ _24131_/Q VGND VGND VPWR VPWR _18643_/A sky130_fd_sc_hd__inv_2
X_15854_ _21064_/B VGND VGND VPWR VPWR _15855_/B sky130_fd_sc_hd__buf_2
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14436__B1 _14392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_26_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_53_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_14805_ _14805_/A VGND VGND VPWR VPWR _14805_/X sky130_fd_sc_hd__buf_2
X_18573_ _18567_/A _18567_/B VGND VGND VPWR VPWR _18574_/C sky130_fd_sc_hd__nand2_4
XANTENNA__21624__A _22199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15785_ _11681_/B _15918_/B VGND VGND VPWR VPWR _15811_/A sky130_fd_sc_hd__or2_4
X_12997_ _12989_/X _13005_/D _12990_/A VGND VGND VPWR VPWR _12997_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16718__A _16365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19375__B1 _19351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17524_ _11717_/A _17523_/A _11717_/Y _17523_/Y VGND VGND VPWR VPWR _17525_/D sky130_fd_sc_hd__o22a_4
XFILLER_45_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15141__A2_N _24584_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14736_ _14718_/A _14724_/Y _14735_/X _22043_/A _14718_/Y VGND VGND VPWR VPWR _14736_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21343__B _21343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11948_ _11948_/A _11948_/B VGND VGND VPWR VPWR _11948_/X sky130_fd_sc_hd__or2_4
XFILLER_189_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17455_ _17453_/X VGND VGND VPWR VPWR _17455_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14667_ _21252_/A VGND VGND VPWR VPWR _22069_/A sky130_fd_sc_hd__buf_2
XANTENNA__15936__B1 _15564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11879_ _11799_/X _11877_/X _11869_/A _11876_/Y VGND VGND VPWR VPWR _25515_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24489__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19127__B1 _19125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16406_ _16418_/A VGND VGND VPWR VPWR _16406_/X sky130_fd_sc_hd__buf_2
X_13618_ _18082_/A _13593_/A _13617_/X _13593_/Y VGND VGND VPWR VPWR _13618_/X sky130_fd_sc_hd__o22a_4
X_17386_ _23977_/Q _17385_/X VGND VGND VPWR VPWR _17386_/X sky130_fd_sc_hd__or2_4
X_14598_ _14550_/X _14597_/Y _14546_/X _14591_/X _25085_/Q VGND VGND VPWR VPWR _25085_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_158_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22277__A3 _21306_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24418__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19125_ _18985_/A VGND VGND VPWR VPWR _19125_/X sky130_fd_sc_hd__buf_2
XFILLER_201_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16337_ _16344_/A VGND VGND VPWR VPWR _16337_/X sky130_fd_sc_hd__buf_2
X_13549_ _13549_/A VGND VGND VPWR VPWR _22695_/A sky130_fd_sc_hd__inv_2
XFILLER_186_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16453__A _16453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19056_ _23871_/Q VGND VGND VPWR VPWR _19056_/Y sky130_fd_sc_hd__inv_2
X_16268_ _16268_/A _16270_/B VGND VGND VPWR VPWR _16268_/X sky130_fd_sc_hd__or2_4
XFILLER_173_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24071__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18007_ _18193_/A _18007_/B VGND VGND VPWR VPWR _18007_/X sky130_fd_sc_hd__or2_4
X_15219_ _15219_/A _15223_/B VGND VGND VPWR VPWR _15219_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__19764__A _19764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16199_ _16197_/Y _16198_/X _15567_/X _16198_/X VGND VGND VPWR VPWR _16199_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24000__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21788__A2 _21786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22190__A _22190_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19958_ _21208_/B _19953_/X _19874_/X _19946_/A VGND VGND VPWR VPWR _19958_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21518__B _21419_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_108_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_108_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16010__A1_N _16009_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22737__B2 _21317_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18909_ _18909_/A VGND VGND VPWR VPWR _18909_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19889_ _19888_/Y _19884_/X _19613_/X _19884_/X VGND VGND VPWR VPWR _19889_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21920_ _21920_/A VGND VGND VPWR VPWR _21926_/A sky130_fd_sc_hd__buf_2
XFILLER_216_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14427__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18651__A2_N _24143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21851_ _21851_/A _21847_/Y _21851_/C _21851_/D VGND VGND VPWR VPWR _21851_/X sky130_fd_sc_hd__and4_4
XFILLER_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20802_ _13106_/B _20797_/X VGND VGND VPWR VPWR _20802_/X sky130_fd_sc_hd__or2_4
X_21782_ _22228_/A _21774_/X _21781_/X VGND VGND VPWR VPWR _21782_/X sky130_fd_sc_hd__or3_4
X_24570_ _24573_/CLK _16478_/X HRESETn VGND VGND VPWR VPWR _16477_/A sky130_fd_sc_hd__dfrtp_4
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23521_ _23912_/CLK _20057_/X VGND VGND VPWR VPWR _13214_/B sky130_fd_sc_hd__dfxtp_4
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20733_ _13118_/A _13117_/X _20732_/Y VGND VGND VPWR VPWR _20733_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24841__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20664_ _20664_/A _17401_/A VGND VGND VPWR VPWR _20664_/X sky130_fd_sc_hd__or2_4
X_23452_ _23452_/CLK _23452_/D VGND VGND VPWR VPWR _13392_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22365__A _22365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24159__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_46_0_HCLK clkbuf_8_47_0_HCLK/A VGND VGND VPWR VPWR _24208_/CLK sky130_fd_sc_hd__clkbuf_1
X_22403_ _21284_/X _22399_/Y _21515_/Y _22402_/X VGND VGND VPWR VPWR _22403_/X sky130_fd_sc_hd__a2bb2o_4
X_23383_ _24413_/CLK _20413_/X VGND VGND VPWR VPWR _20412_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23229__A1_N _12264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20595_ _14083_/A _20595_/B _20595_/C VGND VGND VPWR VPWR _20595_/X sky130_fd_sc_hd__and3_4
XANTENNA__12891__A _12801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16363__A _16363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25122_ _23927_/CLK _25122_/D HRESETn VGND VGND VPWR VPWR _25122_/Q sky130_fd_sc_hd__dfrtp_4
X_22334_ _22327_/Y _22329_/Y _22330_/X _22333_/Y _21556_/Y VGND VGND VPWR VPWR _22334_/X
+ sky130_fd_sc_hd__o41a_4
X_22265_ _21954_/A _22257_/X _22264_/X VGND VGND VPWR VPWR _22265_/X sky130_fd_sc_hd__and3_4
X_25053_ _25052_/CLK _25053_/D HRESETn VGND VGND VPWR VPWR _14812_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__22425__B1 _22424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21216_ _21216_/A _21215_/X VGND VGND VPWR VPWR _21216_/X sky130_fd_sc_hd__or2_4
X_24004_ _24662_/CLK _20695_/Y HRESETn VGND VGND VPWR VPWR _13110_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22196_ _22196_/A VGND VGND VPWR VPWR _22226_/A sky130_fd_sc_hd__buf_2
XFILLER_144_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22440__A3 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21147_ _25488_/Q _12081_/A _25297_/Q _13457_/D VGND VGND VPWR VPWR _21147_/X sky130_fd_sc_hd__o22a_4
XFILLER_160_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14611__A _14610_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21078_ _21078_/A _22423_/A VGND VGND VPWR VPWR _21078_/X sky130_fd_sc_hd__or2_4
X_12920_ _12920_/A _12919_/X VGND VGND VPWR VPWR _12920_/X sky130_fd_sc_hd__or2_4
X_20029_ _20029_/A VGND VGND VPWR VPWR _21201_/B sky130_fd_sc_hd__inv_2
X_24906_ _24907_/CLK _15602_/X HRESETn VGND VGND VPWR VPWR _15600_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13227__A _13421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14418__B1 _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12851_ _12851_/A _12851_/B VGND VGND VPWR VPWR _12851_/X sky130_fd_sc_hd__or2_4
X_24837_ _24809_/CLK _24837_/D HRESETn VGND VGND VPWR VPWR _24837_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16538__A _24546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24929__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11802_/A VGND VGND VPWR VPWR _11802_/Y sky130_fd_sc_hd__inv_2
XPHY_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15553_/A VGND VGND VPWR VPWR _15570_/X sky130_fd_sc_hd__buf_2
XFILLER_199_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _25385_/Q _12780_/Y _12781_/Y _22130_/A VGND VGND VPWR VPWR _12782_/X sky130_fd_sc_hd__a2bb2o_4
X_24768_ _24765_/CLK _24768_/D HRESETn VGND VGND VPWR VPWR _24768_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21164__B1 _14179_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _25102_/Q _14499_/X _23393_/Q _14494_/X VGND VGND VPWR VPWR _14521_/X sky130_fd_sc_hd__o22a_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11766_/A VGND VGND VPWR VPWR _11733_/X sky130_fd_sc_hd__buf_2
X_23719_ _23406_/CLK _23719_/D VGND VGND VPWR VPWR _23719_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24699_ _24753_/CLK _16119_/X HRESETn VGND VGND VPWR VPWR _22870_/A sky130_fd_sc_hd__dfrtp_4
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24582__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _17237_/Y _17346_/C _17345_/A _17240_/D VGND VGND VPWR VPWR _17240_/X sky130_fd_sc_hd__or4_4
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _25125_/Q VGND VGND VPWR VPWR _14452_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _16366_/A _11664_/B VGND VGND VPWR VPWR _16077_/A sky130_fd_sc_hd__or2_4
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22275__A _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24511__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _13264_/X _19666_/A VGND VGND VPWR VPWR _13403_/X sky130_fd_sc_hd__or2_4
XFILLER_186_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17171_ _17171_/A VGND VGND VPWR VPWR _17171_/Y sky130_fd_sc_hd__inv_2
XFILLER_168_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22706__C _21864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22664__B1 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383_ _14083_/A _14370_/B VGND VGND VPWR VPWR _14383_/X sky130_fd_sc_hd__or2_4
XANTENNA__16273__A _16272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16122_ _22778_/A VGND VGND VPWR VPWR _16122_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _13334_/A _13334_/B VGND VGND VPWR VPWR _13334_/X sky130_fd_sc_hd__or2_4
XFILLER_183_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15802__A1_N _12356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15146__B2 _24600_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16053_ _16052_/Y _16050_/X _15754_/X _16050_/X VGND VGND VPWR VPWR _24724_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13265_ _13264_/X _19656_/A VGND VGND VPWR VPWR _13267_/B sky130_fd_sc_hd__or2_4
X_15004_ _25016_/Q _24454_/Q _15254_/A _15003_/Y VGND VGND VPWR VPWR _15007_/C sky130_fd_sc_hd__o22a_4
XFILLER_124_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12216_ _24765_/Q VGND VGND VPWR VPWR _12216_/Y sky130_fd_sc_hd__inv_2
X_13196_ _13289_/A VGND VGND VPWR VPWR _13252_/A sky130_fd_sc_hd__buf_2
X_19812_ _23608_/Q VGND VGND VPWR VPWR _19812_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_HCLK_A HCLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12147_ _12147_/A VGND VGND VPWR VPWR _20971_/B sky130_fd_sc_hd__buf_2
XFILLER_151_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25370__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19743_ HWDATA[6] VGND VGND VPWR VPWR _19743_/X sky130_fd_sc_hd__buf_2
X_12078_ _12078_/A VGND VGND VPWR VPWR _12078_/Y sky130_fd_sc_hd__inv_2
X_16955_ _16044_/Y _24384_/Q _16044_/Y _24384_/Q VGND VGND VPWR VPWR _16955_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15906_ _14764_/X _15904_/Y _15905_/X VGND VGND VPWR VPWR _15906_/X sky130_fd_sc_hd__o21a_4
X_16886_ _16884_/Y _16877_/X _16885_/X _14777_/X VGND VGND VPWR VPWR _16886_/X sky130_fd_sc_hd__a2bb2o_4
X_19674_ _19670_/Y _19673_/X _19652_/X _19673_/X VGND VGND VPWR VPWR _19674_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14409__B1 _14407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15837_ _15642_/X _15761_/X _15770_/X _24819_/Q _15836_/X VGND VGND VPWR VPWR _15837_/X
+ sky130_fd_sc_hd__a32o_4
X_18625_ _24133_/Q VGND VGND VPWR VPWR _18686_/A sky130_fd_sc_hd__inv_2
XANTENNA__15080__A2_N _16404_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16448__A _16721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15768_ _15745_/X _15761_/X _15643_/X _24855_/Q _15706_/X VGND VGND VPWR VPWR _24855_/D
+ sky130_fd_sc_hd__a32o_4
X_18556_ _18556_/A _18556_/B VGND VGND VPWR VPWR _18557_/C sky130_fd_sc_hd__or2_4
XFILLER_206_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14719_ _14697_/A _14664_/X _14715_/Y _13726_/A _14718_/Y VGND VGND VPWR VPWR _25069_/D
+ sky130_fd_sc_hd__a32o_4
X_17507_ _17507_/A VGND VGND VPWR VPWR _17569_/A sky130_fd_sc_hd__inv_2
X_18487_ _18497_/A _18487_/B _18487_/C VGND VGND VPWR VPWR _24189_/D sky130_fd_sc_hd__and3_4
XANTENNA__19759__A _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15699_ _15836_/B VGND VGND VPWR VPWR _15699_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17438_ _14212_/B _17438_/B VGND VGND VPWR VPWR _17438_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__14188__A2 _14185_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24252__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12199__A1 _12197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_5_0_HCLK clkbuf_8_5_0_HCLK/A VGND VGND VPWR VPWR _23406_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_165_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17369_ _24346_/Q _17369_/B VGND VGND VPWR VPWR _17370_/C sky130_fd_sc_hd__or2_4
XANTENNA__17279__A _17333_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22655__B1 _24833_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16183__A _16368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19108_ _23853_/Q VGND VGND VPWR VPWR _19108_/Y sky130_fd_sc_hd__inv_2
X_20380_ _20372_/X _20368_/X _20061_/X _23396_/Q _20370_/X VGND VGND VPWR VPWR _23396_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_118_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19039_ _23877_/Q VGND VGND VPWR VPWR _19039_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22407__B1 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16911__A _24277_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22050_ _21511_/X _23342_/B VGND VGND VPWR VPWR _22050_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22958__B2 _22846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21001_ _21000_/A _21000_/B _24336_/Q _21000_/X VGND VGND VPWR VPWR _21001_/X sky130_fd_sc_hd__o22a_4
XFILLER_99_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25040__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17742__A _24288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22952_ _22952_/A VGND VGND VPWR VPWR _22952_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20197__B2 _20180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21903_ _22225_/A _19907_/Y VGND VGND VPWR VPWR _21903_/X sky130_fd_sc_hd__or2_4
X_22883_ _22883_/A _22800_/B VGND VGND VPWR VPWR _22883_/X sky130_fd_sc_hd__or2_4
XFILLER_216_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16358__A _18951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19339__B1 _19295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24622_ _25521_/CLK _16335_/X HRESETn VGND VGND VPWR VPWR _24622_/Q sky130_fd_sc_hd__dfrtp_4
X_21834_ _13114_/A _21832_/X _15625_/A _21833_/X VGND VGND VPWR VPWR _21834_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_102_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24553_ _24555_/CLK _24553_/D HRESETn VGND VGND VPWR VPWR _16520_/A sky130_fd_sc_hd__dfrtp_4
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21765_ _21761_/X _21764_/X _14744_/X VGND VGND VPWR VPWR _21765_/X sky130_fd_sc_hd__o21a_4
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23504_ _23490_/CLK _20097_/X VGND VGND VPWR VPWR _23504_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20716_ _20716_/A VGND VGND VPWR VPWR _20716_/X sky130_fd_sc_hd__buf_2
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24484_ _24486_/CLK _16705_/X HRESETn VGND VGND VPWR VPWR _24484_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_178_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16573__B1 _16397_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21696_ _21689_/Y _21695_/Y _22041_/A VGND VGND VPWR VPWR _21697_/D sky130_fd_sc_hd__o21a_4
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21449__A1 _17880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23435_ _24317_/CLK _20282_/X VGND VGND VPWR VPWR _23435_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_137_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20647_ _20646_/X VGND VGND VPWR VPWR _23981_/D sky130_fd_sc_hd__inv_2
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20578_ _14417_/Y _20566_/X _20557_/X _20577_/X VGND VGND VPWR VPWR _20578_/X sky130_fd_sc_hd__a211o_4
X_23366_ _21013_/X VGND VGND VPWR VPWR IRQ[22] sky130_fd_sc_hd__buf_2
XANTENNA__12231__A1_N _12418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22823__A _22946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25105_ _25146_/CLK _25105_/D HRESETn VGND VGND VPWR VPWR _25105_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23975__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22317_ _22317_/A VGND VGND VPWR VPWR _22317_/Y sky130_fd_sc_hd__inv_2
X_23297_ _23297_/A _23022_/B VGND VGND VPWR VPWR _23297_/X sky130_fd_sc_hd__or2_4
XFILLER_164_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22949__B2 _22290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13050_ _13048_/A _13046_/X _13050_/C VGND VGND VPWR VPWR _13050_/X sky130_fd_sc_hd__and3_4
X_25036_ _25015_/CLK _25036_/D HRESETn VGND VGND VPWR VPWR _25036_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22248_ _21674_/X _22248_/B _22247_/X VGND VGND VPWR VPWR _22249_/C sky130_fd_sc_hd__and3_4
XFILLER_105_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14351__A2 _14340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25128__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22413__A3 _21306_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16540__B _16540_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12001_ _12001_/A _11981_/A VGND VGND VPWR VPWR _12002_/A sky130_fd_sc_hd__and2_4
X_22179_ _21569_/X _22177_/X _21575_/X _22178_/X VGND VGND VPWR VPWR _22179_/X sky130_fd_sc_hd__o22a_4
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18748__A _18658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16740_ _15037_/Y _16735_/X _16386_/X _16739_/X VGND VGND VPWR VPWR _24470_/D sky130_fd_sc_hd__a2bb2o_4
X_13952_ _14238_/A _13952_/B VGND VGND VPWR VPWR _15424_/C sky130_fd_sc_hd__or2_4
XFILLER_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18467__B _18467_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12903_ _12741_/X _12892_/B VGND VGND VPWR VPWR _12907_/A sky130_fd_sc_hd__or2_4
XFILLER_47_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16671_ _16670_/Y _16668_/X _16397_/X _16668_/X VGND VGND VPWR VPWR _24498_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13883_ _13883_/A VGND VGND VPWR VPWR _13883_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12796__A _12796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24763__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15622_ _15608_/A VGND VGND VPWR VPWR _15622_/X sky130_fd_sc_hd__buf_2
X_18410_ _24655_/Q _18409_/A _16247_/Y _18409_/Y VGND VGND VPWR VPWR _18415_/B sky130_fd_sc_hd__o22a_4
X_12834_ _12834_/A _12755_/Y _12834_/C _12833_/X VGND VGND VPWR VPWR _12834_/X sky130_fd_sc_hd__or4_4
X_19390_ _19386_/Y _19389_/X _19301_/X _19389_/X VGND VGND VPWR VPWR _19390_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18341_ _18341_/A VGND VGND VPWR VPWR _18341_/Y sky130_fd_sc_hd__inv_2
X_15553_ _15553_/A VGND VGND VPWR VPWR _15553_/X sky130_fd_sc_hd__buf_2
X_12765_ _12754_/X _12765_/B _12761_/X _12765_/D VGND VGND VPWR VPWR _12779_/C sky130_fd_sc_hd__or4_4
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14491_/X _14503_/X VGND VGND VPWR VPWR _14504_/X sky130_fd_sc_hd__or2_4
XANTENNA__22717__B _22708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19750__B1 _19702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11713_/Y _11714_/X _11715_/X _11714_/X VGND VGND VPWR VPWR _25539_/D sky130_fd_sc_hd__a2bb2o_4
X_18272_ _13768_/X VGND VGND VPWR VPWR _21281_/B sky130_fd_sc_hd__buf_2
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _24070_/D VGND VGND VPWR VPWR _15511_/A sky130_fd_sc_hd__inv_2
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A _12696_/B VGND VGND VPWR VPWR _12697_/B sky130_fd_sc_hd__or2_4
XFILLER_203_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17223_ _16281_/Y _24371_/Q _16281_/Y _24371_/Q VGND VGND VPWR VPWR _17223_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ _25133_/Q VGND VGND VPWR VPWR _14435_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13420__A _13388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11928__B2 _11897_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17154_ _17125_/A _17153_/B VGND VGND VPWR VPWR _17154_/X sky130_fd_sc_hd__or2_4
X_14366_ _14366_/A _21343_/A VGND VGND VPWR VPWR _14366_/X sky130_fd_sc_hd__or2_4
XANTENNA__16316__B1 _15953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20112__B2 _20088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_92_0_HCLK clkbuf_7_46_0_HCLK/X VGND VGND VPWR VPWR _24809_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22733__A _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22652__A3 _22138_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16105_ _16103_/Y _16099_/X _15939_/X _16104_/X VGND VGND VPWR VPWR _24705_/D sky130_fd_sc_hd__a2bb2o_4
X_13317_ _13350_/A _19791_/A VGND VGND VPWR VPWR _13318_/C sky130_fd_sc_hd__or2_4
X_17085_ _17381_/B _17085_/B _17084_/X VGND VGND VPWR VPWR _17085_/X sky130_fd_sc_hd__or3_4
X_14297_ MSO_S2 _14296_/X _25177_/Q _14291_/X VGND VGND VPWR VPWR _14297_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_170_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16036_ _16035_/Y _16033_/X _11730_/X _16033_/X VGND VGND VPWR VPWR _16036_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15756__A1_N _12524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13248_ _13285_/A _23872_/Q VGND VGND VPWR VPWR _13251_/B sky130_fd_sc_hd__or2_4
XANTENNA__21349__A _21349_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13179_ _13179_/A _13179_/B _13179_/C VGND VGND VPWR VPWR _13179_/X sky130_fd_sc_hd__and3_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17987_ _14639_/A VGND VGND VPWR VPWR _17987_/X sky130_fd_sc_hd__buf_2
XANTENNA__22168__A2 _21365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18658__A _24146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19726_ _19725_/Y _19723_/X _19702_/X _19723_/X VGND VGND VPWR VPWR _23639_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16938_ _24278_/Q VGND VGND VPWR VPWR _16938_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21084__A _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19657_ _19650_/Y VGND VGND VPWR VPWR _19657_/X sky130_fd_sc_hd__buf_2
X_16869_ _16863_/A VGND VGND VPWR VPWR _16869_/X sky130_fd_sc_hd__buf_2
XFILLER_65_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18608_ _16578_/Y _24142_/Q _16578_/Y _24142_/Q VGND VGND VPWR VPWR _18608_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19588_ _19586_/Y _19581_/X _19587_/X _19581_/X VGND VGND VPWR VPWR _23686_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22908__A _22136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24433__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18539_ _18467_/B _18538_/X VGND VGND VPWR VPWR _18540_/B sky130_fd_sc_hd__or2_4
XFILLER_240_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16906__A _16906_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15810__A _11706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21550_ _21346_/A VGND VGND VPWR VPWR _22119_/B sky130_fd_sc_hd__buf_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20501_ _20495_/X _20501_/B VGND VGND VPWR VPWR _20501_/X sky130_fd_sc_hd__or2_4
XFILLER_194_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21481_ _22262_/A VGND VGND VPWR VPWR _21677_/A sky130_fd_sc_hd__buf_2
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20432_ _14369_/B VGND VGND VPWR VPWR _20455_/C sky130_fd_sc_hd__inv_2
X_23220_ _21868_/X _23219_/X _22477_/X _24883_/Q _21871_/X VGND VGND VPWR VPWR _23221_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_165_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16307__B1 _16020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20363_ _21671_/B _20362_/X _19617_/A _20362_/X VGND VGND VPWR VPWR _20363_/X sky130_fd_sc_hd__a2bb2o_4
X_23151_ _16291_/A _22904_/X VGND VGND VPWR VPWR _23151_/X sky130_fd_sc_hd__or2_4
XFILLER_162_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25292__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16641__A _16660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_0_0_HCLK clkbuf_5_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_0_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_22102_ _20462_/A _21849_/X VGND VGND VPWR VPWR _22109_/A sky130_fd_sc_hd__nor2_4
X_23082_ _12759_/Y _21879_/X _16906_/Y _22826_/X VGND VGND VPWR VPWR _23082_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21259__A _22056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20294_ _22034_/B _20288_/X _19970_/X _20293_/X VGND VGND VPWR VPWR _23431_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22033_ _22014_/A _22033_/B VGND VGND VPWR VPWR _22033_/X sky130_fd_sc_hd__or2_4
XANTENNA__11785__A _11785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17807__B1 _16940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18568__A _18400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23984_ _25050_/CLK _20659_/Y HRESETn VGND VGND VPWR VPWR _17393_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22935_ _14922_/A _22807_/X _21737_/X _22934_/X VGND VGND VPWR VPWR _22936_/C sky130_fd_sc_hd__a211o_4
XFILLER_228_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_7_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22866_ _22486_/X _22864_/X _22489_/X _24734_/Q _22865_/X VGND VGND VPWR VPWR _22866_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24174__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24605_ _24551_/CLK _24605_/D HRESETn VGND VGND VPWR VPWR _24605_/Q sky130_fd_sc_hd__dfrtp_4
X_21817_ _21817_/A _21817_/B VGND VGND VPWR VPWR _21818_/C sky130_fd_sc_hd__or2_4
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22797_ _21283_/A _21955_/A _22619_/B _22520_/A VGND VGND VPWR VPWR _22798_/A sky130_fd_sc_hd__a211o_4
XFILLER_197_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24103__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19732__B1 _19708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12550_ _12550_/A VGND VGND VPWR VPWR _12550_/Y sky130_fd_sc_hd__inv_2
X_24536_ _24573_/CLK _16568_/X HRESETn VGND VGND VPWR VPWR _16566_/A sky130_fd_sc_hd__dfrtp_4
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21748_ _21748_/A _21747_/X VGND VGND VPWR VPWR _21748_/Y sky130_fd_sc_hd__nor2_4
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _12475_/B VGND VGND VPWR VPWR _12482_/B sky130_fd_sc_hd__inv_2
X_24467_ _24443_/CLK _24467_/D HRESETn VGND VGND VPWR VPWR _15020_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21679_ _21673_/X _21678_/X _21489_/X VGND VGND VPWR VPWR _21679_/X sky130_fd_sc_hd__o21a_4
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ _25198_/Q VGND VGND VPWR VPWR _14220_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_16_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_16_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23418_ _23425_/CLK _20325_/X VGND VGND VPWR VPWR _21214_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_138_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18299__B1 _17731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24398_ _24377_/CLK _17078_/X HRESETn VGND VGND VPWR VPWR _24398_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_79_0_HCLK clkbuf_7_79_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_79_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14151_ _14102_/C _14087_/X _14102_/C _14087_/X VGND VGND VPWR VPWR _14151_/X sky130_fd_sc_hd__a2bb2o_4
X_23349_ _25325_/Q _25297_/Q VGND VGND VPWR VPWR _23349_/X sky130_fd_sc_hd__and2_4
XFILLER_180_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13102_ _12982_/A _13101_/Y VGND VGND VPWR VPWR _13102_/X sky130_fd_sc_hd__or2_4
XFILLER_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14082_ _24002_/Q _14067_/A _14062_/X _14012_/A _14049_/B VGND VGND VPWR VPWR _25226_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_180_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19799__B1 _19711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13033_ _12357_/Y _13032_/X VGND VGND VPWR VPWR _13033_/X sky130_fd_sc_hd__or2_4
X_17910_ _21993_/A _17910_/B VGND VGND VPWR VPWR _17910_/X sky130_fd_sc_hd__or2_4
X_25019_ _24967_/CLK _15250_/X HRESETn VGND VGND VPWR VPWR _25019_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11695__A HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18890_ _18871_/X _18885_/X _20984_/B _24123_/Q _18888_/X VGND VGND VPWR VPWR _18890_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_121_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17841_ _17756_/Y _17841_/B VGND VGND VPWR VPWR _17842_/A sky130_fd_sc_hd__or2_4
XFILLER_239_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24944__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14984_ _15229_/A _24461_/Q _15229_/A _24461_/Q VGND VGND VPWR VPWR _14984_/X sky130_fd_sc_hd__a2bb2o_4
X_17772_ _17790_/A _17772_/B _17772_/C VGND VGND VPWR VPWR _17772_/X sky130_fd_sc_hd__and3_4
X_19511_ _21948_/B _19508_/X _11915_/X _19508_/X VGND VGND VPWR VPWR _19511_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13935_ _13935_/A _13935_/B _13934_/X _13942_/C VGND VGND VPWR VPWR _13935_/X sky130_fd_sc_hd__or4_4
X_16723_ _24477_/Q VGND VGND VPWR VPWR _16723_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16654_ _24504_/Q VGND VGND VPWR VPWR _16654_/Y sky130_fd_sc_hd__inv_2
X_19442_ _19442_/A VGND VGND VPWR VPWR _19442_/Y sky130_fd_sc_hd__inv_2
X_13866_ _13860_/X _13865_/X _14256_/A _13856_/X VGND VGND VPWR VPWR _13866_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16785__B1 _16435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15605_ _24904_/Q VGND VGND VPWR VPWR _15605_/Y sky130_fd_sc_hd__inv_2
X_12817_ _12816_/Y _24788_/Q _25369_/Q _12783_/Y VGND VGND VPWR VPWR _12823_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16585_ _16598_/A VGND VGND VPWR VPWR _16585_/X sky130_fd_sc_hd__buf_2
X_19373_ _19371_/Y _19367_/X _19282_/X _19372_/X VGND VGND VPWR VPWR _23760_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_222_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13797_ _13797_/A VGND VGND VPWR VPWR _16361_/A sky130_fd_sc_hd__buf_2
XFILLER_90_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15536_ _15535_/Y _15533_/X HADDR[1] _15533_/X VGND VGND VPWR VPWR _15536_/X sky130_fd_sc_hd__a2bb2o_4
X_18324_ _20387_/A VGND VGND VPWR VPWR _19209_/A sky130_fd_sc_hd__buf_2
X_12748_ _12895_/A _12746_/Y _12735_/A _12747_/Y VGND VGND VPWR VPWR _12751_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16537__B1 _16361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20248__A _20243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18255_ _18238_/X _18240_/X _15830_/X _24230_/Q _18241_/X VGND VGND VPWR VPWR _18255_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14891__D _14891_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15467_ _15465_/Y _15463_/X _15466_/X _15463_/X VGND VGND VPWR VPWR _15467_/X sky130_fd_sc_hd__a2bb2o_4
X_12679_ _12678_/X VGND VGND VPWR VPWR _12679_/Y sky130_fd_sc_hd__inv_2
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17206_ _16329_/Y _24353_/Q _16329_/Y _24353_/Q VGND VGND VPWR VPWR _17208_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13150__A _13433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14418_ _14417_/Y _14415_/X _14262_/X _14415_/X VGND VGND VPWR VPWR _25139_/D sky130_fd_sc_hd__a2bb2o_4
X_18186_ _18014_/A _23892_/Q VGND VGND VPWR VPWR _18186_/X sky130_fd_sc_hd__or2_4
X_15398_ _15379_/A _15395_/B _15398_/C VGND VGND VPWR VPWR _15398_/X sky130_fd_sc_hd__and3_4
XFILLER_116_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17137_ _17035_/A _17140_/B VGND VGND VPWR VPWR _17138_/C sky130_fd_sc_hd__nand2_4
XFILLER_162_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14349_ _14349_/A VGND VGND VPWR VPWR _14349_/X sky130_fd_sc_hd__buf_2
XFILLER_143_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17557__A _17602_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17068_ _16965_/A _17072_/B VGND VGND VPWR VPWR _17070_/B sky130_fd_sc_hd__or2_4
XANTENNA__21079__A _11701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16019_ _15998_/A VGND VGND VPWR VPWR _16019_/X sky130_fd_sc_hd__buf_2
XFILLER_143_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24685__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24614__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19709_ _19706_/Y _19707_/X _19708_/X _19707_/X VGND VGND VPWR VPWR _19709_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20981_ _14111_/X _20980_/X _14084_/Y VGND VGND VPWR VPWR _23956_/D sky130_fd_sc_hd__o21a_4
XFILLER_65_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_0_0_HCLK_A clkbuf_3_0_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18765__A1 _18692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22720_ _16128_/Y _22718_/X _22719_/X _11732_/Y _22279_/X VGND VGND VPWR VPWR _22720_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_213_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16776__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21542__A _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22651_ _24625_/Q _22654_/B VGND VGND VPWR VPWR _22651_/X sky130_fd_sc_hd__or2_4
XANTENNA__24121__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19714__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21602_ _22219_/A VGND VGND VPWR VPWR _21769_/A sky130_fd_sc_hd__buf_2
XANTENNA__15540__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25370_ _25375_/CLK _25370_/D HRESETn VGND VGND VPWR VPWR _25370_/Q sky130_fd_sc_hd__dfrtp_4
X_22582_ _22582_/A VGND VGND VPWR VPWR _22619_/B sky130_fd_sc_hd__buf_2
XFILLER_178_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24321_ _24317_/CLK _17595_/Y HRESETn VGND VGND VPWR VPWR _17549_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21533_ _21533_/A VGND VGND VPWR VPWR _23172_/A sky130_fd_sc_hd__buf_2
XFILLER_178_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24252_ _24252_/CLK _24252_/D HRESETn VGND VGND VPWR VPWR _13528_/C sky130_fd_sc_hd__dfrtp_4
X_21464_ _21661_/A _19871_/Y VGND VGND VPWR VPWR _21468_/B sky130_fd_sc_hd__or2_4
XANTENNA__25402__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23203_ _23235_/A _23203_/B VGND VGND VPWR VPWR _23203_/Y sky130_fd_sc_hd__nor2_4
XFILLER_147_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12565__B2 _24870_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20415_ _20409_/Y VGND VGND VPWR VPWR _20415_/X sky130_fd_sc_hd__buf_2
XFILLER_134_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21395_ _14688_/A _21393_/X _21395_/C VGND VGND VPWR VPWR _21395_/X sky130_fd_sc_hd__and3_4
X_24183_ _24188_/CLK _18514_/X HRESETn VGND VGND VPWR VPWR _18461_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_162_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23134_ _16472_/A _22885_/X _23133_/X VGND VGND VPWR VPWR _23134_/X sky130_fd_sc_hd__o21a_4
XFILLER_134_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20346_ _20345_/Y _20341_/X _20008_/X _20328_/Y VGND VGND VPWR VPWR _20346_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16700__B1 _16518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12317__B2 _12316_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20277_ _21792_/B _20272_/X _19977_/X _20272_/X VGND VGND VPWR VPWR _23437_/D sky130_fd_sc_hd__a2bb2o_4
X_23065_ _16477_/A _22885_/X _22802_/X VGND VGND VPWR VPWR _23065_/X sky130_fd_sc_hd__o21a_4
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12404__A _12194_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22016_ _22016_/A _22016_/B VGND VGND VPWR VPWR _22017_/C sky130_fd_sc_hd__or2_4
XANTENNA__21052__A2 _21031_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24355__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11981_ _11981_/A VGND VGND VPWR VPWR _11981_/Y sky130_fd_sc_hd__inv_2
X_23967_ _24973_/CLK _21011_/X HRESETn VGND VGND VPWR VPWR _23967_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15019__B1 _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18756__A1 _18693_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13720_ _11836_/A _13708_/X _13690_/X _13668_/B VGND VGND VPWR VPWR _25281_/D sky130_fd_sc_hd__o22a_4
X_22918_ _17251_/C _22916_/X _12766_/A _22917_/X VGND VGND VPWR VPWR _22918_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16767__B1 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23898_ _23827_/CLK _23898_/D VGND VGND VPWR VPWR _17937_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13651_ _13651_/A _13637_/X _13650_/X VGND VGND VPWR VPWR _13651_/X sky130_fd_sc_hd__or3_4
X_22849_ _22130_/B VGND VGND VPWR VPWR _22849_/X sky130_fd_sc_hd__buf_2
XFILLER_140_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16546__A _24544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19705__B1 _19587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12602_ _12584_/X _12717_/A _12498_/Y _12697_/A VGND VGND VPWR VPWR _12605_/B sky130_fd_sc_hd__or4_4
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16370_ _16370_/A VGND VGND VPWR VPWR _16370_/X sky130_fd_sc_hd__buf_2
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21171__B _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13582_ _19522_/A VGND VGND VPWR VPWR _19570_/A sky130_fd_sc_hd__buf_2
XFILLER_169_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16519__B1 _16518_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ _15315_/A _15320_/X _15313_/A _15316_/Y VGND VGND VPWR VPWR _15322_/A sky130_fd_sc_hd__a211o_4
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23990__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12533_ _12623_/A VGND VGND VPWR VPWR _12624_/A sky130_fd_sc_hd__inv_2
X_24519_ _24520_/CLK _24519_/D HRESETn VGND VGND VPWR VPWR _16610_/A sky130_fd_sc_hd__dfrtp_4
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25499_ _25499_/CLK _25499_/D HRESETn VGND VGND VPWR VPWR _11931_/A sky130_fd_sc_hd__dfrtp_4
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18040_ _18151_/A _18040_/B VGND VGND VPWR VPWR _18041_/C sky130_fd_sc_hd__or2_4
X_15252_ _15246_/C _15251_/X _15185_/A _15248_/B VGND VGND VPWR VPWR _15253_/A sky130_fd_sc_hd__a211o_4
XFILLER_8_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12464_ _12480_/A _12464_/B _12463_/X VGND VGND VPWR VPWR _25444_/D sky130_fd_sc_hd__and3_4
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ _14203_/A VGND VGND VPWR VPWR _14203_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22714__C _21864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17377__A _17242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12556__B2 _24869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15183_ _15165_/A _15181_/X _15183_/C VGND VGND VPWR VPWR _15183_/X sky130_fd_sc_hd__and3_4
XFILLER_126_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12395_ _12170_/A _12400_/B VGND VGND VPWR VPWR _12395_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_4_11_0_HCLK_A clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14134_ _14114_/X _14132_/Y _14091_/A _14133_/X VGND VGND VPWR VPWR _25220_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19991_ _19990_/Y VGND VGND VPWR VPWR _19991_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_103_0_HCLK clkbuf_7_51_0_HCLK/X VGND VGND VPWR VPWR _24763_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_152_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14065_ _14049_/B VGND VGND VPWR VPWR _14065_/X sky130_fd_sc_hd__buf_2
X_18942_ _18942_/A VGND VGND VPWR VPWR _18942_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_166_0_HCLK clkbuf_7_83_0_HCLK/X VGND VGND VPWR VPWR _23889_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_9_0_HCLK clkbuf_7_9_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_13016_ _12971_/Y _12985_/X _12349_/Y _12978_/X VGND VGND VPWR VPWR _13016_/X sky130_fd_sc_hd__or4_4
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21627__A _21627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18873_ _23939_/Q _18872_/X VGND VGND VPWR VPWR _20553_/A sky130_fd_sc_hd__or2_4
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17824_ _17760_/Y _17813_/B VGND VGND VPWR VPWR _17828_/A sky130_fd_sc_hd__or2_4
XFILLER_227_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18001__A _18054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24096__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14967_ _25028_/Q VGND VGND VPWR VPWR _15207_/A sky130_fd_sc_hd__inv_2
X_17755_ _17755_/A VGND VGND VPWR VPWR _17755_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24025__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13145__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16706_ _16706_/A VGND VGND VPWR VPWR _16706_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17840__A _17602_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13918_ _13947_/C VGND VGND VPWR VPWR _13923_/D sky130_fd_sc_hd__buf_2
XFILLER_223_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14898_ _14898_/A VGND VGND VPWR VPWR _14898_/X sky130_fd_sc_hd__buf_2
X_17686_ _17686_/A VGND VGND VPWR VPWR _17687_/B sky130_fd_sc_hd__inv_2
XFILLER_223_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16758__B1 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16993__A1_N _16042_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19425_ _18143_/B VGND VGND VPWR VPWR _19425_/Y sky130_fd_sc_hd__inv_2
X_13849_ _13839_/A VGND VGND VPWR VPWR _13849_/X sky130_fd_sc_hd__buf_2
X_16637_ _16637_/A _15671_/A VGND VGND VPWR VPWR _16640_/A sky130_fd_sc_hd__or2_4
XFILLER_222_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19356_ _19343_/A VGND VGND VPWR VPWR _19356_/X sky130_fd_sc_hd__buf_2
X_16568_ _16566_/Y _16567_/X _16483_/X _16567_/X VGND VGND VPWR VPWR _16568_/X sky130_fd_sc_hd__a2bb2o_4
X_18307_ _21475_/A _18305_/X _18306_/Y VGND VGND VPWR VPWR _24213_/D sky130_fd_sc_hd__o21a_4
X_15519_ _15530_/A VGND VGND VPWR VPWR _15519_/X sky130_fd_sc_hd__buf_2
XFILLER_149_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16499_ _16498_/Y _16496_/X _16226_/X _16496_/X VGND VGND VPWR VPWR _16499_/X sky130_fd_sc_hd__a2bb2o_4
X_19287_ _23790_/Q VGND VGND VPWR VPWR _19287_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18238_ _13807_/D VGND VGND VPWR VPWR _18238_/X sky130_fd_sc_hd__buf_2
XFILLER_176_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23256__B1 _16913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16930__B1 _16131_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18169_ _18030_/A _18169_/B _18168_/X VGND VGND VPWR VPWR _18173_/B sky130_fd_sc_hd__and3_4
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_62_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20200_ _20200_/A VGND VGND VPWR VPWR _20200_/Y sky130_fd_sc_hd__inv_2
X_21180_ _21189_/A _21180_/B VGND VGND VPWR VPWR _21181_/C sky130_fd_sc_hd__or2_4
XFILLER_116_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22921__A _16670_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24866__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15497__B1 HADDR[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20131_ _21411_/B _20128_/X _20109_/X _20128_/X VGND VGND VPWR VPWR _23492_/D sky130_fd_sc_hd__a2bb2o_4
X_20062_ _20054_/A _18328_/A _20061_/X _13367_/B _20055_/A VGND VGND VPWR VPWR _20062_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21537__A _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24870_ _24866_/CLK _24870_/D HRESETn VGND VGND VPWR VPWR _24870_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23821_ _23831_/CLK _19201_/X VGND VGND VPWR VPWR _18161_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_241_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19935__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23752_ _23785_/CLK _19397_/X VGND VGND VPWR VPWR _18036_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20964_ _11985_/X _20964_/B VGND VGND VPWR VPWR _20964_/X sky130_fd_sc_hd__and2_4
XANTENNA__20545__A1 _14158_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21742__B1 _21582_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22703_ _24428_/Q _21336_/X _15663_/A _22702_/X VGND VGND VPWR VPWR _22704_/C sky130_fd_sc_hd__a211o_4
XPHY_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23683_ _23706_/CLK _19595_/X VGND VGND VPWR VPWR _19594_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ _13650_/C _20889_/X _20894_/Y VGND VGND VPWR VPWR _20895_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__16366__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25422_ _24872_/CLK _25422_/D HRESETn VGND VGND VPWR VPWR _12657_/A sky130_fd_sc_hd__dfrtp_4
X_22634_ _21294_/X _22633_/X _21300_/A _24832_/Q _22490_/X VGND VGND VPWR VPWR _22634_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_241_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25353_ _25344_/CLK _13048_/X HRESETn VGND VGND VPWR VPWR _12324_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22565_ _22149_/X _22564_/X _22134_/A _25530_/Q _22554_/X VGND VGND VPWR VPWR _22565_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_166_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24304_ _23411_/CLK _24304_/D HRESETn VGND VGND VPWR VPWR _17659_/A sky130_fd_sc_hd__dfrtp_4
X_21516_ _21515_/Y VGND VGND VPWR VPWR _22041_/A sky130_fd_sc_hd__buf_2
X_25284_ _25285_/CLK _25284_/D HRESETn VGND VGND VPWR VPWR _11816_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23247__B1 _23235_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22496_ _11681_/B _22494_/X _22495_/X _25529_/Q _15983_/X VGND VGND VPWR VPWR _22496_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_154_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24235_ _25091_/CLK _18248_/X HRESETn VGND VGND VPWR VPWR _22517_/A sky130_fd_sc_hd__dfrtp_4
X_21447_ _11664_/B VGND VGND VPWR VPWR _21447_/X sky130_fd_sc_hd__buf_2
XANTENNA__17477__A1 _18900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12180_ _25443_/Q _12178_/Y _12278_/A _23144_/A VGND VGND VPWR VPWR _12180_/X sky130_fd_sc_hd__a2bb2o_4
X_24166_ _24650_/CLK _24166_/D HRESETn VGND VGND VPWR VPWR _18409_/A sky130_fd_sc_hd__dfrtp_4
X_21378_ _21377_/X VGND VGND VPWR VPWR _21378_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22470__B2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22831__A _23075_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15488__B1 HADDR[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23117_ _17236_/A _22916_/X _12878_/A _22917_/X VGND VGND VPWR VPWR _23117_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20329_ _20328_/Y VGND VGND VPWR VPWR _20329_/X sky130_fd_sc_hd__buf_2
X_24097_ _23388_/CLK _24097_/D HRESETn VGND VGND VPWR VPWR _24097_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24536__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_239_0_HCLK clkbuf_8_239_0_HCLK/A VGND VGND VPWR VPWR _25052_/CLK sky130_fd_sc_hd__clkbuf_1
X_23048_ _23047_/X VGND VGND VPWR VPWR _23048_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21447__A _11664_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15870_ _15843_/X _15850_/X _15725_/X _24808_/Q _15857_/X VGND VGND VPWR VPWR _24808_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_76_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21166__B _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14821_ _14830_/A VGND VGND VPWR VPWR _14826_/A sky130_fd_sc_hd__buf_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24999_ _24953_/CLK _15341_/X HRESETn VGND VGND VPWR VPWR _24999_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_236_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23183__C1 _23182_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14752_ _22202_/A VGND VGND VPWR VPWR _22225_/A sky130_fd_sc_hd__buf_2
X_17540_ _11694_/Y _24313_/Q _25530_/Q _17499_/Y VGND VGND VPWR VPWR _17540_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ _11962_/X VGND VGND VPWR VPWR _11964_/Y sky130_fd_sc_hd__inv_2
X_13703_ _11832_/Y _13675_/B VGND VGND VPWR VPWR _13703_/Y sky130_fd_sc_hd__nand2_4
X_17471_ _18911_/B _17462_/X _17469_/Y _17470_/Y VGND VGND VPWR VPWR _17472_/D sky130_fd_sc_hd__a211o_4
XFILLER_72_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14683_ _14683_/A _13736_/A VGND VGND VPWR VPWR _14683_/X sky130_fd_sc_hd__or2_4
XFILLER_205_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11895_ _19600_/A VGND VGND VPWR VPWR _11895_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16276__A _22505_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25395__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19210_ _19209_/X VGND VGND VPWR VPWR _19224_/A sky130_fd_sc_hd__inv_2
XFILLER_232_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13634_ _25300_/Q _13627_/X _13633_/Y VGND VGND VPWR VPWR _25300_/D sky130_fd_sc_hd__o21a_4
X_16422_ _16418_/A VGND VGND VPWR VPWR _16422_/X sky130_fd_sc_hd__buf_2
XANTENNA__15963__A1 _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25324__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15963__B2 _15925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16353_ _14392_/A VGND VGND VPWR VPWR _16353_/X sky130_fd_sc_hd__buf_2
X_19141_ _19411_/A _19141_/B _13615_/A _13613_/A VGND VGND VPWR VPWR _19141_/X sky130_fd_sc_hd__or4_4
X_13565_ _13565_/A _13565_/B _13561_/X _13564_/X VGND VGND VPWR VPWR _13575_/C sky130_fd_sc_hd__or4_4
XANTENNA__19587__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15304_ _15315_/A _15326_/A _15304_/C _15303_/X VGND VGND VPWR VPWR _15304_/X sky130_fd_sc_hd__or4_4
X_12516_ _12657_/A _12514_/Y _12503_/A _12515_/Y VGND VGND VPWR VPWR _12516_/X sky130_fd_sc_hd__a2bb2o_4
X_19072_ _13753_/X _13754_/X _19072_/C _13741_/D VGND VGND VPWR VPWR _19073_/A sky130_fd_sc_hd__or4_4
X_16284_ _16318_/A VGND VGND VPWR VPWR _16284_/X sky130_fd_sc_hd__buf_2
XFILLER_157_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13496_ _25310_/Q VGND VGND VPWR VPWR _13496_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15235_ _15234_/X VGND VGND VPWR VPWR _15236_/B sky130_fd_sc_hd__inv_2
X_18023_ _15691_/X _17997_/X _18021_/X _24249_/Q _18022_/X VGND VGND VPWR VPWR _18023_/X
+ sky130_fd_sc_hd__o32a_4
X_12447_ _12271_/X _12494_/A VGND VGND VPWR VPWR _12447_/X sky130_fd_sc_hd__or2_4
XFILLER_173_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_49_0_HCLK clkbuf_5_24_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_99_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15166_ _14981_/A _15242_/B VGND VGND VPWR VPWR _15167_/B sky130_fd_sc_hd__and2_4
XFILLER_5_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12378_ _12370_/X _12261_/X VGND VGND VPWR VPWR _12378_/X sky130_fd_sc_hd__and2_4
X_14117_ _14117_/A VGND VGND VPWR VPWR _14117_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15097_ _24604_/Q VGND VGND VPWR VPWR _15097_/Y sky130_fd_sc_hd__inv_2
X_19974_ _19974_/A VGND VGND VPWR VPWR _19974_/X sky130_fd_sc_hd__buf_2
XFILLER_153_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15058__C _15246_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24277__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14048_ _14073_/A VGND VGND VPWR VPWR _14049_/B sky130_fd_sc_hd__buf_2
X_18925_ _18925_/A VGND VGND VPWR VPWR _18925_/X sky130_fd_sc_hd__buf_2
XANTENNA__24206__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18856_ _18852_/X _18853_/X _18854_/X _18855_/X VGND VGND VPWR VPWR _18856_/X sky130_fd_sc_hd__or4_4
XANTENNA__16979__B1 _15995_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17807_ _17763_/X _17773_/X _16940_/Y VGND VGND VPWR VPWR _17807_/X sky130_fd_sc_hd__o21a_4
XFILLER_82_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_HCLK clkbuf_3_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_9_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_18787_ _18787_/A _18786_/X VGND VGND VPWR VPWR _18810_/A sky130_fd_sc_hd__or2_4
X_15999_ _15995_/Y _15990_/X _15996_/X _15998_/X VGND VGND VPWR VPWR _24745_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17738_ _17703_/X _17706_/A _21822_/A VGND VGND VPWR VPWR _17738_/X sky130_fd_sc_hd__or3_4
XFILLER_224_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21724__B1 _15468_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17669_ _17513_/Y _17669_/B VGND VGND VPWR VPWR _17670_/B sky130_fd_sc_hd__or2_4
XFILLER_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19408_ _17440_/A VGND VGND VPWR VPWR _19408_/X sky130_fd_sc_hd__buf_2
XANTENNA__13603__A _18095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20680_ _20675_/X _20679_/X _20613_/B VGND VGND VPWR VPWR _20680_/X sky130_fd_sc_hd__o21a_4
XFILLER_195_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25065__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22916__A _22429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12768__A1 _12766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21820__A _21954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19339_ _19338_/Y _19334_/X _19295_/X _19327_/A VGND VGND VPWR VPWR _23771_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22635__B _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22350_ _21935_/A _22350_/B VGND VGND VPWR VPWR _22350_/X sky130_fd_sc_hd__or2_4
XFILLER_137_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21301_ _21292_/X _21295_/X _21306_/C VGND VGND VPWR VPWR _21301_/X sky130_fd_sc_hd__and3_4
XFILLER_136_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22281_ _24618_/Q _22280_/X VGND VGND VPWR VPWR _22281_/X sky130_fd_sc_hd__or2_4
X_24020_ _24051_/CLK _20766_/X HRESETn VGND VGND VPWR VPWR _13107_/A sky130_fd_sc_hd__dfrtp_4
X_21232_ _15981_/A VGND VGND VPWR VPWR _21232_/X sky130_fd_sc_hd__buf_2
XFILLER_191_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14390__B1 _14389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20058__A3 _13829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17745__A _24283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21163_ _21343_/B _21162_/X _17438_/B VGND VGND VPWR VPWR _21163_/X sky130_fd_sc_hd__o21a_4
X_20114_ _20136_/A _13741_/D _19803_/X VGND VGND VPWR VPWR _20115_/A sky130_fd_sc_hd__or3_4
X_21094_ _21015_/A _21048_/Y VGND VGND VPWR VPWR _21094_/X sky130_fd_sc_hd__and2_4
XFILLER_131_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20171__A _20158_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12889__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15890__B1 _13818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11793__A _13459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20045_ _23525_/Q VGND VGND VPWR VPWR _21634_/B sky130_fd_sc_hd__inv_2
X_24922_ _24032_/CLK _15558_/X HRESETn VGND VGND VPWR VPWR _15556_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_69_0_HCLK clkbuf_7_34_0_HCLK/X VGND VGND VPWR VPWR _25444_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24853_ _24910_/CLK _15774_/X HRESETn VGND VGND VPWR VPWR _20684_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_46_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23804_ _23859_/CLK _23804_/D VGND VGND VPWR VPWR _19247_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__23929__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24784_ _24889_/CLK _24784_/D HRESETn VGND VGND VPWR VPWR _24784_/Q sky130_fd_sc_hd__dfrtp_4
X_21996_ _17893_/Y _23420_/Q _21997_/A _20318_/X VGND VGND VPWR VPWR _21996_/X sky130_fd_sc_hd__o22a_4
XPHY_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _23735_/CLK _23735_/D VGND VGND VPWR VPWR _19442_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _20947_/A VGND VGND VPWR VPWR _20947_/Y sky130_fd_sc_hd__inv_2
XFILLER_214_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14609__A _14608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _22136_/B VGND VGND VPWR VPWR _11681_/B sky130_fd_sc_hd__buf_2
X_23666_ _25326_/CLK _19653_/X VGND VGND VPWR VPWR _23666_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _20877_/Y _20871_/Y _13648_/X VGND VGND VPWR VPWR _20878_/X sky130_fd_sc_hd__o21a_4
XFILLER_198_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25405_ _24032_/CLK _12715_/Y HRESETn VGND VGND VPWR VPWR _12569_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22617_ _16831_/A _21031_/X _22533_/X _22616_/X VGND VGND VPWR VPWR _22618_/C sky130_fd_sc_hd__a211o_4
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21730__A _21730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23597_ _23526_/CLK _19848_/X VGND VGND VPWR VPWR _23597_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_197_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13350_ _13350_/A _13350_/B VGND VGND VPWR VPWR _13351_/C sky130_fd_sc_hd__or2_4
X_25336_ _25341_/CLK _25336_/D HRESETn VGND VGND VPWR VPWR _12982_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19200__A _19063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22548_ _22548_/A _16368_/A VGND VGND VPWR VPWR _22548_/X sky130_fd_sc_hd__or2_4
XFILLER_6_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12301_ _12301_/A _12295_/X _12298_/X _12301_/D VGND VGND VPWR VPWR _12328_/B sky130_fd_sc_hd__or4_4
XFILLER_127_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24788__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13281_ _13353_/A _13272_/X _13280_/X VGND VGND VPWR VPWR _13281_/X sky130_fd_sc_hd__and3_4
X_25267_ _24172_/CLK _13815_/X HRESETn VGND VGND VPWR VPWR _25267_/Q sky130_fd_sc_hd__dfrtp_4
X_22479_ _22474_/X _22476_/X _22477_/X _24829_/Q _22478_/X VGND VGND VPWR VPWR _22479_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_155_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15020_ _15020_/A VGND VGND VPWR VPWR _15020_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24717__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12232_ _25456_/Q VGND VGND VPWR VPWR _12232_/Y sky130_fd_sc_hd__inv_2
X_24218_ _25285_/CLK _24218_/D HRESETn VGND VGND VPWR VPWR _18279_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__14381__B1 _14380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25198_ _25043_/CLK _14221_/X HRESETn VGND VGND VPWR VPWR _25198_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA_clkbuf_5_3_0_HCLK_A clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12163_ _12163_/A VGND VGND VPWR VPWR _14318_/A sky130_fd_sc_hd__inv_2
X_24149_ _24146_/CLK _24149_/D HRESETn VGND VGND VPWR VPWR _24149_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24370__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21177__A _21177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12094_ _12094_/A VGND VGND VPWR VPWR _12119_/A sky130_fd_sc_hd__inv_2
X_16971_ _24381_/Q VGND VGND VPWR VPWR _16971_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18710_ _18700_/C _18707_/X _18703_/B _18709_/X VGND VGND VPWR VPWR _18710_/X sky130_fd_sc_hd__a211o_4
X_15922_ _15665_/X _15783_/X _15920_/X _12728_/A _15921_/X VGND VGND VPWR VPWR _24780_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_39_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19690_ _19689_/Y _19685_/X _19646_/X _19672_/Y VGND VGND VPWR VPWR _23651_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18641_ _18641_/A VGND VGND VPWR VPWR _18815_/A sky130_fd_sc_hd__inv_2
X_15853_ _22638_/B VGND VGND VPWR VPWR _21064_/B sky130_fd_sc_hd__buf_2
XFILLER_49_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15633__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14804_ _14830_/A VGND VGND VPWR VPWR _14805_/A sky130_fd_sc_hd__inv_2
X_18572_ _18572_/A _18568_/X _18571_/Y VGND VGND VPWR VPWR _18572_/X sky130_fd_sc_hd__and3_4
X_12996_ _13059_/A _12494_/A VGND VGND VPWR VPWR _13005_/D sky130_fd_sc_hd__and2_4
X_15784_ _15783_/X VGND VGND VPWR VPWR _15784_/X sky130_fd_sc_hd__buf_2
XFILLER_80_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25505__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17523_ _17523_/A VGND VGND VPWR VPWR _17523_/Y sky130_fd_sc_hd__inv_2
X_11947_ _11947_/A VGND VGND VPWR VPWR _11948_/A sky130_fd_sc_hd__buf_2
X_14735_ _22044_/A _14735_/B VGND VGND VPWR VPWR _14735_/X sky130_fd_sc_hd__or2_4
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14666_ _14672_/A VGND VGND VPWR VPWR _14666_/X sky130_fd_sc_hd__buf_2
X_17454_ _17451_/X VGND VGND VPWR VPWR _18342_/A sky130_fd_sc_hd__inv_2
XFILLER_220_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11878_ _11799_/X _11877_/X _11869_/A _11875_/X VGND VGND VPWR VPWR _25516_/D sky130_fd_sc_hd__a22oi_4
XFILLER_177_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13617_ _25078_/Q VGND VGND VPWR VPWR _13617_/X sky130_fd_sc_hd__buf_2
X_16405_ _16375_/A VGND VGND VPWR VPWR _16418_/A sky130_fd_sc_hd__buf_2
XFILLER_177_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_25_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_14597_ _14550_/A _14550_/B VGND VGND VPWR VPWR _14597_/Y sky130_fd_sc_hd__nand2_4
X_17385_ _17385_/A _17385_/B VGND VGND VPWR VPWR _17385_/X sky130_fd_sc_hd__or2_4
XFILLER_220_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22131__B1 _12551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19124_ _18053_/B VGND VGND VPWR VPWR _19124_/Y sky130_fd_sc_hd__inv_2
X_13548_ _25260_/Q _14553_/A _25266_/Q _14561_/A VGND VGND VPWR VPWR _13548_/X sky130_fd_sc_hd__a2bb2o_4
X_16336_ _24621_/Q VGND VGND VPWR VPWR _16336_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16267_ _13797_/A VGND VGND VPWR VPWR _16267_/X sky130_fd_sc_hd__buf_2
X_19055_ _19053_/Y _19049_/X _18985_/X _19054_/X VGND VGND VPWR VPWR _23872_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_185_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13479_ _13478_/Y _13476_/X _12076_/X _13476_/X VGND VGND VPWR VPWR _13479_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24458__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15218_ _15214_/B _15221_/A VGND VGND VPWR VPWR _15223_/B sky130_fd_sc_hd__or2_4
X_18006_ _18017_/A VGND VGND VPWR VPWR _18193_/A sky130_fd_sc_hd__buf_2
XFILLER_173_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16198_ _16190_/X VGND VGND VPWR VPWR _16198_/X sky130_fd_sc_hd__buf_2
XANTENNA__22471__A _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12383__C1 _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15149_ _15148_/Y _16432_/A _15417_/A _15120_/Y VGND VGND VPWR VPWR _15149_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24088__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21877__A1_N _22435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21087__A _21087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19957_ _19957_/A VGND VGND VPWR VPWR _21208_/B sky130_fd_sc_hd__inv_2
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24040__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22737__A2 _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_222_0_HCLK clkbuf_8_222_0_HCLK/A VGND VGND VPWR VPWR _24443_/CLK sky130_fd_sc_hd__clkbuf_1
X_18908_ _17503_/Y _11683_/X HWDATA[27] _11683_/X VGND VGND VPWR VPWR _18908_/X sky130_fd_sc_hd__a2bb2o_4
X_19888_ _19888_/A VGND VGND VPWR VPWR _19888_/Y sky130_fd_sc_hd__inv_2
XFILLER_228_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18839_ _24549_/Q _24128_/Q _16532_/Y _18819_/A VGND VGND VPWR VPWR _18839_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21815__A _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15624__B1 _15623_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21850_ _20506_/D _21849_/X _14450_/Y _17412_/X VGND VGND VPWR VPWR _21851_/D sky130_fd_sc_hd__o22a_4
XANTENNA__12438__B1 _12390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21534__B _23172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20801_ _20797_/X VGND VGND VPWR VPWR _20801_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21781_ _21777_/X _21780_/X _14744_/X VGND VGND VPWR VPWR _21781_/X sky130_fd_sc_hd__o21a_4
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17916__A2 _14764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22370__B1 _21773_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12336__A2_N _24832_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23520_ _23912_/CLK _23520_/D VGND VGND VPWR VPWR _13260_/B sky130_fd_sc_hd__dfxtp_4
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20732_ _13119_/B VGND VGND VPWR VPWR _20732_/Y sky130_fd_sc_hd__inv_2
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21550__A _21346_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23451_ _23452_/CLK _23451_/D VGND VGND VPWR VPWR _13424_/B sky130_fd_sc_hd__dfxtp_4
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20663_ _20663_/A VGND VGND VPWR VPWR _20663_/Y sky130_fd_sc_hd__inv_2
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22402_ _22395_/Y _22400_/X _22401_/X _24233_/Q _13807_/D VGND VGND VPWR VPWR _22402_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_195_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23382_ _23610_/CLK _23382_/D VGND VGND VPWR VPWR _20414_/A sky130_fd_sc_hd__dfxtp_4
X_20594_ _23948_/Q _18882_/B _20593_/Y _20543_/A VGND VGND VPWR VPWR _20595_/C sky130_fd_sc_hd__a211o_4
XANTENNA__12891__B _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24881__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25121_ _25109_/CLK _25121_/D HRESETn VGND VGND VPWR VPWR _25121_/Q sky130_fd_sc_hd__dfrtp_4
X_22333_ _22333_/A VGND VGND VPWR VPWR _22333_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11788__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21881__C1 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24199__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24810__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25052_ _25052_/CLK _14835_/X HRESETn VGND VGND VPWR VPWR _25052_/Q sky130_fd_sc_hd__dfrtp_4
X_22264_ _18296_/A _22260_/X _22263_/X VGND VGND VPWR VPWR _22264_/X sky130_fd_sc_hd__or3_4
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22381__A _22381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24128__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24003_ _24662_/CLK _24003_/D HRESETn VGND VGND VPWR VPWR _13110_/B sky130_fd_sc_hd__dfrtp_4
X_21215_ _21215_/A _21346_/A VGND VGND VPWR VPWR _21215_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_32_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_65_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22195_ _22195_/A _22195_/B _22195_/C _22194_/X VGND VGND VPWR VPWR _22195_/X sky130_fd_sc_hd__or4_4
X_21146_ _12087_/B _21144_/X _13482_/B _21145_/X VGND VGND VPWR VPWR _21146_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15863__B1 _15557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21077_ _21077_/A VGND VGND VPWR VPWR _21077_/X sky130_fd_sc_hd__buf_2
XFILLER_47_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20028_ _21467_/B _20025_/X _19984_/X _20025_/X VGND VGND VPWR VPWR _20028_/X sky130_fd_sc_hd__a2bb2o_4
X_24905_ _24903_/CLK _15604_/X HRESETn VGND VGND VPWR VPWR _24905_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_247_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12850_ _12588_/X _12825_/X VGND VGND VPWR VPWR _12851_/B sky130_fd_sc_hd__and2_4
XFILLER_246_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16132__A1_N _16131_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12429__B1 _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24836_ _24834_/CLK _15812_/X HRESETn VGND VGND VPWR VPWR _24836_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _25519_/Q _11860_/A _11802_/A VGND VGND VPWR VPWR _11801_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__23321__A1_N _17261_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _25373_/Q VGND VGND VPWR VPWR _12781_/Y sky130_fd_sc_hd__inv_2
X_24767_ _24766_/CLK _15950_/X HRESETn VGND VGND VPWR VPWR _22898_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _21979_/A _20322_/Y VGND VGND VPWR VPWR _21979_/X sky130_fd_sc_hd__and2_4
XFILLER_42_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14510_/X _14519_/X _14477_/A _14495_/Y VGND VGND VPWR VPWR _14520_/X sky130_fd_sc_hd__o22a_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13243__A _11950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _25534_/Q VGND VGND VPWR VPWR _11732_/Y sky130_fd_sc_hd__inv_2
X_23718_ _23691_/CLK _23718_/D VGND VGND VPWR VPWR _19491_/A sky130_fd_sc_hd__dfxtp_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24698_ _24753_/CLK _24698_/D HRESETn VGND VGND VPWR VPWR _24698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_214_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24969__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14450_/Y _14448_/X _14380_/X _14448_/X VGND VGND VPWR VPWR _25126_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _15984_/A _14178_/B _14365_/C _15984_/D VGND VGND VPWR VPWR _11664_/B sky130_fd_sc_hd__or4_4
X_23649_ _23644_/CLK _19697_/X VGND VGND VPWR VPWR _13233_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22113__B1 _21111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13434_/A _13402_/B _13402_/C VGND VGND VPWR VPWR _13402_/X sky130_fd_sc_hd__and3_4
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ _16317_/Y _24357_/Q _16317_/Y _24357_/Q VGND VGND VPWR VPWR _17170_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ _25149_/Q VGND VGND VPWR VPWR _14382_/Y sky130_fd_sc_hd__inv_2
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16121_ _16120_/Y _16116_/X _15953_/X _16116_/X VGND VGND VPWR VPWR _24698_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_114_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_229_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13333_ _13365_/A _13331_/X _13333_/C VGND VGND VPWR VPWR _13333_/X sky130_fd_sc_hd__and3_4
X_25319_ _25479_/CLK _13477_/X HRESETn VGND VGND VPWR VPWR _13475_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17540__B1 _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24551__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16052_ _16052_/A VGND VGND VPWR VPWR _16052_/Y sky130_fd_sc_hd__inv_2
X_13264_ _13289_/A VGND VGND VPWR VPWR _13264_/X sky130_fd_sc_hd__buf_2
X_15003_ _24454_/Q VGND VGND VPWR VPWR _15003_/Y sky130_fd_sc_hd__inv_2
X_12215_ _12174_/X _12186_/X _12215_/C _12215_/D VGND VGND VPWR VPWR _12261_/A sky130_fd_sc_hd__or4_4
XFILLER_142_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13195_ _13189_/A VGND VGND VPWR VPWR _13289_/A sky130_fd_sc_hd__buf_2
XANTENNA__19293__B1 _19203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14802__A _20628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19811_ _19809_/Y _19806_/X _19810_/X _19806_/X VGND VGND VPWR VPWR _19811_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12146_ _18372_/D VGND VGND VPWR VPWR _12147_/A sky130_fd_sc_hd__buf_2
XFILLER_111_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19742_ _23633_/Q VGND VGND VPWR VPWR _19742_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19045__B1 _18998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12077_ _12074_/Y _12072_/X _12076_/X _12072_/X VGND VGND VPWR VPWR _25480_/D sky130_fd_sc_hd__a2bb2o_4
X_16954_ _21014_/B _16952_/X _16953_/Y VGND VGND VPWR VPWR _16954_/X sky130_fd_sc_hd__o21a_4
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12322__A _24822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_238_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15905_ _24784_/Q _13527_/B VGND VGND VPWR VPWR _15905_/X sky130_fd_sc_hd__or2_4
XANTENNA__21635__A _22380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19673_ _19672_/Y VGND VGND VPWR VPWR _19673_/X sky130_fd_sc_hd__buf_2
X_16885_ _19827_/A VGND VGND VPWR VPWR _16885_/X sky130_fd_sc_hd__buf_2
XFILLER_92_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15606__B1 _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18624_ _24539_/Q _24150_/Q _16559_/Y _18677_/A VGND VGND VPWR VPWR _18627_/C sky130_fd_sc_hd__o22a_4
XFILLER_92_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_52_0_HCLK clkbuf_7_26_0_HCLK/X VGND VGND VPWR VPWR _25524_/CLK sky130_fd_sc_hd__clkbuf_1
X_15836_ _15771_/B _15836_/B VGND VGND VPWR VPWR _15836_/X sky130_fd_sc_hd__or2_4
XFILLER_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16448__B _16721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18555_ _24171_/Q _18555_/B VGND VGND VPWR VPWR _18557_/B sky130_fd_sc_hd__or2_4
X_12979_ _13074_/A _13073_/A _13072_/A _12979_/D VGND VGND VPWR VPWR _12984_/A sky130_fd_sc_hd__or4_4
X_15767_ _12550_/Y _15759_/X _14479_/X _15713_/X VGND VGND VPWR VPWR _15767_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17506_ _17506_/A _17501_/X _17504_/X _17505_/X VGND VGND VPWR VPWR _17506_/X sky130_fd_sc_hd__or4_4
XANTENNA__13153__A _13168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24952__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14718_ _14718_/A VGND VGND VPWR VPWR _14718_/Y sky130_fd_sc_hd__inv_2
X_18486_ _24189_/Q _18484_/Y VGND VGND VPWR VPWR _18487_/C sky130_fd_sc_hd__nand2_4
X_15698_ _15698_/A VGND VGND VPWR VPWR _15836_/B sky130_fd_sc_hd__buf_2
XANTENNA__22466__A _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17437_ _17436_/X VGND VGND VPWR VPWR _17438_/B sky130_fd_sc_hd__buf_2
X_14649_ _25073_/Q VGND VGND VPWR VPWR _19002_/B sky130_fd_sc_hd__buf_2
XANTENNA__16464__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24639__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22655__A1 _16539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17368_ _17346_/D VGND VGND VPWR VPWR _17369_/B sky130_fd_sc_hd__inv_2
XANTENNA__22655__B2 _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16183__B _16540_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19107_ _19105_/Y _19101_/X _19106_/X _19101_/X VGND VGND VPWR VPWR _23854_/D sky130_fd_sc_hd__a2bb2o_4
X_16319_ _16344_/A VGND VGND VPWR VPWR _16319_/X sky130_fd_sc_hd__buf_2
X_17299_ _17230_/X _17299_/B _17299_/C VGND VGND VPWR VPWR _24364_/D sky130_fd_sc_hd__and3_4
XANTENNA__17531__B1 _25525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24292__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19038_ _19037_/Y _19033_/X _18965_/X _19033_/X VGND VGND VPWR VPWR _19038_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22407__A1 _25527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24221__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22958__A2 _22718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19284__B1 _19282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23080__A1 _24740_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_19_0_HCLK clkbuf_4_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_19_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21000_ _21000_/A _21000_/B VGND VGND VPWR VPWR _21000_/X sky130_fd_sc_hd__and2_4
XFILLER_130_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25498__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19036__B1 _18942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15246__C _15246_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22951_ _21421_/A _22949_/X _22831_/X _22950_/X VGND VGND VPWR VPWR _22952_/A sky130_fd_sc_hd__o22a_4
XFILLER_56_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21902_ _21902_/A _20145_/Y VGND VGND VPWR VPWR _21902_/X sky130_fd_sc_hd__or2_4
XANTENNA__15543__A _14366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22882_ _23062_/A _22882_/B VGND VGND VPWR VPWR _22882_/Y sky130_fd_sc_hd__nor2_4
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25080__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24621_ _24623_/CLK _24621_/D HRESETn VGND VGND VPWR VPWR _24621_/Q sky130_fd_sc_hd__dfrtp_4
X_21833_ _21325_/X VGND VGND VPWR VPWR _21833_/X sky130_fd_sc_hd__buf_2
XFILLER_24_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24552_ _24555_/CLK _16526_/X HRESETn VGND VGND VPWR VPWR _24552_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21764_ _21764_/A _21762_/X _21763_/X VGND VGND VPWR VPWR _21764_/X sky130_fd_sc_hd__and3_4
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23503_ _23808_/CLK _23503_/D VGND VGND VPWR VPWR _23503_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20715_ _20715_/A VGND VGND VPWR VPWR _20715_/Y sky130_fd_sc_hd__inv_2
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24483_ _24594_/CLK _24483_/D HRESETn VGND VGND VPWR VPWR _16706_/A sky130_fd_sc_hd__dfrtp_4
X_21695_ _21695_/A VGND VGND VPWR VPWR _21695_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23434_ _23675_/CLK _23434_/D VGND VGND VPWR VPWR _23434_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20646_ _14229_/Y _20638_/X _20629_/X _20645_/X VGND VGND VPWR VPWR _20646_/X sky130_fd_sc_hd__a211o_4
XFILLER_11_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24309__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23365_ _21012_/X VGND VGND VPWR VPWR IRQ[21] sky130_fd_sc_hd__buf_2
XFILLER_176_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20577_ _20580_/B _20576_/Y _20572_/X VGND VGND VPWR VPWR _20577_/X sky130_fd_sc_hd__and3_4
XFILLER_20_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25104_ _25146_/CLK _14518_/X HRESETn VGND VGND VPWR VPWR _25104_/Q sky130_fd_sc_hd__dfrtp_4
X_22316_ _14096_/A _17411_/X _20601_/A _22181_/B VGND VGND VPWR VPWR _22316_/X sky130_fd_sc_hd__a2bb2o_4
X_23296_ _23169_/A _23296_/B VGND VGND VPWR VPWR _23296_/Y sky130_fd_sc_hd__nor2_4
X_25035_ _25035_/CLK _15183_/X HRESETn VGND VGND VPWR VPWR _14886_/A sky130_fd_sc_hd__dfrtp_4
X_22247_ _22255_/A _22247_/B VGND VGND VPWR VPWR _22247_/X sky130_fd_sc_hd__or2_4
XFILLER_152_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12898__B1 _12862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12000_ _25315_/Q VGND VGND VPWR VPWR _12000_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16089__B1 _15554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22178_ _12097_/Y _12086_/A _18376_/Y _12057_/A VGND VGND VPWR VPWR _22178_/X sky130_fd_sc_hd__o22a_4
XFILLER_120_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21129_ _21040_/X _21126_/X _21127_/X _21128_/Y VGND VGND VPWR VPWR _21129_/X sky130_fd_sc_hd__a211o_4
XANTENNA__13238__A _13421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23944__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13951_ _13957_/A _13943_/X _13950_/X VGND VGND VPWR VPWR _13952_/B sky130_fd_sc_hd__o21ai_4
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12902_ _12766_/Y _12906_/B _12901_/Y VGND VGND VPWR VPWR _12902_/X sky130_fd_sc_hd__o21a_4
XFILLER_86_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_39_0_HCLK clkbuf_7_39_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_79_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13882_ _13902_/A _14232_/C _13924_/A _15421_/B VGND VGND VPWR VPWR _13883_/A sky130_fd_sc_hd__or4_4
X_16670_ _16670_/A VGND VGND VPWR VPWR _16670_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12833_ _12816_/Y _12775_/Y _12833_/C VGND VGND VPWR VPWR _12833_/X sky130_fd_sc_hd__or3_4
X_15621_ _24898_/Q VGND VGND VPWR VPWR _15621_/Y sky130_fd_sc_hd__inv_2
X_24819_ _24819_/CLK _15837_/X HRESETn VGND VGND VPWR VPWR _24819_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22334__B1 _21556_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18340_ _18900_/A _18326_/B _17473_/Y VGND VGND VPWR VPWR _18341_/A sky130_fd_sc_hd__o21a_4
X_12764_ _12762_/A _22420_/A _12762_/Y _12763_/Y VGND VGND VPWR VPWR _12765_/D sky130_fd_sc_hd__o22a_4
X_15552_ _15608_/A VGND VGND VPWR VPWR _15553_/A sky130_fd_sc_hd__buf_2
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16013__B1 _15939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ HWDATA[19] VGND VGND VPWR VPWR _11715_/X sky130_fd_sc_hd__buf_2
X_14503_ _14490_/B _14500_/X _14501_/Y _14502_/X VGND VGND VPWR VPWR _14503_/X sky130_fd_sc_hd__o22a_4
XFILLER_230_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _15483_/A VGND VGND VPWR VPWR _24070_/D sky130_fd_sc_hd__buf_2
X_18271_ _13783_/D _18256_/X _16267_/X _23348_/A _18264_/X VGND VGND VPWR VPWR _24221_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_15_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12695_ _12704_/A _12707_/B VGND VGND VPWR VPWR _12696_/B sky130_fd_sc_hd__or2_4
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24732__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _16352_/Y _17241_/A _24613_/Q _17203_/X VGND VGND VPWR VPWR _17226_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_202_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14434_ _14433_/Y _14431_/X _14380_/X _14431_/X VGND VGND VPWR VPWR _14434_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ _15984_/A _14365_/B _14365_/C _14365_/D VGND VGND VPWR VPWR _21343_/A sky130_fd_sc_hd__or4_4
X_17153_ _17125_/A _17153_/B VGND VGND VPWR VPWR _17153_/Y sky130_fd_sc_hd__nand2_4
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13316_ _13445_/A _19749_/A VGND VGND VPWR VPWR _13318_/B sky130_fd_sc_hd__or2_4
X_16104_ _16111_/A VGND VGND VPWR VPWR _16104_/X sky130_fd_sc_hd__buf_2
X_17084_ _17045_/D _17062_/X _17006_/Y VGND VGND VPWR VPWR _17084_/X sky130_fd_sc_hd__o21a_4
XFILLER_7_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14296_ _14296_/A VGND VGND VPWR VPWR _14296_/X sky130_fd_sc_hd__buf_2
XFILLER_115_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13247_ _13247_/A VGND VGND VPWR VPWR _13390_/A sky130_fd_sc_hd__buf_2
X_16035_ _16035_/A VGND VGND VPWR VPWR _16035_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13178_ _13175_/A _13178_/B VGND VGND VPWR VPWR _13179_/C sky130_fd_sc_hd__or2_4
XFILLER_111_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18939__A _18947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12129_ _12129_/A VGND VGND VPWR VPWR _12129_/Y sky130_fd_sc_hd__inv_2
X_17986_ _17985_/X _17986_/B VGND VGND VPWR VPWR _17986_/X sky130_fd_sc_hd__or2_4
XANTENNA__25520__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19725_ _19725_/A VGND VGND VPWR VPWR _19725_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16039__A1_N _16037_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21365__A _21365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16937_ _16154_/Y _24262_/Q _23225_/A _16945_/A VGND VGND VPWR VPWR _16937_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16459__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19656_ _19656_/A VGND VGND VPWR VPWR _19656_/Y sky130_fd_sc_hd__inv_2
X_16868_ _16867_/X VGND VGND VPWR VPWR _16868_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18607_ _18600_/X _18607_/B _18607_/C _18607_/D VGND VGND VPWR VPWR _18638_/A sky130_fd_sc_hd__or4_4
X_15819_ _15818_/X _15813_/X _16240_/A _24831_/Q _15786_/X VGND VGND VPWR VPWR _15819_/X
+ sky130_fd_sc_hd__a32o_4
X_19587_ _11780_/A VGND VGND VPWR VPWR _19587_/X sky130_fd_sc_hd__buf_2
XFILLER_241_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16799_ _16799_/A VGND VGND VPWR VPWR _16799_/X sky130_fd_sc_hd__buf_2
XFILLER_203_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18538_ _18466_/B _18538_/B VGND VGND VPWR VPWR _18538_/X sky130_fd_sc_hd__or2_4
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22196__A _22196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18469_ _24171_/Q VGND VGND VPWR VPWR _18556_/A sky130_fd_sc_hd__inv_2
XFILLER_194_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14707__A _22205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24473__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20500_ _13962_/A _20500_/B VGND VGND VPWR VPWR _20501_/B sky130_fd_sc_hd__nor2_4
XFILLER_178_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21480_ _21809_/A _21480_/B VGND VGND VPWR VPWR _21483_/B sky130_fd_sc_hd__or2_4
XFILLER_165_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24402__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20431_ _20430_/X VGND VGND VPWR VPWR _23926_/D sky130_fd_sc_hd__buf_2
XFILLER_174_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23150_ _23280_/A _23150_/B VGND VGND VPWR VPWR _23160_/C sky130_fd_sc_hd__and2_4
XFILLER_180_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20362_ _20349_/Y VGND VGND VPWR VPWR _20362_/X sky130_fd_sc_hd__buf_2
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14869__A1 _14863_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22101_ _22708_/A _22097_/X _22101_/C VGND VGND VPWR VPWR _22101_/X sky130_fd_sc_hd__and3_4
X_23081_ _22141_/X _23081_/B _23080_/X VGND VGND VPWR VPWR _23081_/X sky130_fd_sc_hd__and3_4
X_20293_ _20287_/Y VGND VGND VPWR VPWR _20293_/X sky130_fd_sc_hd__buf_2
X_22032_ _22028_/X _22031_/X _21686_/X VGND VGND VPWR VPWR _22032_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_103_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19009__B1 _18981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16491__B1 _16400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23983_ _25050_/CLK _23983_/D HRESETn VGND VGND VPWR VPWR _17392_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_228_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22934_ _24465_/Q _22431_/X _22891_/X VGND VGND VPWR VPWR _22934_/X sky130_fd_sc_hd__o21a_4
XFILLER_17_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16243__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22865_ _21127_/X VGND VGND VPWR VPWR _22865_/X sky130_fd_sc_hd__buf_2
XFILLER_83_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22316__B1 _20601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21816_ _21657_/A _21816_/B VGND VGND VPWR VPWR _21816_/X sky130_fd_sc_hd__or2_4
X_24604_ _25005_/CLK _24604_/D HRESETn VGND VGND VPWR VPWR _24604_/Q sky130_fd_sc_hd__dfrtp_4
X_22796_ _23328_/A _22796_/B VGND VGND VPWR VPWR _22796_/Y sky130_fd_sc_hd__nor2_4
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24535_ _24573_/CLK _24535_/D HRESETn VGND VGND VPWR VPWR _16569_/A sky130_fd_sc_hd__dfrtp_4
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21747_ _21597_/A _21745_/X _21121_/A _21746_/X VGND VGND VPWR VPWR _21747_/X sky130_fd_sc_hd__o22a_4
XFILLER_52_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13521__A _14262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12480_ _12480_/A _12480_/B _12479_/Y VGND VGND VPWR VPWR _12480_/X sky130_fd_sc_hd__and3_4
X_24466_ _24443_/CLK _16747_/X HRESETn VGND VGND VPWR VPWR _15047_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_169_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21678_ _22021_/A _21676_/X _21678_/C VGND VGND VPWR VPWR _21678_/X sky130_fd_sc_hd__and3_4
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24143__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23417_ _23415_/CLK _23417_/D VGND VGND VPWR VPWR _20326_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20629_ _20629_/A VGND VGND VPWR VPWR _20629_/X sky130_fd_sc_hd__buf_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24397_ _24377_/CLK _17080_/X HRESETn VGND VGND VPWR VPWR _24397_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14150_ _14135_/X _14149_/Y _25135_/Q _14100_/X VGND VGND VPWR VPWR _25215_/D sky130_fd_sc_hd__a2bb2o_4
X_23348_ _23348_/A _23347_/X VGND VGND VPWR VPWR _23348_/X sky130_fd_sc_hd__and2_4
XFILLER_165_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13101_ _13068_/D VGND VGND VPWR VPWR _13101_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081_ _14012_/A _20453_/C _14058_/X _14022_/B _14049_/B VGND VGND VPWR VPWR _25227_/D
+ sky130_fd_sc_hd__a32o_4
X_23279_ _21868_/X _23278_/X _22477_/X _24885_/Q _21871_/X VGND VGND VPWR VPWR _23280_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25349__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13032_ _12977_/X _13032_/B VGND VGND VPWR VPWR _13032_/X sky130_fd_sc_hd__or2_4
X_25018_ _25015_/CLK _25018_/D HRESETn VGND VGND VPWR VPWR _15026_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__15809__B1 _11721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17840_ _17602_/B _17811_/D VGND VGND VPWR VPWR _17841_/B sky130_fd_sc_hd__or2_4
XFILLER_154_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17771_ _23320_/A _17769_/Y VGND VGND VPWR VPWR _17772_/C sky130_fd_sc_hd__nand2_4
X_14983_ _15219_/A _24464_/Q _15219_/A _24464_/Q VGND VGND VPWR VPWR _14983_/X sky130_fd_sc_hd__a2bb2o_4
X_19510_ _23711_/Q VGND VGND VPWR VPWR _21948_/B sky130_fd_sc_hd__inv_2
X_16722_ _15323_/A _16721_/X _16716_/X _16721_/X VGND VGND VPWR VPWR _16722_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15183__A _15165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13934_ _24975_/Q _13934_/B _13934_/C VGND VGND VPWR VPWR _13934_/X sky130_fd_sc_hd__or3_4
XANTENNA__19420__B1 _19395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16234__B1 _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24984__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19441_ _19439_/Y _19435_/X _19395_/X _19440_/X VGND VGND VPWR VPWR _19441_/X sky130_fd_sc_hd__a2bb2o_4
X_16653_ _16652_/Y _16648_/X _16382_/X _16648_/X VGND VGND VPWR VPWR _16653_/X sky130_fd_sc_hd__a2bb2o_4
X_13865_ _21723_/A _13849_/X _21559_/A _13844_/X VGND VGND VPWR VPWR _13865_/X sky130_fd_sc_hd__o22a_4
XFILLER_234_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24913__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15604_ _15603_/Y _15601_/X _11743_/X _15601_/X VGND VGND VPWR VPWR _15604_/X sky130_fd_sc_hd__a2bb2o_4
X_12816_ _25371_/Q VGND VGND VPWR VPWR _12816_/Y sky130_fd_sc_hd__inv_2
X_19372_ _19372_/A VGND VGND VPWR VPWR _19372_/X sky130_fd_sc_hd__buf_2
X_16584_ _24529_/Q VGND VGND VPWR VPWR _16584_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13796_ _25271_/Q VGND VGND VPWR VPWR _13796_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_126_0_HCLK clkbuf_7_63_0_HCLK/X VGND VGND VPWR VPWR _24508_/CLK sky130_fd_sc_hd__clkbuf_1
X_18323_ _21822_/A _18322_/Y _17894_/Y VGND VGND VPWR VPWR _24211_/D sky130_fd_sc_hd__o21a_4
X_15535_ _13581_/A VGND VGND VPWR VPWR _15535_/Y sky130_fd_sc_hd__inv_2
X_12747_ _23187_/A VGND VGND VPWR VPWR _12747_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_189_0_HCLK clkbuf_7_94_0_HCLK/X VGND VGND VPWR VPWR _25226_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15032__A2_N _24453_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18254_ _11824_/Y _18252_/X _17421_/X _18252_/X VGND VGND VPWR VPWR _24231_/D sky130_fd_sc_hd__a2bb2o_4
X_12678_ _12555_/Y _12662_/B _12627_/X _12675_/Y VGND VGND VPWR VPWR _12678_/X sky130_fd_sc_hd__a211o_4
X_15466_ _14380_/A VGND VGND VPWR VPWR _15466_/X sky130_fd_sc_hd__buf_2
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14246__B _14212_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17205_ _24613_/Q _17203_/X _24617_/Q _17346_/C VGND VGND VPWR VPWR _17208_/B sky130_fd_sc_hd__a2bb2o_4
X_14417_ _14417_/A VGND VGND VPWR VPWR _14417_/Y sky130_fd_sc_hd__inv_2
X_18185_ _18053_/A _23772_/Q VGND VGND VPWR VPWR _18185_/X sky130_fd_sc_hd__or2_4
XFILLER_156_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15397_ _15294_/B _15400_/B VGND VGND VPWR VPWR _15398_/C sky130_fd_sc_hd__nand2_4
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17136_ _17142_/A _17132_/X _17136_/C VGND VGND VPWR VPWR _17136_/X sky130_fd_sc_hd__and3_4
X_14348_ _25160_/Q _14340_/X _25159_/Q _14345_/X VGND VGND VPWR VPWR _14348_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11782__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14279_ _13513_/B _12013_/B _13509_/X VGND VGND VPWR VPWR _14283_/B sky130_fd_sc_hd__or3_4
X_17067_ _17069_/B VGND VGND VPWR VPWR _17072_/B sky130_fd_sc_hd__inv_2
XFILLER_144_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14262__A _14262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16018_ _24737_/Q VGND VGND VPWR VPWR _16018_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25019__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16473__B1 _16295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15815__A3 _15741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17969_ _13597_/A VGND VGND VPWR VPWR _18027_/A sky130_fd_sc_hd__buf_2
XANTENNA__22546__B1 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19708_ _11785_/A VGND VGND VPWR VPWR _19708_/X sky130_fd_sc_hd__buf_2
X_20980_ scl_oen_o_S4 _20979_/Y VGND VGND VPWR VPWR _20980_/X sky130_fd_sc_hd__and2_4
XFILLER_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22919__A _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19639_ _19638_/Y _19634_/X _19587_/X _19634_/X VGND VGND VPWR VPWR _23670_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16531__A1_N _16530_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_22_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16917__A _16917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24654__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22638__B _22638_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_85_0_HCLK clkbuf_7_85_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_85_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22650_ _22618_/X _22650_/B _22650_/C _22649_/Y VGND VGND VPWR VPWR HRDATA[12] sky130_fd_sc_hd__or4_4
XFILLER_241_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21601_ _21601_/A _21601_/B _21601_/C _21600_/X VGND VGND VPWR VPWR _21601_/X sky130_fd_sc_hd__or4_4
XFILLER_241_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22581_ _22539_/A _22581_/B _22581_/C VGND VGND VPWR VPWR _22581_/X sky130_fd_sc_hd__and3_4
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24320_ _24315_/CLK _24320_/D HRESETn VGND VGND VPWR VPWR _17516_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21532_ _21531_/X VGND VGND VPWR VPWR _21532_/X sky130_fd_sc_hd__buf_2
XFILLER_166_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22654__A _24761_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24251_ _23747_/CLK _17929_/X HRESETn VGND VGND VPWR VPWR _24251_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_239_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21463_ _21463_/A VGND VGND VPWR VPWR _21661_/A sky130_fd_sc_hd__buf_2
XFILLER_166_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17748__A _24262_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23202_ _23120_/X _23200_/X _23123_/X _23201_/X VGND VGND VPWR VPWR _23203_/B sky130_fd_sc_hd__o22a_4
X_20414_ _20414_/A VGND VGND VPWR VPWR _22070_/B sky130_fd_sc_hd__inv_2
XANTENNA__21285__B1 _21284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24182_ _24675_/CLK _18516_/X HRESETn VGND VGND VPWR VPWR _18411_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_147_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21394_ _21385_/X _19088_/Y VGND VGND VPWR VPWR _21395_/C sky130_fd_sc_hd__or2_4
XFILLER_135_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23133_ _23178_/A VGND VGND VPWR VPWR _23133_/X sky130_fd_sc_hd__buf_2
XANTENNA__15268__A _25013_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20345_ _20345_/A VGND VGND VPWR VPWR _20345_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19963__A _19962_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23064_ _23064_/A _23063_/X VGND VGND VPWR VPWR _23064_/X sky130_fd_sc_hd__or2_4
XFILLER_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20276_ _20276_/A VGND VGND VPWR VPWR _21792_/B sky130_fd_sc_hd__inv_2
XFILLER_115_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22015_ _22015_/A VGND VGND VPWR VPWR _22016_/A sky130_fd_sc_hd__buf_2
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20260__B2 _20243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11980_ _24095_/Q _11979_/X VGND VGND VPWR VPWR _11981_/A sky130_fd_sc_hd__and2_4
X_23966_ _25243_/CLK _23966_/D HRESETn VGND VGND VPWR VPWR _23966_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16216__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22829__A _22829_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22917_ _21022_/A VGND VGND VPWR VPWR _22917_/X sky130_fd_sc_hd__buf_2
XFILLER_72_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23897_ _23827_/CLK _23897_/D VGND VGND VPWR VPWR _18007_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_232_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22548__B _16368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24395__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15731__A _15713_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19203__A _19360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18745__C _18745_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13650_ _24048_/Q _13649_/X _13650_/C _20889_/A VGND VGND VPWR VPWR _13650_/X sky130_fd_sc_hd__or4_4
X_22848_ _23094_/A _22848_/B VGND VGND VPWR VPWR _22848_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__20349__A _20348_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _25411_/Q VGND VGND VPWR VPWR _12697_/A sky130_fd_sc_hd__inv_2
X_13581_ _13581_/A _13581_/B VGND VGND VPWR VPWR _19522_/A sky130_fd_sc_hd__or2_4
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ _11681_/B _22778_/X _22495_/X _25536_/Q _15983_/X VGND VGND VPWR VPWR _22779_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21171__C _21327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12532_ _12532_/A _12532_/B _12528_/X _12532_/D VGND VGND VPWR VPWR _12532_/X sky130_fd_sc_hd__or4_4
X_15320_ _15082_/Y _15320_/B _15326_/A _15320_/D VGND VGND VPWR VPWR _15320_/X sky130_fd_sc_hd__or4_4
X_24518_ _24520_/CLK _24518_/D HRESETn VGND VGND VPWR VPWR _24518_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25498_ _25499_/CLK _11968_/X HRESETn VGND VGND VPWR VPWR _11932_/C sky130_fd_sc_hd__dfrtp_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22564__A _22564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12463_ _12266_/A _12461_/A VGND VGND VPWR VPWR _12463_/X sky130_fd_sc_hd__or2_4
X_15251_ _15251_/A _15254_/A _15254_/B VGND VGND VPWR VPWR _15251_/X sky130_fd_sc_hd__or3_4
XFILLER_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24449_ _24419_/CLK _16784_/X HRESETn VGND VGND VPWR VPWR _16781_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14202_ _14201_/Y _14199_/X _13521_/X _14190_/A VGND VGND VPWR VPWR _14202_/X sky130_fd_sc_hd__a2bb2o_4
X_15182_ _15182_/A _15180_/A VGND VGND VPWR VPWR _15183_/C sky130_fd_sc_hd__or2_4
XANTENNA__22473__C1 _22472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12394_ _12396_/B VGND VGND VPWR VPWR _12400_/B sky130_fd_sc_hd__inv_2
X_14133_ _14113_/X VGND VGND VPWR VPWR _14133_/X sky130_fd_sc_hd__buf_2
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23017__A1 _12240_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19990_ _19989_/X VGND VGND VPWR VPWR _19990_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14064_ _13986_/X _14054_/X _14046_/X _13978_/X _14055_/X VGND VGND VPWR VPWR _14064_/X
+ sky130_fd_sc_hd__a32o_4
X_18941_ _23911_/Q VGND VGND VPWR VPWR _18941_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18489__A _18823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13015_ _13015_/A VGND VGND VPWR VPWR _13015_/Y sky130_fd_sc_hd__inv_2
XFILLER_239_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18872_ _18872_/A _20544_/A VGND VGND VPWR VPWR _18872_/X sky130_fd_sc_hd__or2_4
XFILLER_67_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16455__B1 _15545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17823_ _16911_/Y _17827_/B _17822_/Y VGND VGND VPWR VPWR _17823_/X sky130_fd_sc_hd__o21a_4
XFILLER_79_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17754_ _16908_/Y _16889_/Y _17750_/X _17753_/X VGND VGND VPWR VPWR _17811_/D sky130_fd_sc_hd__or4_4
X_14966_ _14966_/A VGND VGND VPWR VPWR _14966_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16705_ _16703_/Y _16704_/X _16525_/X _16704_/X VGND VGND VPWR VPWR _16705_/X sky130_fd_sc_hd__a2bb2o_4
X_13917_ _13942_/C _13917_/B VGND VGND VPWR VPWR _13947_/C sky130_fd_sc_hd__or2_4
X_17685_ _17669_/B _17685_/B _17688_/C VGND VGND VPWR VPWR _17685_/X sky130_fd_sc_hd__and3_4
XFILLER_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14897_ _15026_/A _14895_/Y _15066_/A _24440_/Q VGND VGND VPWR VPWR _14897_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19424_ _19423_/Y _19419_/X _19377_/X _19419_/X VGND VGND VPWR VPWR _23742_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_223_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15641__A _15644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16636_ _13728_/B _16635_/X _16631_/X VGND VGND VPWR VPWR _24511_/D sky130_fd_sc_hd__o21a_4
XFILLER_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13848_ _20476_/A _13846_/X _13841_/X _13847_/Y VGND VGND VPWR VPWR _13848_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24065__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19355_ _18135_/B VGND VGND VPWR VPWR _19355_/Y sky130_fd_sc_hd__inv_2
X_16567_ _16548_/A VGND VGND VPWR VPWR _16567_/X sky130_fd_sc_hd__buf_2
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13779_ _19570_/A _14243_/A VGND VGND VPWR VPWR _13779_/X sky130_fd_sc_hd__or2_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18306_ _18306_/A VGND VGND VPWR VPWR _18306_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15518_ _15518_/A VGND VGND VPWR VPWR _15518_/Y sky130_fd_sc_hd__inv_2
X_19286_ _19285_/Y _19283_/X _19194_/X _19283_/X VGND VGND VPWR VPWR _23791_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16498_ _24562_/Q VGND VGND VPWR VPWR _16498_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22474__A _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18237_ _22735_/A _18236_/X _15739_/X _18236_/X VGND VGND VPWR VPWR _18237_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15449_ _24074_/Q _15444_/X _15436_/Y _13935_/A _15447_/X VGND VGND VPWR VPWR _15449_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_148_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23256__A1 _12769_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18168_ _18104_/A _18168_/B VGND VGND VPWR VPWR _18168_/X sky130_fd_sc_hd__or2_4
XANTENNA__14941__B1 _25013_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17119_ _24386_/Q _17118_/Y VGND VGND VPWR VPWR _17119_/X sky130_fd_sc_hd__or2_4
XFILLER_117_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18099_ _18099_/A _18099_/B _18099_/C VGND VGND VPWR VPWR _18100_/C sky130_fd_sc_hd__or3_4
XFILLER_171_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20130_ _23492_/Q VGND VGND VPWR VPWR _21411_/B sky130_fd_sc_hd__inv_2
XFILLER_143_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20061_ _11785_/A VGND VGND VPWR VPWR _20061_/X sky130_fd_sc_hd__buf_2
XFILLER_225_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24835__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23820_ _23827_/CLK _23820_/D VGND VGND VPWR VPWR _18193_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23751_ _23785_/CLK _19399_/X VGND VGND VPWR VPWR _18073_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_242_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20963_ _11977_/A _13507_/Y VGND VGND VPWR VPWR _24091_/D sky130_fd_sc_hd__nor2_4
XFILLER_241_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21742__A1 _16613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22702_ _24460_/Q _21843_/B _21741_/B VGND VGND VPWR VPWR _22702_/X sky130_fd_sc_hd__and3_4
XPHY_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23682_ _23559_/CLK _23682_/D VGND VGND VPWR VPWR _23682_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ _20921_/C VGND VGND VPWR VPWR _20894_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22633_ _24760_/Q _22487_/X VGND VGND VPWR VPWR _22633_/X sky130_fd_sc_hd__or2_4
X_25421_ _24872_/CLK _25421_/D HRESETn VGND VGND VPWR VPWR _12575_/A sky130_fd_sc_hd__dfrtp_4
X_25352_ _25344_/CLK _13050_/X HRESETn VGND VGND VPWR VPWR _12344_/A sky130_fd_sc_hd__dfrtp_4
X_22564_ _22564_/A _21101_/A VGND VGND VPWR VPWR _22564_/X sky130_fd_sc_hd__or2_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_172_0_HCLK clkbuf_7_86_0_HCLK/X VGND VGND VPWR VPWR _23827_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_167_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21515_ _21955_/A VGND VGND VPWR VPWR _21515_/Y sky130_fd_sc_hd__inv_2
X_24303_ _23411_/CLK _17663_/Y HRESETn VGND VGND VPWR VPWR _24303_/Q sky130_fd_sc_hd__dfrtp_4
X_25283_ _24227_/CLK _25283_/D HRESETn VGND VGND VPWR VPWR _11840_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22495_ _21436_/X VGND VGND VPWR VPWR _22495_/X sky130_fd_sc_hd__buf_2
XFILLER_182_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16382__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_29_0_HCLK clkbuf_8_29_0_HCLK/A VGND VGND VPWR VPWR _24315_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_108_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24234_ _24236_/CLK _24234_/D HRESETn VGND VGND VPWR VPWR _24234_/Q sky130_fd_sc_hd__dfrtp_4
X_21446_ _21019_/X VGND VGND VPWR VPWR _21446_/X sky130_fd_sc_hd__buf_2
X_24165_ _24650_/CLK _18578_/X HRESETn VGND VGND VPWR VPWR _24165_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21377_ _13780_/Y _19523_/Y _19572_/A VGND VGND VPWR VPWR _21377_/X sky130_fd_sc_hd__or3_4
XANTENNA__22470__A2 _21596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23116_ _12172_/Y _22984_/X _24283_/Q _22914_/X VGND VGND VPWR VPWR _23118_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20328_ _20328_/A VGND VGND VPWR VPWR _20328_/Y sky130_fd_sc_hd__inv_2
X_24096_ _23916_/CLK _24096_/D HRESETn VGND VGND VPWR VPWR _12001_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23047_ _23044_/X _23045_/X _23046_/X _16014_/A _22865_/X VGND VGND VPWR VPWR _23047_/X
+ sky130_fd_sc_hd__a32o_4
X_20259_ _23443_/Q VGND VGND VPWR VPWR _21266_/B sky130_fd_sc_hd__inv_2
XANTENNA__16437__B1 _16358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21166__C _21327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24576__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14820_ _14838_/A VGND VGND VPWR VPWR _14820_/X sky130_fd_sc_hd__buf_2
XFILLER_236_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12150__A _18372_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24998_ _24953_/CLK _24998_/D HRESETn VGND VGND VPWR VPWR _24998_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22559__A _21127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23183__B1 _23167_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24505__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21463__A _21463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14751_ _21239_/A VGND VGND VPWR VPWR _22202_/A sky130_fd_sc_hd__buf_2
X_11963_ _11956_/X _11962_/X VGND VGND VPWR VPWR _11963_/X sky130_fd_sc_hd__and2_4
X_23949_ _25211_/CLK _20598_/Y HRESETn VGND VGND VPWR VPWR _23949_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_245_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13702_ _13677_/B _13694_/X _13699_/Y _13701_/X _25290_/Q VGND VGND VPWR VPWR _13702_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_189_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17470_ _18911_/B _17462_/X VGND VGND VPWR VPWR _17470_/Y sky130_fd_sc_hd__nor2_4
X_11894_ _19964_/A VGND VGND VPWR VPWR _19600_/A sky130_fd_sc_hd__buf_2
X_14682_ _22219_/A VGND VGND VPWR VPWR _21764_/A sky130_fd_sc_hd__buf_2
XFILLER_189_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20079__A _20067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16276__B _15986_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16421_ _15081_/Y _16418_/X _16420_/X _16418_/X VGND VGND VPWR VPWR _24590_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13633_ _25300_/Q _14294_/A _13632_/X VGND VGND VPWR VPWR _13633_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_189_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19140_ _19140_/A VGND VGND VPWR VPWR _19140_/Y sky130_fd_sc_hd__inv_2
X_16352_ _24615_/Q VGND VGND VPWR VPWR _16352_/Y sky130_fd_sc_hd__inv_2
X_13564_ _13562_/A _13563_/A _13562_/Y _13563_/Y VGND VGND VPWR VPWR _13564_/X sky130_fd_sc_hd__o22a_4
XFILLER_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22294__A _22451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15303_ _15082_/Y _15320_/B VGND VGND VPWR VPWR _15303_/X sky130_fd_sc_hd__or2_4
XFILLER_200_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12515_ _12515_/A VGND VGND VPWR VPWR _12515_/Y sky130_fd_sc_hd__inv_2
X_19071_ _23866_/Q VGND VGND VPWR VPWR _19071_/Y sky130_fd_sc_hd__inv_2
X_13495_ _11986_/Y _13494_/X _11775_/X _13494_/X VGND VGND VPWR VPWR _13495_/X sky130_fd_sc_hd__a2bb2o_4
X_16283_ _23253_/A VGND VGND VPWR VPWR _16283_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25364__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18022_ _18022_/A VGND VGND VPWR VPWR _18022_/X sky130_fd_sc_hd__buf_2
X_12446_ _12446_/A VGND VGND VPWR VPWR _25447_/D sky130_fd_sc_hd__inv_2
X_15234_ _15204_/B _15233_/X VGND VGND VPWR VPWR _15234_/X sky130_fd_sc_hd__or2_4
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12377_ _12413_/A _12377_/B _12377_/C VGND VGND VPWR VPWR _25464_/D sky130_fd_sc_hd__and3_4
X_15165_ _15165_/A _15163_/X _15164_/X VGND VGND VPWR VPWR _25039_/D sky130_fd_sc_hd__and3_4
XFILLER_176_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16676__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14116_ _14086_/A _14092_/X _14095_/A _14093_/Y VGND VGND VPWR VPWR _14116_/X sky130_fd_sc_hd__o22a_4
X_15096_ _25000_/Q VGND VGND VPWR VPWR _15333_/A sky130_fd_sc_hd__inv_2
X_19973_ _19973_/A VGND VGND VPWR VPWR _21944_/B sky130_fd_sc_hd__inv_2
XANTENNA__22749__B1 _24835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18924_ _23917_/Q VGND VGND VPWR VPWR _18924_/Y sky130_fd_sc_hd__inv_2
X_14047_ _14044_/X VGND VGND VPWR VPWR _14073_/A sky130_fd_sc_hd__inv_2
XANTENNA__14540__A HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16428__B1 _16062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18855_ _16505_/Y _24138_/Q _16505_/Y _24138_/Q VGND VGND VPWR VPWR _18855_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16979__A1 _24745_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18947__A _18947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17806_ _17790_/A _17796_/X _17806_/C VGND VGND VPWR VPWR _24281_/D sky130_fd_sc_hd__and3_4
XFILLER_227_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18786_ _18786_/A _18815_/B VGND VGND VPWR VPWR _18786_/X sky130_fd_sc_hd__or2_4
X_15998_ _15998_/A VGND VGND VPWR VPWR _15998_/X sky130_fd_sc_hd__buf_2
XANTENNA__22469__A _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24246__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21373__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17737_ _17736_/X VGND VGND VPWR VPWR _17737_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19917__B2 _19900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14949_ _15204_/A _24427_/Q _15204_/A _24427_/Q VGND VGND VPWR VPWR _14949_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_20_0_HCLK_A clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12995__A _13028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16467__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17668_ _17574_/D _17668_/B VGND VGND VPWR VPWR _17669_/B sky130_fd_sc_hd__or2_4
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19407_ _23747_/Q VGND VGND VPWR VPWR _19407_/Y sky130_fd_sc_hd__inv_2
X_16619_ _24515_/Q VGND VGND VPWR VPWR _16619_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25134__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17599_ _17516_/A _17598_/Y VGND VGND VPWR VPWR _17599_/X sky130_fd_sc_hd__or2_4
XANTENNA__25197__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_195_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19338_ _23771_/Q VGND VGND VPWR VPWR _19338_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_245_0_HCLK clkbuf_7_122_0_HCLK/X VGND VGND VPWR VPWR _25015_/CLK sky130_fd_sc_hd__clkbuf_1
X_19269_ _19268_/Y _19266_/X _16885_/X _19266_/X VGND VGND VPWR VPWR _19269_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23229__B2 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21300_ _21300_/A VGND VGND VPWR VPWR _21306_/C sky130_fd_sc_hd__buf_2
X_22280_ _22130_/B VGND VGND VPWR VPWR _22280_/X sky130_fd_sc_hd__buf_2
XFILLER_148_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25034__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21231_ _15661_/A _21230_/X _13658_/Y _15661_/A VGND VGND VPWR VPWR _21231_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22651__B _22654_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21162_ _21155_/X _21157_/X _21162_/C _21161_/X VGND VGND VPWR VPWR _21162_/X sky130_fd_sc_hd__and4_4
XFILLER_132_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21660__B1 _17725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20113_ _23498_/Q VGND VGND VPWR VPWR _20113_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18408__A1 _22927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21093_ _21583_/A VGND VGND VPWR VPWR _21864_/C sky130_fd_sc_hd__buf_2
XFILLER_120_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16419__B1 _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20044_ _20043_/Y _20039_/X _19820_/X _20039_/X VGND VGND VPWR VPWR _20044_/X sky130_fd_sc_hd__a2bb2o_4
X_24921_ _24032_/CLK _15562_/X HRESETn VGND VGND VPWR VPWR _15559_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_219_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25413__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24852_ _24907_/CLK _24852_/D HRESETn VGND VGND VPWR VPWR _13129_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22379__A _22379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24336__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23803_ _23806_/CLK _23803_/D VGND VGND VPWR VPWR _19249_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_85_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21283__A _21283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _21994_/X VGND VGND VPWR VPWR _21995_/Y sky130_fd_sc_hd__inv_2
X_24783_ _24889_/CLK _24783_/D HRESETn VGND VGND VPWR VPWR _13527_/B sky130_fd_sc_hd__dfrtp_4
XPHY_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _16650_/Y _20846_/A _20919_/A _20945_/Y VGND VGND VPWR VPWR _20947_/A sky130_fd_sc_hd__o22a_4
X_23734_ _25073_/CLK _23734_/D VGND VGND VPWR VPWR _19444_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14609__B _15694_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23969__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _24046_/Q VGND VGND VPWR VPWR _20877_/Y sky130_fd_sc_hd__inv_2
X_23665_ _23665_/CLK _19655_/X VGND VGND VPWR VPWR _13221_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_55_0_HCLK clkbuf_6_54_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_55_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25404_ _24032_/CLK _12720_/X HRESETn VGND VGND VPWR VPWR _12578_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22616_ _16763_/A _22534_/X _22535_/X VGND VGND VPWR VPWR _22616_/X sky130_fd_sc_hd__o21a_4
XFILLER_186_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23596_ _23525_/CLK _23596_/D VGND VGND VPWR VPWR _23596_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22547_ _22546_/X VGND VGND VPWR VPWR _22577_/B sky130_fd_sc_hd__inv_2
X_25335_ _25346_/CLK _13105_/Y HRESETn VGND VGND VPWR VPWR _12299_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12300_ _12983_/D _24820_/Q _12983_/D _24820_/Q VGND VGND VPWR VPWR _12301_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_6_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13280_ _13150_/X _13276_/X _13280_/C VGND VGND VPWR VPWR _13280_/X sky130_fd_sc_hd__or3_4
XFILLER_154_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22478_ _21080_/X VGND VGND VPWR VPWR _22478_/X sky130_fd_sc_hd__buf_2
X_25266_ _24172_/CLK _13816_/X HRESETn VGND VGND VPWR VPWR _25266_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_212_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11719__B1 _11718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12231_ _12418_/A _24761_/Q _12418_/A _24761_/Q VGND VGND VPWR VPWR _12239_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21429_ _21424_/X _21425_/X _21427_/X _12550_/A _21428_/X VGND VGND VPWR VPWR _21430_/B
+ sky130_fd_sc_hd__a32o_4
X_24217_ _25285_/CLK _24217_/D HRESETn VGND VGND VPWR VPWR _24217_/Q sky130_fd_sc_hd__dfrtp_4
X_25197_ _25043_/CLK _14223_/X HRESETn VGND VGND VPWR VPWR _25197_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_135_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22561__B _21337_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16658__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12162_ SSn_S3 _12161_/Y _12076_/X _12161_/Y VGND VGND VPWR VPWR _25466_/D sky130_fd_sc_hd__a2bb2o_4
X_24148_ _24148_/CLK _24148_/D HRESETn VGND VGND VPWR VPWR _24148_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21458__A _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16992__A1_N _24717_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24757__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12093_ _12092_/Y _12090_/X _11757_/X _12090_/X VGND VGND VPWR VPWR _25477_/D sky130_fd_sc_hd__a2bb2o_4
X_16970_ _24735_/Q _24392_/Q _16024_/Y _16969_/Y VGND VGND VPWR VPWR _16977_/A sky130_fd_sc_hd__o22a_4
X_24079_ _24073_/CLK _24079_/D HRESETn VGND VGND VPWR VPWR _20479_/B sky130_fd_sc_hd__dfrtp_4
X_15921_ _15670_/X _15918_/B VGND VGND VPWR VPWR _15921_/X sky130_fd_sc_hd__or2_4
XANTENNA__22746__A3 _22296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18640_ _16576_/A _18755_/B _16608_/Y _24131_/Q VGND VGND VPWR VPWR _18647_/A sky130_fd_sc_hd__a2bb2o_4
X_15852_ _15851_/X VGND VGND VPWR VPWR _22638_/B sky130_fd_sc_hd__buf_2
XFILLER_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14803_ _14803_/A VGND VGND VPWR VPWR _14830_/A sky130_fd_sc_hd__buf_2
XANTENNA__16830__B1 _15743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18571_ _18400_/Y _18567_/X VGND VGND VPWR VPWR _18571_/Y sky130_fd_sc_hd__nand2_4
XFILLER_92_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15783_ _15813_/A VGND VGND VPWR VPWR _15783_/X sky130_fd_sc_hd__buf_2
X_12995_ _13028_/A VGND VGND VPWR VPWR _12998_/A sky130_fd_sc_hd__buf_2
XFILLER_205_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17522_ _25522_/Q _17521_/A _11783_/Y _17521_/Y VGND VGND VPWR VPWR _17525_/C sky130_fd_sc_hd__o22a_4
XFILLER_45_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14734_ _14726_/X _14733_/Y _14720_/A _14718_/Y VGND VGND VPWR VPWR _25067_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16930__A1_N _16131_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11946_ _11929_/A VGND VGND VPWR VPWR _11947_/A sky130_fd_sc_hd__inv_2
XFILLER_55_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17453_ _17452_/A _13284_/A _20387_/A _13385_/A VGND VGND VPWR VPWR _17453_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14665_ _14705_/A VGND VGND VPWR VPWR _14672_/A sky130_fd_sc_hd__buf_2
XANTENNA__20390__B1 _18250_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11877_ _11869_/A _11896_/B _11876_/Y VGND VGND VPWR VPWR _11877_/X sky130_fd_sc_hd__o21a_4
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25545__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16404_ _16404_/A VGND VGND VPWR VPWR _16404_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13616_ _25078_/Q VGND VGND VPWR VPWR _18082_/A sky130_fd_sc_hd__inv_2
X_17384_ _17384_/A VGND VGND VPWR VPWR _17384_/X sky130_fd_sc_hd__buf_2
X_14596_ _14551_/X _14595_/Y _14588_/X _14591_/X _13560_/A VGND VGND VPWR VPWR _25086_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__22131__A1 _22129_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22131__B2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19123_ _19121_/Y _19119_/X _19122_/X _19119_/X VGND VGND VPWR VPWR _19123_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16335_ _16334_/Y _16332_/X _15965_/X _16332_/X VGND VGND VPWR VPWR _16335_/X sky130_fd_sc_hd__a2bb2o_4
X_13547_ _25094_/Q VGND VGND VPWR VPWR _14561_/A sky130_fd_sc_hd__inv_2
XFILLER_71_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19054_ _19054_/A VGND VGND VPWR VPWR _19054_/X sky130_fd_sc_hd__buf_2
X_16266_ _16265_/Y _16184_/X _15475_/X _16184_/X VGND VGND VPWR VPWR _16266_/X sky130_fd_sc_hd__a2bb2o_4
X_13478_ _25318_/Q VGND VGND VPWR VPWR _13478_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_12_0_HCLK clkbuf_7_6_0_HCLK/X VGND VGND VPWR VPWR _23526_/CLK sky130_fd_sc_hd__clkbuf_1
X_18005_ _18004_/X _23777_/Q VGND VGND VPWR VPWR _18008_/B sky130_fd_sc_hd__or2_4
X_15217_ _15214_/C _15214_/D VGND VGND VPWR VPWR _15221_/A sky130_fd_sc_hd__or2_4
XFILLER_161_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12429_ _12201_/Y _12428_/X _12382_/X VGND VGND VPWR VPWR _12429_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__23092__C1 _23091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_75_0_HCLK clkbuf_8_74_0_HCLK/A VGND VGND VPWR VPWR _24639_/CLK sky130_fd_sc_hd__clkbuf_1
X_16197_ _23170_/A VGND VGND VPWR VPWR _16197_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16649__B1 _16464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15148_ _24979_/Q VGND VGND VPWR VPWR _15148_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21368__A _21368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24498__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15079_ _15078_/Y VGND VGND VPWR VPWR _15366_/A sky130_fd_sc_hd__buf_2
X_19956_ _19955_/Y _19953_/X _19620_/X _19953_/X VGND VGND VPWR VPWR _23556_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21518__D _21518_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24427__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18907_ _17541_/Y _11794_/X HWDATA[28] _11794_/X VGND VGND VPWR VPWR _18907_/X sky130_fd_sc_hd__a2bb2o_4
X_19887_ _19886_/Y _19884_/X _19610_/X _19884_/X VGND VGND VPWR VPWR _23583_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18838_ _24555_/Q _24134_/Q _16515_/Y _18797_/A VGND VGND VPWR VPWR _18838_/X sky130_fd_sc_hd__o22a_4
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22199__A _22199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24080__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18769_ _18769_/A _18768_/Y VGND VGND VPWR VPWR _18769_/X sky130_fd_sc_hd__or2_4
XFILLER_64_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20800_ _13106_/B VGND VGND VPWR VPWR _20800_/Y sky130_fd_sc_hd__inv_2
X_21780_ _21769_/A _21778_/X _21779_/X VGND VGND VPWR VPWR _21780_/X sky130_fd_sc_hd__and3_4
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22927__A _22927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20731_ _20780_/A VGND VGND VPWR VPWR _20731_/X sky130_fd_sc_hd__buf_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15927__A2 _15887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23450_ _24413_/CLK _23450_/D VGND VGND VPWR VPWR _23450_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19301__A _19006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20662_ _14220_/Y _20615_/A _20629_/A _20661_/X VGND VGND VPWR VPWR _20663_/A sky130_fd_sc_hd__a211o_4
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22401_ _23401_/Q _22397_/B VGND VGND VPWR VPWR _22401_/X sky130_fd_sc_hd__or2_4
X_23381_ _23808_/CLK _23381_/D VGND VGND VPWR VPWR _23381_/Q sky130_fd_sc_hd__dfxtp_4
X_20593_ _20593_/A VGND VGND VPWR VPWR _20593_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22332_ _22331_/Y _21349_/A _14207_/Y _14209_/X VGND VGND VPWR VPWR _22333_/A sky130_fd_sc_hd__o22a_4
X_25120_ _25109_/CLK _25120_/D HRESETn VGND VGND VPWR VPWR _25120_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25051_ _25052_/CLK _14839_/X HRESETn VGND VGND VPWR VPWR _25051_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22263_ _21462_/A _22263_/B _22263_/C VGND VGND VPWR VPWR _22263_/X sky130_fd_sc_hd__and3_4
XFILLER_247_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18629__B2 _18693_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16660__A _16660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24002_ _25226_/CLK _24002_/D HRESETn VGND VGND VPWR VPWR _24002_/Q sky130_fd_sc_hd__dfrtp_4
X_21214_ _21214_/A _19570_/X VGND VGND VPWR VPWR _21214_/X sky130_fd_sc_hd__or2_4
XFILLER_151_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22194_ _22194_/A _22190_/X _22193_/X VGND VGND VPWR VPWR _22194_/X sky130_fd_sc_hd__and3_4
XANTENNA__24850__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21145_ _13523_/A _12082_/A _13452_/Y _12082_/A VGND VGND VPWR VPWR _21145_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19971__A _19962_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24168__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21076_ _21075_/Y VGND VGND VPWR VPWR _21077_/A sky130_fd_sc_hd__buf_2
XFILLER_101_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20027_ _23532_/Q VGND VGND VPWR VPWR _21467_/B sky130_fd_sc_hd__inv_2
X_24904_ _24903_/CLK _15606_/X HRESETn VGND VGND VPWR VPWR _24904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16812__B1 HWDATA[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18404__A1_N _22996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24835_ _24855_/CLK _15814_/X HRESETn VGND VGND VPWR VPWR _24835_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13626__B1 _14610_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11797_/Y _11799_/X VGND VGND VPWR VPWR _11802_/A sky130_fd_sc_hd__or2_4
XPHY_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _24802_/Q VGND VGND VPWR VPWR _12780_/Y sky130_fd_sc_hd__inv_2
X_24766_ _24766_/CLK _15952_/X HRESETn VGND VGND VPWR VPWR _22857_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _18354_/A _20324_/Y _21979_/A _20322_/Y VGND VGND VPWR VPWR _21978_/X sky130_fd_sc_hd__o22a_4
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22361__A1 _17709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21741__A _16530_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11728_/Y _11723_/X _11730_/X _11723_/X VGND VGND VPWR VPWR _11731_/X sky130_fd_sc_hd__a2bb2o_4
X_23717_ _23427_/CLK _19495_/X VGND VGND VPWR VPWR _23717_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _20928_/Y _20925_/Y _20932_/B VGND VGND VPWR VPWR _20929_/X sky130_fd_sc_hd__o21a_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24697_ _24696_/CLK _24697_/D HRESETn VGND VGND VPWR VPWR _22778_/A sky130_fd_sc_hd__dfrtp_4
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _25126_/Q VGND VGND VPWR VPWR _14450_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _15541_/A _12038_/B VGND VGND VPWR VPWR _15984_/D sky130_fd_sc_hd__or2_4
X_23648_ _23644_/CLK _23648_/D VGND VGND VPWR VPWR _13273_/B sky130_fd_sc_hd__dfxtp_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13433_/A _13397_/X _13401_/C VGND VGND VPWR VPWR _13402_/C sky130_fd_sc_hd__or3_4
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14381_ _20506_/D _14371_/X _14380_/X _14373_/X VGND VGND VPWR VPWR _14381_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23579_ _23555_/CLK _23579_/D VGND VGND VPWR VPWR _19895_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16120_ _24698_/Q VGND VGND VPWR VPWR _16120_/Y sky130_fd_sc_hd__inv_2
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ _13396_/A _18944_/A VGND VGND VPWR VPWR _13333_/C sky130_fd_sc_hd__or2_4
X_25318_ _25479_/CLK _13479_/X HRESETn VGND VGND VPWR VPWR _25318_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21872__B1 _24859_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22572__A _21019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24938__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16051_ _16049_/Y _16045_/X _15752_/X _16050_/X VGND VGND VPWR VPWR _24725_/D sky130_fd_sc_hd__a2bb2o_4
X_13263_ _13263_/A _13263_/B _13262_/X VGND VGND VPWR VPWR _13263_/X sky130_fd_sc_hd__and3_4
X_25249_ _25249_/CLK _13862_/X HRESETn VGND VGND VPWR VPWR _25249_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22291__B _22417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15002_ _15002_/A VGND VGND VPWR VPWR _15254_/A sky130_fd_sc_hd__buf_2
X_12214_ _12203_/X _12214_/B _12214_/C _12213_/X VGND VGND VPWR VPWR _12215_/D sky130_fd_sc_hd__or4_4
XANTENNA__20427__B2 _20409_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13194_ _13288_/A VGND VGND VPWR VPWR _13254_/A sky130_fd_sc_hd__buf_2
XFILLER_123_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24591__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12145_ _12145_/A _12145_/B _12145_/C _12144_/X VGND VGND VPWR VPWR _18372_/D sky130_fd_sc_hd__or4_4
X_19810_ _16858_/X VGND VGND VPWR VPWR _19810_/X sky130_fd_sc_hd__buf_2
XFILLER_123_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24520__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12076_ _14262_/A VGND VGND VPWR VPWR _12076_/X sky130_fd_sc_hd__buf_2
X_16953_ _24713_/Q VGND VGND VPWR VPWR _16953_/Y sky130_fd_sc_hd__inv_2
X_19741_ _19737_/Y _19740_/X _19652_/X _19740_/X VGND VGND VPWR VPWR _19741_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21916__A _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15904_ _24784_/Q _15904_/B VGND VGND VPWR VPWR _15904_/Y sky130_fd_sc_hd__nor2_4
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19672_ _19672_/A VGND VGND VPWR VPWR _19672_/Y sky130_fd_sc_hd__inv_2
X_16884_ _19852_/A VGND VGND VPWR VPWR _16884_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18623_ _24150_/Q VGND VGND VPWR VPWR _18677_/A sky130_fd_sc_hd__inv_2
XFILLER_77_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15835_ _15818_/X _15829_/X _15770_/X _24820_/Q _15786_/X VGND VGND VPWR VPWR _15835_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_65_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18554_ _18556_/B VGND VGND VPWR VPWR _18555_/B sky130_fd_sc_hd__inv_2
X_15766_ _12540_/Y _15759_/X _15472_/X _15759_/X VGND VGND VPWR VPWR _15766_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12978_ _12975_/Y _12357_/Y _12977_/X VGND VGND VPWR VPWR _12978_/X sky130_fd_sc_hd__or3_4
XFILLER_206_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17505_ _11790_/Y _24291_/Q _11790_/Y _24291_/Q VGND VGND VPWR VPWR _17505_/X sky130_fd_sc_hd__a2bb2o_4
X_14717_ _14702_/X _14716_/X VGND VGND VPWR VPWR _14718_/A sky130_fd_sc_hd__or2_4
X_11929_ _11929_/A VGND VGND VPWR VPWR _11929_/X sky130_fd_sc_hd__buf_2
X_18485_ _24189_/Q _18484_/Y VGND VGND VPWR VPWR _18487_/B sky130_fd_sc_hd__or2_4
XANTENNA__20363__B1 _19617_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15697_ _14366_/A _15697_/B VGND VGND VPWR VPWR _15698_/A sky130_fd_sc_hd__or2_4
XANTENNA__15909__A2 _14764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17436_ _12084_/A _17436_/B _17436_/C VGND VGND VPWR VPWR _17436_/X sky130_fd_sc_hd__or3_4
X_14648_ _14648_/A _14784_/A VGND VGND VPWR VPWR _14648_/X sky130_fd_sc_hd__or2_4
XFILLER_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17367_ _17351_/A _17367_/B _17366_/Y VGND VGND VPWR VPWR _24347_/D sky130_fd_sc_hd__and3_4
X_14579_ _13757_/Y VGND VGND VPWR VPWR _14579_/X sky130_fd_sc_hd__buf_2
XANTENNA__18859__B2 _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19106_ _18965_/A VGND VGND VPWR VPWR _19106_/X sky130_fd_sc_hd__buf_2
X_16318_ _16318_/A VGND VGND VPWR VPWR _16344_/A sky130_fd_sc_hd__buf_2
X_17298_ _17298_/A _17301_/B VGND VGND VPWR VPWR _17299_/C sky130_fd_sc_hd__or2_4
XFILLER_158_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19037_ _19037_/A VGND VGND VPWR VPWR _19037_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24679__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16249_ _24654_/Q VGND VGND VPWR VPWR _16249_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22407__A2 _22282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24608__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22812__C1 _22811_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22958__A3 _22719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17295__B1 _17276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12108__B1 _11786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24261__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21826__A _13772_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19939_ _19939_/A _19939_/B _19479_/X VGND VGND VPWR VPWR _19939_/X sky130_fd_sc_hd__or3_4
XFILLER_228_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22950_ _16667_/Y _22794_/A _15583_/Y _22832_/X VGND VGND VPWR VPWR _22950_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21901_ _21901_/A _21891_/X _21900_/X VGND VGND VPWR VPWR _21901_/X sky130_fd_sc_hd__or3_4
XFILLER_233_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15543__B _21290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22881_ _20767_/Y _21122_/X _20906_/Y _21227_/X VGND VGND VPWR VPWR _22882_/B sky130_fd_sc_hd__o22a_4
XANTENNA__11882__A2 _11934_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24620_ _24346_/CLK _24620_/D HRESETn VGND VGND VPWR VPWR _24620_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_7_120_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_241_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21832_ _21832_/A VGND VGND VPWR VPWR _21832_/X sky130_fd_sc_hd__buf_2
XANTENNA__18848__A2_N _24143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22657__A _21087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21763_ _14753_/X _20101_/Y VGND VGND VPWR VPWR _21763_/X sky130_fd_sc_hd__or2_4
X_24551_ _24551_/CLK _16529_/X HRESETn VGND VGND VPWR VPWR _16527_/A sky130_fd_sc_hd__dfrtp_4
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16655__A _16655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20714_ _22291_/A _20708_/X _20696_/X _20713_/Y VGND VGND VPWR VPWR _20715_/A sky130_fd_sc_hd__o22a_4
X_23502_ _23494_/CLK _23502_/D VGND VGND VPWR VPWR _23502_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21694_ _18274_/A _21692_/X _21510_/X _21693_/Y VGND VGND VPWR VPWR _21695_/A sky130_fd_sc_hd__a211o_4
X_24482_ _24486_/CLK _16710_/X HRESETn VGND VGND VPWR VPWR _16708_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_178_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20645_ _20645_/A _20643_/Y _20661_/C VGND VGND VPWR VPWR _20645_/X sky130_fd_sc_hd__and3_4
X_23433_ _23441_/CLK _23433_/D VGND VGND VPWR VPWR _23433_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23364_ _23364_/A VGND VGND VPWR VPWR IRQ[20] sky130_fd_sc_hd__buf_2
X_20576_ _23944_/Q _18877_/X VGND VGND VPWR VPWR _20576_/Y sky130_fd_sc_hd__nand2_4
XFILLER_165_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17522__A1 _25522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25103_ _25146_/CLK _14520_/X HRESETn VGND VGND VPWR VPWR _21347_/A sky130_fd_sc_hd__dfrtp_4
X_22315_ _22314_/X VGND VGND VPWR VPWR _22315_/Y sky130_fd_sc_hd__inv_2
X_23295_ _20817_/Y _22290_/X _20956_/Y _22794_/X VGND VGND VPWR VPWR _23296_/B sky130_fd_sc_hd__o22a_4
XFILLER_106_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24349__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22246_ _22251_/A _22246_/B VGND VGND VPWR VPWR _22248_/B sky130_fd_sc_hd__or2_4
X_25034_ _25035_/CLK _25034_/D HRESETn VGND VGND VPWR VPWR _25034_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12898__A1 _12813_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22177_ _13490_/Y _12086_/A _12017_/Y _12057_/A VGND VGND VPWR VPWR _22177_/X sky130_fd_sc_hd__o22a_4
XFILLER_239_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21128_ _25334_/Q _21128_/B VGND VGND VPWR VPWR _21128_/Y sky130_fd_sc_hd__nor2_4
XFILLER_120_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21736__A _21736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13950_ _13949_/A _13948_/Y _13949_/Y _13947_/X VGND VGND VPWR VPWR _13950_/X sky130_fd_sc_hd__o22a_4
X_21059_ _21059_/A _21058_/X VGND VGND VPWR VPWR _21059_/X sky130_fd_sc_hd__or2_4
XFILLER_87_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21231__A1_N _15661_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12901_ _12766_/Y _12906_/B _12854_/X VGND VGND VPWR VPWR _12901_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_207_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23984__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13881_ _13880_/X VGND VGND VPWR VPWR _15421_/B sky130_fd_sc_hd__buf_2
X_15620_ _22291_/A _15613_/X _15619_/X _15613_/X VGND VGND VPWR VPWR _24899_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13254__A _13254_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12832_ _25369_/Q VGND VGND VPWR VPWR _12833_/C sky130_fd_sc_hd__inv_2
X_24818_ _24855_/CLK _15840_/X HRESETn VGND VGND VPWR VPWR _12592_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22567__A _16691_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15551_ _15550_/Y VGND VGND VPWR VPWR _15608_/A sky130_fd_sc_hd__buf_2
XFILLER_61_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12763_ _22420_/A VGND VGND VPWR VPWR _12763_/Y sky130_fd_sc_hd__inv_2
X_24749_ _24696_/CLK _24749_/D HRESETn VGND VGND VPWR VPWR _21442_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14490_/C VGND VGND VPWR VPWR _14502_/X sky130_fd_sc_hd__buf_2
XFILLER_230_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11683_/X VGND VGND VPWR VPWR _11714_/X sky130_fd_sc_hd__buf_2
X_18270_ _13783_/D _18256_/X _11788_/X _21504_/A _18264_/X VGND VGND VPWR VPWR _24222_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_187_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _24069_/D _15482_/B VGND VGND VPWR VPWR _15483_/A sky130_fd_sc_hd__or2_4
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12706_/A _12693_/X VGND VGND VPWR VPWR _12707_/B sky130_fd_sc_hd__or2_4
XFILLER_230_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_25_0_HCLK clkbuf_5_25_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _17214_/X _17221_/B _17218_/X _17220_/X VGND VGND VPWR VPWR _17221_/X sky130_fd_sc_hd__or4_4
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14433_/A VGND VGND VPWR VPWR _14433_/Y sky130_fd_sc_hd__inv_2
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14085__A scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17152_ _16982_/Y _17151_/X VGND VGND VPWR VPWR _17153_/B sky130_fd_sc_hd__or2_4
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14364_ _14364_/A VGND VGND VPWR VPWR _14366_/A sky130_fd_sc_hd__buf_2
XFILLER_155_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16103_ _24705_/Q VGND VGND VPWR VPWR _16103_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24772__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13315_ _13225_/A VGND VGND VPWR VPWR _13445_/A sky130_fd_sc_hd__buf_2
XANTENNA__22733__C _22732_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17083_ _17070_/A _17075_/X _17083_/C VGND VGND VPWR VPWR _24396_/D sky130_fd_sc_hd__and3_4
XFILLER_128_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14295_ _14295_/A VGND VGND VPWR VPWR _14295_/X sky130_fd_sc_hd__buf_2
XFILLER_155_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24701__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16034_ _16031_/Y _16033_/X _11726_/X _16033_/X VGND VGND VPWR VPWR _24732_/D sky130_fd_sc_hd__a2bb2o_4
X_13246_ _13186_/X _13244_/X _25332_/Q _13245_/X VGND VGND VPWR VPWR _25332_/D sky130_fd_sc_hd__o22a_4
XFILLER_171_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24019__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17277__B1 _17276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13429__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13177_ _13157_/X _18909_/A VGND VGND VPWR VPWR _13179_/B sky130_fd_sc_hd__or2_4
XFILLER_184_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12333__A _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_149_0_HCLK clkbuf_7_74_0_HCLK/X VGND VGND VPWR VPWR _24188_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12128_ _25474_/Q _12127_/Y _25474_/Q _12127_/Y VGND VGND VPWR VPWR _12128_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17985_ _17999_/A VGND VGND VPWR VPWR _17985_/X sky130_fd_sc_hd__buf_2
XANTENNA__13838__B1 _13798_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12059_ _12058_/X VGND VGND VPWR VPWR _12060_/A sky130_fd_sc_hd__inv_2
X_16936_ _24286_/Q VGND VGND VPWR VPWR _16945_/A sky130_fd_sc_hd__inv_2
X_19724_ _19722_/Y _19718_/X _19633_/X _19723_/X VGND VGND VPWR VPWR _23640_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15644__A _15644_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18020__A _18020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22573__A1 _16895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16867_ _20099_/A VGND VGND VPWR VPWR _16867_/X sky130_fd_sc_hd__buf_2
X_19655_ _19654_/Y _19651_/X _19630_/X _19651_/X VGND VGND VPWR VPWR _19655_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15818_ _11706_/X VGND VGND VPWR VPWR _15818_/X sky130_fd_sc_hd__buf_2
X_18606_ _16557_/Y _18732_/A _16557_/Y _18732_/A VGND VGND VPWR VPWR _18607_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19586_ _19585_/X VGND VGND VPWR VPWR _19586_/Y sky130_fd_sc_hd__inv_2
X_16798_ _16793_/A VGND VGND VPWR VPWR _16799_/A sky130_fd_sc_hd__buf_2
XFILLER_80_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14263__B1 _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22477__A _22146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18537_ _18407_/Y _18541_/B _18536_/Y VGND VGND VPWR VPWR _24177_/D sky130_fd_sc_hd__o21a_4
X_15749_ _15745_/X _15738_/X _15748_/X _24866_/Q _15706_/X VGND VGND VPWR VPWR _15749_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_179_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18468_ _18468_/A _18442_/Y _18468_/C VGND VGND VPWR VPWR _18510_/D sky130_fd_sc_hd__or3_4
XFILLER_178_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17419_ _17417_/Y _17414_/X _17418_/X _17414_/X VGND VGND VPWR VPWR _24332_/D sky130_fd_sc_hd__a2bb2o_4
X_18399_ _16221_/Y _24174_/Q _16221_/Y _24174_/Q VGND VGND VPWR VPWR _18399_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22628__A2 _21098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15763__B1 _24859_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18690__A _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20430_ _20430_/A _20467_/C VGND VGND VPWR VPWR _20430_/X sky130_fd_sc_hd__or2_4
XFILLER_146_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20361_ _20361_/A VGND VGND VPWR VPWR _21671_/B sky130_fd_sc_hd__inv_2
XANTENNA__15515__B1 HADDR[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22100_ _24520_/Q _21863_/X _22098_/X _22099_/X VGND VGND VPWR VPWR _22101_/C sky130_fd_sc_hd__a211o_4
XANTENNA__24442__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23080_ _24740_/Q _21061_/X _21062_/X _23079_/X VGND VGND VPWR VPWR _23080_/X sky130_fd_sc_hd__a211o_4
X_20292_ _23431_/Q VGND VGND VPWR VPWR _22034_/B sky130_fd_sc_hd__inv_2
XFILLER_115_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22940__A _16485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_45_0_HCLK clkbuf_7_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22031_ _22024_/A _22029_/X _22030_/X VGND VGND VPWR VPWR _22031_/X sky130_fd_sc_hd__and3_4
XFILLER_114_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21556__A _21556_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16146__A1_N _16144_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15554__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23982_ _23986_/CLK _20651_/Y HRESETn VGND VGND VPWR VPWR _23982_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22933_ _15091_/A _23177_/B VGND VGND VPWR VPWR _22933_/X sky130_fd_sc_hd__or2_4
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22864_ _24630_/Q _22487_/X VGND VGND VPWR VPWR _22864_/X sky130_fd_sc_hd__or2_4
XFILLER_37_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25230__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22316__B2 _22181_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24603_ _25005_/CLK _16390_/X HRESETn VGND VGND VPWR VPWR _24603_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21815_ _21484_/X _21813_/X _21814_/X VGND VGND VPWR VPWR _21815_/X sky130_fd_sc_hd__and3_4
X_22795_ _20759_/Y _22290_/X _20898_/Y _22794_/X VGND VGND VPWR VPWR _22796_/B sky130_fd_sc_hd__o22a_4
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24534_ _24573_/CLK _16573_/X HRESETn VGND VGND VPWR VPWR _16571_/A sky130_fd_sc_hd__dfrtp_4
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21746_ _21746_/A _21745_/B VGND VGND VPWR VPWR _21746_/X sky130_fd_sc_hd__and2_4
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18940__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24465_ _24443_/CLK _16750_/X HRESETn VGND VGND VPWR VPWR _24465_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21677_ _21677_/A _21677_/B VGND VGND VPWR VPWR _21678_/C sky130_fd_sc_hd__or2_4
XANTENNA__12418__A _12418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12568__B1 _25411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23416_ _23575_/CLK _23416_/D VGND VGND VPWR VPWR _20331_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20628_ _20628_/A VGND VGND VPWR VPWR _20629_/A sky130_fd_sc_hd__buf_2
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24396_ _24377_/CLK _24396_/D HRESETn VGND VGND VPWR VPWR _17024_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20559_ _18874_/X _20559_/B _20553_/C VGND VGND VPWR VPWR _20559_/X sky130_fd_sc_hd__and3_4
X_23347_ _24224_/Q _21985_/X _23345_/X _23346_/Y VGND VGND VPWR VPWR _23347_/X sky130_fd_sc_hd__a211o_4
XFILLER_153_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13100_ _13097_/B _13100_/B _13091_/C VGND VGND VPWR VPWR _13100_/X sky130_fd_sc_hd__and3_4
XANTENNA__24183__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14080_ _14053_/A VGND VGND VPWR VPWR _20453_/C sky130_fd_sc_hd__buf_2
X_23278_ _24815_/Q _23278_/B VGND VGND VPWR VPWR _23278_/X sky130_fd_sc_hd__or2_4
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24112__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13031_ _12971_/Y _12985_/X VGND VGND VPWR VPWR _13032_/B sky130_fd_sc_hd__or2_4
X_25017_ _24967_/CLK _15258_/X HRESETn VGND VGND VPWR VPWR _25017_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22229_ _19578_/A _22229_/B VGND VGND VPWR VPWR _22229_/X sky130_fd_sc_hd__and2_4
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25389__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_2_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17770_ _23320_/A _17769_/Y VGND VGND VPWR VPWR _17772_/B sky130_fd_sc_hd__or2_4
X_14982_ _14982_/A VGND VGND VPWR VPWR _15185_/A sky130_fd_sc_hd__buf_2
XFILLER_66_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16721_ _16721_/A _16721_/B _22539_/A _21327_/B VGND VGND VPWR VPWR _16721_/X sky130_fd_sc_hd__and4_4
X_13933_ _13932_/X VGND VGND VPWR VPWR _13939_/B sky130_fd_sc_hd__inv_2
X_19440_ _19447_/A VGND VGND VPWR VPWR _19440_/X sky130_fd_sc_hd__buf_2
XFILLER_90_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16652_ _24505_/Q VGND VGND VPWR VPWR _16652_/Y sky130_fd_sc_hd__inv_2
X_13864_ _13860_/X _13863_/X _25189_/Q _13856_/X VGND VGND VPWR VPWR _13864_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22307__A1 _24522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15603_ _24905_/Q VGND VGND VPWR VPWR _15603_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12815_ _12805_/X _12815_/B _12811_/X _12814_/X VGND VGND VPWR VPWR _12815_/X sky130_fd_sc_hd__or4_4
X_19371_ _23760_/Q VGND VGND VPWR VPWR _19371_/Y sky130_fd_sc_hd__inv_2
X_16583_ _16582_/Y _16580_/X _16226_/X _16580_/X VGND VGND VPWR VPWR _24530_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13795_ _13794_/Y _13792_/X _13521_/X _13792_/X VGND VGND VPWR VPWR _13795_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16295__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18322_ _18322_/A VGND VGND VPWR VPWR _18322_/Y sky130_fd_sc_hd__inv_2
X_15534_ _17436_/B _15530_/X HADDR[2] _15533_/X VGND VGND VPWR VPWR _24927_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12746_ _22972_/A VGND VGND VPWR VPWR _12746_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18253_ _11808_/Y _18252_/X _17418_/X _18252_/X VGND VGND VPWR VPWR _18253_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15465_ _15465_/A VGND VGND VPWR VPWR _15465_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18850__A1_N _16492_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12677_ _12677_/A _12663_/X _12677_/C VGND VGND VPWR VPWR _25416_/D sky130_fd_sc_hd__and3_4
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _24346_/Q VGND VGND VPWR VPWR _17346_/C sky130_fd_sc_hd__inv_2
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ _14414_/Y _14415_/X _14384_/X _14415_/X VGND VGND VPWR VPWR _14416_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18184_ _17990_/X _18184_/B _18183_/X VGND VGND VPWR VPWR _18184_/X sky130_fd_sc_hd__and3_4
X_15396_ _15379_/A _15390_/B _15395_/Y VGND VGND VPWR VPWR _24985_/D sky130_fd_sc_hd__and3_4
XFILLER_129_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ _17038_/D _17131_/X VGND VGND VPWR VPWR _17136_/C sky130_fd_sc_hd__nand2_4
XFILLER_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14347_ _14344_/X _14346_/Y _12049_/A _14344_/X VGND VGND VPWR VPWR _14347_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22491__B1 _24725_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18015__A _18056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17066_ _17066_/A VGND VGND VPWR VPWR _24401_/D sky130_fd_sc_hd__inv_2
X_14278_ _14278_/A VGND VGND VPWR VPWR _14283_/A sky130_fd_sc_hd__inv_2
XFILLER_171_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16017_ _16016_/Y _16012_/X _15942_/X _16012_/X VGND VGND VPWR VPWR _24738_/D sky130_fd_sc_hd__a2bb2o_4
X_13229_ _13172_/A _13229_/B _13228_/X VGND VGND VPWR VPWR _13230_/C sky130_fd_sc_hd__and3_4
XFILLER_170_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12731__B1 _12830_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15374__A _15331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17968_ _18026_/A VGND VGND VPWR VPWR _17968_/X sky130_fd_sc_hd__buf_2
XANTENNA__25059__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19707_ _19694_/A VGND VGND VPWR VPWR _19707_/X sky130_fd_sc_hd__buf_2
X_16919_ _16919_/A _16919_/B _16919_/C _16918_/X VGND VGND VPWR VPWR _16920_/D sky130_fd_sc_hd__or4_4
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17899_ _17896_/Y _17906_/B _17898_/Y VGND VGND VPWR VPWR _17899_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_66_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19638_ _13343_/B VGND VGND VPWR VPWR _19638_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19569_ _14180_/A _12043_/Y _13765_/A _15657_/X VGND VGND VPWR VPWR _21159_/A sky130_fd_sc_hd__or4_4
XFILLER_179_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19175__B1 _19106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21600_ _21119_/X _21595_/Y _21596_/X _21599_/X VGND VGND VPWR VPWR _21600_/X sky130_fd_sc_hd__o22a_4
XFILLER_179_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22580_ _24425_/Q _21031_/X _22533_/X _22579_/X VGND VGND VPWR VPWR _22581_/C sky130_fd_sc_hd__a211o_4
XFILLER_61_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24694__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21531_ _15780_/B VGND VGND VPWR VPWR _21531_/X sky130_fd_sc_hd__buf_2
XANTENNA__12227__A2_N _24762_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22654__B _22654_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24623__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21462_ _21462_/A VGND VGND VPWR VPWR _21472_/A sky130_fd_sc_hd__buf_2
X_24250_ _23747_/CLK _24250_/D HRESETn VGND VGND VPWR VPWR _24250_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20413_ _22217_/B _20410_/X _16858_/X _20410_/X VGND VGND VPWR VPWR _20413_/X sky130_fd_sc_hd__a2bb2o_4
X_23201_ _15563_/Y _23292_/B VGND VGND VPWR VPWR _23201_/X sky130_fd_sc_hd__and2_4
XANTENNA__21285__A1 _21275_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21393_ _22197_/A _19268_/Y VGND VGND VPWR VPWR _21393_/X sky130_fd_sc_hd__or2_4
X_24181_ _24188_/CLK _24181_/D HRESETn VGND VGND VPWR VPWR _24181_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20344_ _20343_/Y _20341_/X _19620_/A _20341_/X VGND VGND VPWR VPWR _20344_/X sky130_fd_sc_hd__a2bb2o_4
X_23132_ _23132_/A _23063_/X VGND VGND VPWR VPWR _23132_/X sky130_fd_sc_hd__or2_4
XANTENNA__23026__A2 _23017_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23063_ _22530_/A VGND VGND VPWR VPWR _23063_/X sky130_fd_sc_hd__buf_2
X_20275_ _21921_/B _20272_/X _19974_/X _20272_/X VGND VGND VPWR VPWR _23438_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22014_ _22014_/A _19861_/Y VGND VGND VPWR VPWR _22017_/B sky130_fd_sc_hd__or2_4
XFILLER_161_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18989__B1 _18942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25482__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_132_0_HCLK clkbuf_7_66_0_HCLK/X VGND VGND VPWR VPWR _23391_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_124_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22537__A1 _15018_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_195_0_HCLK clkbuf_7_97_0_HCLK/X VGND VGND VPWR VPWR _24592_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_130_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23965_ _25249_/CLK _23965_/D HRESETn VGND VGND VPWR VPWR _23965_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23289__A1_N _17232_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22916_ _22429_/X VGND VGND VPWR VPWR _22916_/X sky130_fd_sc_hd__buf_2
XFILLER_44_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23896_ _23827_/CLK _23896_/D VGND VGND VPWR VPWR _18983_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_44_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22847_ _12216_/Y _21082_/X _16724_/A _12329_/Y _22846_/X VGND VGND VPWR VPWR _22848_/B
+ sky130_fd_sc_hd__o32a_4
XANTENNA__15975__B1 _24751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19166__B1 _19144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12600_ _12696_/A _12704_/A _12706_/A _12693_/A VGND VGND VPWR VPWR _12600_/X sky130_fd_sc_hd__or4_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _15636_/A _13453_/A _11659_/A _12039_/D VGND VGND VPWR VPWR _21283_/A sky130_fd_sc_hd__or4_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22778_ _22778_/A _22654_/B VGND VGND VPWR VPWR _22778_/X sky130_fd_sc_hd__or2_4
XFILLER_242_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13450__B2 _11950_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12531_ _25408_/Q _24862_/Q _12706_/A _12530_/Y VGND VGND VPWR VPWR _12532_/D sky130_fd_sc_hd__o22a_4
X_24517_ _24520_/CLK _16616_/X HRESETn VGND VGND VPWR VPWR _16615_/A sky130_fd_sc_hd__dfrtp_4
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21729_ _16259_/Y _16180_/A _16432_/A _16719_/A VGND VGND VPWR VPWR _21730_/B sky130_fd_sc_hd__a2bb2o_4
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15727__B1 _11695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25497_ _25499_/CLK _25497_/D HRESETn VGND VGND VPWR VPWR _11967_/A sky130_fd_sc_hd__dfrtp_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24364__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15250_ _15269_/A _15250_/B _15249_/X VGND VGND VPWR VPWR _15250_/X sky130_fd_sc_hd__and3_4
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12462_ _25444_/Q _12461_/Y VGND VGND VPWR VPWR _12464_/B sky130_fd_sc_hd__or2_4
X_24448_ _24477_/CLK _16785_/X HRESETn VGND VGND VPWR VPWR _24448_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15742__A3 _15741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14201_ _14201_/A VGND VGND VPWR VPWR _14201_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15181_ _14886_/A _15180_/Y VGND VGND VPWR VPWR _15181_/X sky130_fd_sc_hd__or2_4
XFILLER_153_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22473__B1 _22457_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12393_ _12279_/B _12494_/A VGND VGND VPWR VPWR _12396_/B sky130_fd_sc_hd__or2_4
X_24379_ _24725_/CLK _17145_/X HRESETn VGND VGND VPWR VPWR _16957_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14132_ _14099_/X _14131_/X _14414_/A _14125_/X VGND VGND VPWR VPWR _14132_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_153_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14063_ _20522_/A _14058_/X _14062_/X _14028_/B _14055_/X VGND VGND VPWR VPWR _14063_/X
+ sky130_fd_sc_hd__a32o_4
X_18940_ _18938_/Y _18934_/X _17421_/X _18939_/X VGND VGND VPWR VPWR _23912_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13014_ _13028_/A _13009_/Y _13013_/X VGND VGND VPWR VPWR _13015_/A sky130_fd_sc_hd__or3_4
XANTENNA__22776__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18871_ _18871_/A VGND VGND VPWR VPWR _18871_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_91_0_HCLK clkbuf_7_91_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17822_ _16911_/Y _17827_/B _16952_/X VGND VGND VPWR VPWR _17822_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_95_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14466__B1 _14403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14965_ _15066_/A _24440_/Q _25028_/Q _14964_/Y VGND VGND VPWR VPWR _14969_/C sky130_fd_sc_hd__a2bb2o_4
X_17753_ _16915_/Y _16904_/Y _16895_/A _17753_/D VGND VGND VPWR VPWR _17753_/X sky130_fd_sc_hd__or4_4
XFILLER_181_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13916_ _13902_/A _13876_/A _13916_/C _13903_/B VGND VGND VPWR VPWR _13942_/C sky130_fd_sc_hd__or4_4
X_16704_ _16692_/A VGND VGND VPWR VPWR _16704_/X sky130_fd_sc_hd__buf_2
XFILLER_47_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17684_ _17627_/A VGND VGND VPWR VPWR _17688_/C sky130_fd_sc_hd__buf_2
XFILLER_47_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14896_ _25034_/Q VGND VGND VPWR VPWR _15066_/A sky130_fd_sc_hd__inv_2
XFILLER_62_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16635_ _16170_/B _16621_/X VGND VGND VPWR VPWR _16635_/X sky130_fd_sc_hd__and2_4
X_19423_ _18111_/B VGND VGND VPWR VPWR _19423_/Y sky130_fd_sc_hd__inv_2
X_13847_ _13842_/B VGND VGND VPWR VPWR _13847_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15966__B1 _15965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19157__B1 _19063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16566_ _16566_/A VGND VGND VPWR VPWR _16566_/Y sky130_fd_sc_hd__inv_2
X_19354_ _19353_/Y _19348_/X _19221_/X _19348_/X VGND VGND VPWR VPWR _19354_/X sky130_fd_sc_hd__a2bb2o_4
X_13778_ _14395_/A _14462_/A VGND VGND VPWR VPWR _14243_/A sky130_fd_sc_hd__or2_4
XANTENNA__18904__B1 _24114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15517_ _15516_/Y _15512_/X HADDR[10] _15512_/X VGND VGND VPWR VPWR _15517_/X sky130_fd_sc_hd__a2bb2o_4
X_18305_ _21473_/A _18302_/Y VGND VGND VPWR VPWR _18305_/X sky130_fd_sc_hd__and2_4
X_12729_ _21015_/A _12382_/X _12728_/Y VGND VGND VPWR VPWR _25400_/D sky130_fd_sc_hd__o21a_4
X_19285_ _19285_/A VGND VGND VPWR VPWR _19285_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15718__B1 _15564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16497_ _16494_/Y _16496_/X _16320_/X _16496_/X VGND VGND VPWR VPWR _16497_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12058__A _16181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20711__B1 _20696_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18236_ _18236_/A VGND VGND VPWR VPWR _18236_/X sky130_fd_sc_hd__buf_2
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15448_ _13935_/A _15444_/X _15441_/X _13934_/C _15447_/X VGND VGND VPWR VPWR _24965_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24034__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18167_ _18103_/A _23764_/Q VGND VGND VPWR VPWR _18169_/B sky130_fd_sc_hd__or2_4
X_15379_ _15379_/A _15377_/X _15378_/X VGND VGND VPWR VPWR _24989_/D sky130_fd_sc_hd__and3_4
XFILLER_191_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17118_ _17120_/B VGND VGND VPWR VPWR _17118_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15800__A1_N _12309_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18098_ _18098_/A _18098_/B _18098_/C VGND VGND VPWR VPWR _18099_/C sky130_fd_sc_hd__and3_4
XANTENNA__16143__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22490__A _21127_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17049_ _17050_/A _17050_/B VGND VGND VPWR VPWR _17051_/B sky130_fd_sc_hd__or2_4
XFILLER_171_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20060_ _20053_/X _18328_/A _18257_/X _13335_/B _20055_/X VGND VGND VPWR VPWR _23518_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_205_0_HCLK clkbuf_8_205_0_HCLK/A VGND VGND VPWR VPWR _24558_/CLK sky130_fd_sc_hd__clkbuf_1
X_23750_ _23785_/CLK _23750_/D VGND VGND VPWR VPWR _18110_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_54_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20962_ _24242_/Q _14608_/Y _15907_/Y _24784_/Q _15681_/X VGND VGND VPWR VPWR _20962_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_242_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21742__A2 _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22701_ _22701_/A _22701_/B VGND VGND VPWR VPWR _22701_/X sky130_fd_sc_hd__or2_4
XFILLER_241_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24875__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ _23575_/CLK _23681_/D VGND VGND VPWR VPWR _23681_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15957__B1 _24764_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ _13650_/X VGND VGND VPWR VPWR _20921_/C sky130_fd_sc_hd__buf_2
XANTENNA__14448__A _14455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25420_ _25409_/CLK _12666_/X HRESETn VGND VGND VPWR VPWR _25420_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24804__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22632_ _22632_/A _22631_/X VGND VGND VPWR VPWR _22632_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12166__A2_N _22597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25351_ _25344_/CLK _13052_/X HRESETn VGND VGND VPWR VPWR _12290_/A sky130_fd_sc_hd__dfrtp_4
X_22563_ _21077_/A _22560_/X _21114_/X _22562_/X VGND VGND VPWR VPWR _22563_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__20702__B1 _20696_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24302_ _24302_/CLK _24302_/D HRESETn VGND VGND VPWR VPWR _24302_/Q sky130_fd_sc_hd__dfrtp_4
X_21514_ _21513_/X VGND VGND VPWR VPWR _21514_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25282_ _24227_/CLK _25282_/D HRESETn VGND VGND VPWR VPWR _11829_/A sky130_fd_sc_hd__dfrtp_4
X_22494_ _22494_/A _22654_/B VGND VGND VPWR VPWR _22494_/X sky130_fd_sc_hd__or2_4
XANTENNA__20185__A _20180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23199__C _22140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24233_ _24233_/CLK _18251_/X HRESETn VGND VGND VPWR VPWR _24233_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22455__B1 _16600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21445_ _21034_/X VGND VGND VPWR VPWR _21445_/X sky130_fd_sc_hd__buf_2
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14183__A _14182_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21376_ _19592_/A _21959_/B _19542_/Y _21959_/B VGND VGND VPWR VPWR _21376_/X sky130_fd_sc_hd__a2bb2o_4
X_24164_ _24654_/CLK _18581_/X HRESETn VGND VGND VPWR VPWR _18395_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16134__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20327_ _19939_/A _19939_/B _19455_/X VGND VGND VPWR VPWR _20328_/A sky130_fd_sc_hd__or3_4
X_23115_ _23160_/A _23103_/X _23115_/C _23115_/D VGND VGND VPWR VPWR _23115_/X sky130_fd_sc_hd__or4_4
XANTENNA__17882__B1 _16952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24095_ _23916_/CLK _24095_/D HRESETn VGND VGND VPWR VPWR _24095_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_15_0_HCLK clkbuf_5_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_20258_ _21408_/B _20255_/X _19827_/A _20255_/X VGND VGND VPWR VPWR _23444_/D sky130_fd_sc_hd__a2bb2o_4
X_23046_ _21311_/X VGND VGND VPWR VPWR _23046_/X sky130_fd_sc_hd__buf_2
XFILLER_88_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19623__B2 _19598_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20189_ _20189_/A VGND VGND VPWR VPWR _20189_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24997_ _25005_/CLK _15352_/X HRESETn VGND VGND VPWR VPWR _24997_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_236_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14750_ _25061_/Q VGND VGND VPWR VPWR _21239_/A sky130_fd_sc_hd__inv_2
X_11962_ _11962_/A _11962_/B VGND VGND VPWR VPWR _11962_/X sky130_fd_sc_hd__and2_4
X_23948_ _25224_/CLK _20595_/X HRESETn VGND VGND VPWR VPWR _23948_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_1_1_HCLK clkbuf_1_1_0_HCLK/X VGND VGND VPWR VPWR clkbuf_2_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13701_ _13700_/X VGND VGND VPWR VPWR _13701_/X sky130_fd_sc_hd__buf_2
XFILLER_245_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14681_ _14681_/A VGND VGND VPWR VPWR _22219_/A sky130_fd_sc_hd__buf_2
XFILLER_45_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11893_ _11848_/B _11891_/Y _11892_/Y VGND VGND VPWR VPWR _11893_/X sky130_fd_sc_hd__o21a_4
X_23879_ _23844_/CLK _19036_/X VGND VGND VPWR VPWR _23879_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19139__B1 _19138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16420_ HWDATA[10] VGND VGND VPWR VPWR _16420_/X sky130_fd_sc_hd__buf_2
XFILLER_32_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24545__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13632_ _25298_/Q _13510_/X _13627_/X VGND VGND VPWR VPWR _13632_/X sky130_fd_sc_hd__a21o_4
XFILLER_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15963__A3 _16240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16351_ _16348_/Y _16344_/X _16349_/X _16350_/X VGND VGND VPWR VPWR _16351_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13563_ _13563_/A VGND VGND VPWR VPWR _13563_/Y sky130_fd_sc_hd__inv_2
X_15302_ _15130_/Y _15137_/Y _15302_/C _15301_/X VGND VGND VPWR VPWR _15320_/B sky130_fd_sc_hd__or4_4
XFILLER_12_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12514_ _12514_/A VGND VGND VPWR VPWR _12514_/Y sky130_fd_sc_hd__inv_2
X_19070_ _19069_/Y _19062_/X _18998_/X _19054_/A VGND VGND VPWR VPWR _23867_/D sky130_fd_sc_hd__a2bb2o_4
X_16282_ _16281_/Y _16279_/X _15554_/X _16279_/X VGND VGND VPWR VPWR _16282_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13494_ _13499_/A VGND VGND VPWR VPWR _13494_/X sky130_fd_sc_hd__buf_2
XFILLER_200_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16912__A2 _24277_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18021_ _18062_/A _18021_/B _18021_/C VGND VGND VPWR VPWR _18021_/X sky130_fd_sc_hd__and3_4
X_15233_ _15059_/X _15311_/B VGND VGND VPWR VPWR _15233_/X sky130_fd_sc_hd__or2_4
X_12445_ _12226_/X _12418_/X _12390_/X _12442_/B VGND VGND VPWR VPWR _12446_/A sky130_fd_sc_hd__a211o_4
XANTENNA__19311__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22997__A1 _24568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15164_ _14883_/Y _15162_/A VGND VGND VPWR VPWR _15164_/X sky130_fd_sc_hd__or2_4
XANTENNA__16125__B1 _11726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12376_ _12376_/A _12374_/A VGND VGND VPWR VPWR _12377_/C sky130_fd_sc_hd__or2_4
X_14115_ _14115_/A VGND VGND VPWR VPWR _14115_/X sky130_fd_sc_hd__buf_2
XFILLER_141_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15095_ _15093_/A _24588_/Q _15294_/B _15094_/Y VGND VGND VPWR VPWR _15095_/X sky130_fd_sc_hd__o22a_4
X_19972_ _19969_/Y _19963_/X _19970_/X _19971_/X VGND VGND VPWR VPWR _23552_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25333__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22749__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14046_ _14067_/A VGND VGND VPWR VPWR _14046_/X sky130_fd_sc_hd__buf_2
X_18923_ _18922_/Y _18918_/X _16783_/X _18918_/X VGND VGND VPWR VPWR _18923_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13437__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18854_ _16517_/Y _24133_/Q _16517_/Y _24133_/Q VGND VGND VPWR VPWR _18854_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14439__B1 _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17805_ _17744_/A _17804_/Y VGND VGND VPWR VPWR _17806_/C sky130_fd_sc_hd__or2_4
X_15997_ _15988_/X VGND VGND VPWR VPWR _15998_/A sky130_fd_sc_hd__buf_2
X_18785_ _18682_/D _18745_/C VGND VGND VPWR VPWR _18815_/B sky130_fd_sc_hd__or2_4
XFILLER_227_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19378__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15652__A _15648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14948_ _15063_/A VGND VGND VPWR VPWR _15204_/A sky130_fd_sc_hd__buf_2
X_17736_ _18313_/A _17736_/B _17736_/C _17735_/X VGND VGND VPWR VPWR _17736_/X sky130_fd_sc_hd__or4_4
XANTENNA__21373__B _21372_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_35_0_HCLK clkbuf_8_35_0_HCLK/A VGND VGND VPWR VPWR _23497_/CLK sky130_fd_sc_hd__clkbuf_1
X_14879_ pwm_S6 VGND VGND VPWR VPWR _14879_/Y sky130_fd_sc_hd__inv_2
X_17667_ _17530_/Y _17686_/A VGND VGND VPWR VPWR _17668_/B sky130_fd_sc_hd__or2_4
Xclkbuf_8_98_0_HCLK clkbuf_8_98_0_HCLK/A VGND VGND VPWR VPWR _24629_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_63_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24286__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19406_ _19405_/Y _19403_/X _19360_/X _19403_/X VGND VGND VPWR VPWR _23748_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16618_ _16617_/Y _16541_/X _16358_/X _16541_/X VGND VGND VPWR VPWR _24516_/D sky130_fd_sc_hd__a2bb2o_4
X_17598_ _17600_/B VGND VGND VPWR VPWR _17598_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22485__A _22429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24215__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16549_ _16546_/Y _16542_/X _16459_/X _16548_/X VGND VGND VPWR VPWR _24544_/D sky130_fd_sc_hd__a2bb2o_4
X_19337_ _19336_/Y _19334_/X _19203_/X _19334_/X VGND VGND VPWR VPWR _19337_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22685__B1 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16483__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19268_ _23796_/Q VGND VGND VPWR VPWR _19268_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16903__A2 _24276_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18219_ _18056_/A _18219_/B _18218_/X VGND VGND VPWR VPWR _18220_/C sky130_fd_sc_hd__and3_4
X_19199_ _19191_/A VGND VGND VPWR VPWR _19199_/X sky130_fd_sc_hd__buf_2
XFILLER_191_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19302__B1 _19301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21230_ _21018_/B _16268_/A _15651_/A _20822_/A _16270_/A VGND VGND VPWR VPWR _21230_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_191_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21829__A _21714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19853__B2 _19835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21161_ _14229_/Y _14209_/A _17433_/Y _21368_/A VGND VGND VPWR VPWR _21161_/X sky130_fd_sc_hd__o22a_4
XANTENNA__25074__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20112_ _20111_/Y _20105_/X _19852_/X _20088_/A VGND VGND VPWR VPWR _20112_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21092_ _21041_/X _21091_/Y _12728_/A _21041_/X VGND VGND VPWR VPWR _21092_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25003__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20043_ _20043_/A VGND VGND VPWR VPWR _20043_/Y sky130_fd_sc_hd__inv_2
X_24920_ _24032_/CLK _15565_/X HRESETn VGND VGND VPWR VPWR _15563_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_131_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24851_ _25390_/CLK _24851_/D HRESETn VGND VGND VPWR VPWR _24851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23802_ _23610_/CLK _23802_/D VGND VGND VPWR VPWR _23802_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24782_ _24819_/CLK _24782_/D HRESETn VGND VGND VPWR VPWR _21015_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_100_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ _17893_/A _20320_/Y _21991_/X _21993_/X VGND VGND VPWR VPWR _21994_/X sky130_fd_sc_hd__o22a_4
XPHY_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23733_ _23747_/CLK _19448_/X VGND VGND VPWR VPWR _19446_/A sky130_fd_sc_hd__dfxtp_4
XPHY_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ _13635_/A _20941_/X _20949_/B VGND VGND VPWR VPWR _20945_/Y sky130_fd_sc_hd__a21oi_4
XPHY_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14609__C _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ _23665_/CLK _23664_/D VGND VGND VPWR VPWR _19656_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_6_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _20870_/X _20872_/Y _24489_/Q _20875_/X VGND VGND VPWR VPWR _20876_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25403_ _25403_/CLK _25403_/D HRESETn VGND VGND VPWR VPWR _25403_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22615_ _16415_/A _22532_/B VGND VGND VPWR VPWR _22615_/X sky130_fd_sc_hd__or2_4
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23595_ _23525_/CLK _19853_/X VGND VGND VPWR VPWR _19851_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19541__B1 _19540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25334_ _24907_/CLK _13130_/X HRESETn VGND VGND VPWR VPWR _25334_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22546_ _22521_/B _22542_/X _22423_/X _22545_/X VGND VGND VPWR VPWR _22546_/X sky130_fd_sc_hd__o22a_4
XFILLER_195_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25265_ _25089_/CLK _25265_/D HRESETn VGND VGND VPWR VPWR _13567_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23938__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22477_ _22146_/X VGND VGND VPWR VPWR _22477_/X sky130_fd_sc_hd__buf_2
XFILLER_148_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12230_ _12275_/A VGND VGND VPWR VPWR _12418_/A sky130_fd_sc_hd__buf_2
X_24216_ _25285_/CLK _24216_/D HRESETn VGND VGND VPWR VPWR _19455_/B sky130_fd_sc_hd__dfrtp_4
X_21428_ _21030_/A VGND VGND VPWR VPWR _21428_/X sky130_fd_sc_hd__buf_2
XANTENNA__16107__B1 _11691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25196_ _25043_/CLK _14226_/X HRESETn VGND VGND VPWR VPWR _25196_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_205_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12161_ _12160_/X VGND VGND VPWR VPWR _12161_/Y sky130_fd_sc_hd__inv_2
X_24147_ _24340_/CLK _24147_/D HRESETn VGND VGND VPWR VPWR _24147_/Q sky130_fd_sc_hd__dfrtp_4
X_21359_ _18388_/Y _21571_/A _12154_/A _21570_/A VGND VGND VPWR VPWR _21359_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23376__D HSEL VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12092_ _25477_/Q VGND VGND VPWR VPWR _12092_/Y sky130_fd_sc_hd__inv_2
X_24078_ _24959_/CLK _20481_/X HRESETn VGND VGND VPWR VPWR _20525_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15920_ _19646_/A VGND VGND VPWR VPWR _15920_/X sky130_fd_sc_hd__buf_2
X_23029_ _12812_/Y _21437_/X _22280_/X _12574_/Y _21085_/X VGND VGND VPWR VPWR _23029_/X
+ sky130_fd_sc_hd__o32a_4
XANTENNA__22600__B1 _24727_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25140__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15851_ _15845_/A VGND VGND VPWR VPWR _15851_/X sky130_fd_sc_hd__buf_2
XFILLER_237_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24797__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14802_ _20628_/A _14802_/B _14802_/C VGND VGND VPWR VPWR _14803_/A sky130_fd_sc_hd__or3_4
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22289__B _22416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24726__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15782_ _15918_/B VGND VGND VPWR VPWR _15813_/A sky130_fd_sc_hd__inv_2
X_18570_ _18473_/Y _18568_/X _18569_/Y VGND VGND VPWR VPWR _24169_/D sky130_fd_sc_hd__o21a_4
XFILLER_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_251_0_HCLK clkbuf_8_251_0_HCLK/A VGND VGND VPWR VPWR _23972_/CLK sky130_fd_sc_hd__clkbuf_1
X_12994_ _12970_/X _12992_/X _12994_/C VGND VGND VPWR VPWR _25366_/D sky130_fd_sc_hd__and3_4
XFILLER_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21167__B1 _11701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14733_ _14721_/X _14725_/Y VGND VGND VPWR VPWR _14733_/Y sky130_fd_sc_hd__nor2_4
X_17521_ _17521_/A VGND VGND VPWR VPWR _17521_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11945_ _11945_/A VGND VGND VPWR VPWR _11945_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ _17452_/A VGND VGND VPWR VPWR _20387_/A sky130_fd_sc_hd__inv_2
X_14664_ _14664_/A _17703_/B _13584_/X _21283_/A VGND VGND VPWR VPWR _14664_/X sky130_fd_sc_hd__or4_4
XFILLER_221_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11876_ _11875_/X VGND VGND VPWR VPWR _11876_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16403_ _15117_/Y _16398_/X _16402_/X _16398_/X VGND VGND VPWR VPWR _24597_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13615_ _13615_/A VGND VGND VPWR VPWR _19117_/A sky130_fd_sc_hd__buf_2
X_17383_ _17399_/A VGND VGND VPWR VPWR _17384_/A sky130_fd_sc_hd__inv_2
X_14595_ _13560_/Y _14550_/X VGND VGND VPWR VPWR _14595_/Y sky130_fd_sc_hd__nand2_4
XFILLER_186_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19532__B1 _19395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16334_ _24622_/Q VGND VGND VPWR VPWR _16334_/Y sky130_fd_sc_hd__inv_2
X_19122_ _18981_/A VGND VGND VPWR VPWR _19122_/X sky130_fd_sc_hd__buf_2
X_13546_ _25088_/Q VGND VGND VPWR VPWR _14553_/A sky130_fd_sc_hd__inv_2
XFILLER_187_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19053_ _23872_/Q VGND VGND VPWR VPWR _19053_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16265_ _16265_/A VGND VGND VPWR VPWR _16265_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13477_ _13475_/Y _13476_/X _11786_/X _13476_/X VGND VGND VPWR VPWR _13477_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25514__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15216_ _14921_/X _15214_/X _15215_/Y VGND VGND VPWR VPWR _25027_/D sky130_fd_sc_hd__o21a_4
X_18004_ _18057_/A VGND VGND VPWR VPWR _18004_/X sky130_fd_sc_hd__buf_2
XFILLER_173_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12428_ _12187_/Y _12428_/B _12428_/C _12428_/D VGND VGND VPWR VPWR _12428_/X sky130_fd_sc_hd__or4_4
X_16196_ _16195_/Y _16191_/X _16004_/X _16191_/X VGND VGND VPWR VPWR _24674_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12383__A1 _12254_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15147_ _15138_/X _15141_/X _15143_/X _15147_/D VGND VGND VPWR VPWR _15157_/C sky130_fd_sc_hd__or4_4
X_12359_ _12350_/X _12359_/B _12355_/X _12358_/X VGND VGND VPWR VPWR _12359_/X sky130_fd_sc_hd__or4_4
XFILLER_153_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15078_ _24992_/Q VGND VGND VPWR VPWR _15078_/Y sky130_fd_sc_hd__inv_2
X_19955_ _23556_/Q VGND VGND VPWR VPWR _19955_/Y sky130_fd_sc_hd__inv_2
X_14029_ _13978_/X _14029_/B _13980_/X _14019_/D VGND VGND VPWR VPWR _14029_/X sky130_fd_sc_hd__or4_4
X_18906_ _17517_/Y _11794_/X HWDATA[29] _11794_/X VGND VGND VPWR VPWR _24112_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17862__A _17849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19886_ _23583_/Q VGND VGND VPWR VPWR _19886_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_61_0_HCLK clkbuf_5_30_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_61_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18837_ _24576_/Q _24155_/Q _16458_/Y _18707_/A VGND VGND VPWR VPWR _18840_/B sky130_fd_sc_hd__o22a_4
XFILLER_228_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24467__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18768_ _18770_/B VGND VGND VPWR VPWR _18768_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16499__A1_N _16498_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17719_ _21924_/A VGND VGND VPWR VPWR _17720_/A sky130_fd_sc_hd__buf_2
XFILLER_236_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18699_ _18745_/C _18706_/A VGND VGND VPWR VPWR _18699_/X sky130_fd_sc_hd__or2_4
XANTENNA__18693__A _18760_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20730_ _20729_/X VGND VGND VPWR VPWR _24012_/D sky130_fd_sc_hd__inv_2
XANTENNA__15927__A3 _15702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_211_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20661_ _17394_/X _20660_/Y _20661_/C VGND VGND VPWR VPWR _20661_/X sky130_fd_sc_hd__and3_4
XFILLER_196_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22122__A2 _21721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22400_ _22400_/A _22396_/B VGND VGND VPWR VPWR _22400_/X sky130_fd_sc_hd__or2_4
XFILLER_51_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20592_ _20592_/A _18888_/A VGND VGND VPWR VPWR _20595_/B sky130_fd_sc_hd__or2_4
X_23380_ _23806_/CLK _23380_/D VGND VGND VPWR VPWR _20419_/A sky130_fd_sc_hd__dfxtp_4
X_22331_ _22331_/A VGND VGND VPWR VPWR _22331_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21881__A1 _25437_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16888__B2 _23320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22662__B _22661_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25050_ _25050_/CLK _25050_/D HRESETn VGND VGND VPWR VPWR _14811_/A sky130_fd_sc_hd__dfrtp_4
X_22262_ _22262_/A _22262_/B VGND VGND VPWR VPWR _22263_/C sky130_fd_sc_hd__or2_4
XFILLER_247_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24001_ _25226_/CLK _20508_/X HRESETn VGND VGND VPWR VPWR _24001_/Q sky130_fd_sc_hd__dfrtp_4
X_21213_ _21178_/X _21196_/X _21212_/X VGND VGND VPWR VPWR _21213_/X sky130_fd_sc_hd__and3_4
XANTENNA__15557__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22193_ _25526_/Q _22417_/B _21118_/X _22192_/X VGND VGND VPWR VPWR _22193_/X sky130_fd_sc_hd__a211o_4
XFILLER_144_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23196__D _23195_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21144_ _12163_/A _12082_/A _12032_/Y _12082_/A VGND VGND VPWR VPWR _21144_/X sky130_fd_sc_hd__a2bb2o_4
X_21075_ _15780_/B VGND VGND VPWR VPWR _21075_/Y sky130_fd_sc_hd__inv_2
X_20026_ _21658_/B _20025_/X _19981_/X _20025_/X VGND VGND VPWR VPWR _23533_/D sky130_fd_sc_hd__a2bb2o_4
X_24903_ _24903_/CLK _15609_/X HRESETn VGND VGND VPWR VPWR _15607_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21294__A _21864_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24890__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24834_ _24834_/CLK _24834_/D HRESETn VGND VGND VPWR VPWR _24834_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13626__A1 _13525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21149__B1 _21568_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24137__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24765_ _24765_/CLK _24765_/D HRESETn VGND VGND VPWR VPWR _24765_/Q sky130_fd_sc_hd__dfrtp_4
X_21977_ _21962_/A _21977_/B VGND VGND VPWR VPWR _21977_/Y sky130_fd_sc_hd__nand2_4
XPHY_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _16226_/A VGND VGND VPWR VPWR _11730_/X sky130_fd_sc_hd__buf_2
X_23716_ _23427_/CLK _19497_/X VGND VGND VPWR VPWR _23716_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ _13651_/A VGND VGND VPWR VPWR _20928_/Y sky130_fd_sc_hd__inv_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21741__B _21741_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24696_ _24696_/CLK _16127_/X HRESETn VGND VGND VPWR VPWR _22753_/A sky130_fd_sc_hd__dfrtp_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_81_0_HCLK clkbuf_7_40_0_HCLK/X VGND VGND VPWR VPWR _25382_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _14177_/A VGND VGND VPWR VPWR _15541_/A sky130_fd_sc_hd__inv_2
X_23647_ _23644_/CLK _23647_/D VGND VGND VPWR VPWR _13311_/B sky130_fd_sc_hd__dfxtp_4
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20859_ _16699_/Y _20846_/X _20855_/X _20858_/X VGND VGND VPWR VPWR _20859_/X sky130_fd_sc_hd__o22a_4
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _13193_/A _13400_/B _13399_/X VGND VGND VPWR VPWR _13401_/C sky130_fd_sc_hd__and3_4
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ _14380_/A VGND VGND VPWR VPWR _14380_/X sky130_fd_sc_hd__buf_2
XANTENNA__16328__B1 _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23578_ _24199_/CLK _23578_/D VGND VGND VPWR VPWR _19897_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__19947__A1_N _19945_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ _13363_/A _13331_/B VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__or2_4
X_25317_ _25479_/CLK _25317_/D HRESETn VGND VGND VPWR VPWR _13480_/A sky130_fd_sc_hd__dfrtp_4
X_22529_ _22498_/X _22502_/X _22508_/Y _22528_/X VGND VGND VPWR VPWR HRDATA[9] sky130_fd_sc_hd__a211o_4
XFILLER_127_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21872__A1 _24789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_HCLK clkbuf_1_0_1_HCLK/X VGND VGND VPWR VPWR clkbuf_3_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21872__B2 _21871_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16050_ _16038_/A VGND VGND VPWR VPWR _16050_/X sky130_fd_sc_hd__buf_2
X_13262_ _13369_/A _13262_/B _13261_/X VGND VGND VPWR VPWR _13262_/X sky130_fd_sc_hd__or3_4
X_25248_ _25249_/CLK _13864_/X HRESETn VGND VGND VPWR VPWR _25248_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15001_ _25037_/Q _24475_/Q _15168_/A _15000_/Y VGND VGND VPWR VPWR _15007_/B sky130_fd_sc_hd__o22a_4
XFILLER_136_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12213_ _25435_/Q _21534_/A _12211_/Y _12212_/Y VGND VGND VPWR VPWR _12213_/X sky130_fd_sc_hd__o22a_4
XFILLER_157_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13193_ _13193_/A _13193_/B _13193_/C VGND VGND VPWR VPWR _13202_/B sky130_fd_sc_hd__and3_4
X_25179_ _25171_/CLK _25179_/D HRESETn VGND VGND VPWR VPWR _14278_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_151_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12144_ _12080_/Y _12143_/X _12080_/Y _12143_/X VGND VGND VPWR VPWR _12144_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24978__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19740_ _19740_/A VGND VGND VPWR VPWR _19740_/X sky130_fd_sc_hd__buf_2
XANTENNA__24907__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12075_ HWDATA[1] VGND VGND VPWR VPWR _14262_/A sky130_fd_sc_hd__buf_2
X_16952_ _17791_/A VGND VGND VPWR VPWR _16952_/X sky130_fd_sc_hd__buf_2
XFILLER_1_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15903_ _15701_/X _15887_/X _15838_/X _24785_/Q _15857_/A VGND VGND VPWR VPWR _24785_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__18253__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19671_ _20052_/A _20220_/D _19094_/C VGND VGND VPWR VPWR _19672_/A sky130_fd_sc_hd__or3_4
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16883_ _16881_/Y _16877_/X _16882_/X _16877_/X VGND VGND VPWR VPWR _24407_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24560__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18622_ _16600_/A _24134_/Q _16600_/Y _18783_/A VGND VGND VPWR VPWR _18622_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15834_ _12332_/Y _15827_/X _14479_/X _15792_/X VGND VGND VPWR VPWR _15834_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_237_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21932__A _21936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18553_ _18479_/B _18553_/B VGND VGND VPWR VPWR _18556_/B sky130_fd_sc_hd__or2_4
XANTENNA__16448__D _21327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12977_ _12324_/Y _13046_/A _12976_/X VGND VGND VPWR VPWR _12977_/X sky130_fd_sc_hd__or3_4
X_15765_ _15745_/X _15761_/X _15764_/X _24858_/Q _15706_/X VGND VGND VPWR VPWR _15765_/X
+ sky130_fd_sc_hd__a32o_4
X_17504_ _25541_/Q _17502_/Y _17494_/A _17503_/Y VGND VGND VPWR VPWR _17504_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15930__A _15924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11928_ _11926_/Y _11919_/X _11927_/X _11897_/X VGND VGND VPWR VPWR _25503_/D sky130_fd_sc_hd__a2bb2o_4
X_14716_ _13731_/X _14699_/B _21787_/A VGND VGND VPWR VPWR _14716_/X sky130_fd_sc_hd__and3_4
XFILLER_73_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15696_ _16364_/A _14178_/B _15636_/C _15984_/D VGND VGND VPWR VPWR _15697_/B sky130_fd_sc_hd__or4_4
X_18484_ _18457_/Y _18483_/X VGND VGND VPWR VPWR _18484_/Y sky130_fd_sc_hd__nor2_4
XFILLER_205_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21560__B1 _14863_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14647_ _13612_/A _14647_/B VGND VGND VPWR VPWR _14784_/A sky130_fd_sc_hd__or2_4
X_17435_ _21012_/A VGND VGND VPWR VPWR _17435_/Y sky130_fd_sc_hd__inv_2
X_11859_ _11802_/Y _11851_/X _11799_/X _11854_/X _11858_/Y VGND VGND VPWR VPWR _11864_/B
+ sky130_fd_sc_hd__a2111o_4
Xclkbuf_8_109_0_HCLK clkbuf_7_54_0_HCLK/X VGND VGND VPWR VPWR _24645_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_33_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12565__A2_N _24870_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14578_ _25093_/Q _14559_/B VGND VGND VPWR VPWR _14578_/X sky130_fd_sc_hd__or2_4
X_17366_ _17366_/A _17366_/B VGND VGND VPWR VPWR _17366_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__22655__A3 _22138_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19105_ _23854_/Q VGND VGND VPWR VPWR _19105_/Y sky130_fd_sc_hd__inv_2
X_13529_ _17914_/A _13528_/X VGND VGND VPWR VPWR _15904_/B sky130_fd_sc_hd__and2_4
X_16317_ _24628_/Q VGND VGND VPWR VPWR _16317_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17297_ _17288_/X VGND VGND VPWR VPWR _17301_/B sky130_fd_sc_hd__inv_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16248_ _16247_/Y _16245_/X _16145_/X _16245_/X VGND VGND VPWR VPWR _24655_/D sky130_fd_sc_hd__a2bb2o_4
X_19036_ _19035_/Y _19033_/X _18942_/X _19033_/X VGND VGND VPWR VPWR _19036_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17167__A1_N _24618_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16179_ _16179_/A VGND VGND VPWR VPWR _16180_/A sky130_fd_sc_hd__buf_2
XFILLER_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22812__B1 _22793_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18688__A _24138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24648__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19938_ _23562_/Q VGND VGND VPWR VPWR _22346_/B sky130_fd_sc_hd__inv_2
XANTENNA__22040__A1 _22393_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22040__B2 _22039_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19869_ _19856_/Y VGND VGND VPWR VPWR _19869_/X sky130_fd_sc_hd__buf_2
XFILLER_228_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21900_ _21895_/X _21899_/X _22212_/A VGND VGND VPWR VPWR _21900_/X sky130_fd_sc_hd__o21a_4
XANTENNA__22591__A2 _22432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22880_ _23060_/A _22880_/B VGND VGND VPWR VPWR _22880_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__12518__A2_N _24855_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16001__A HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17735__A1_N _17731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24230__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21831_ _21830_/Y _21319_/X _16706_/A _11706_/X VGND VGND VPWR VPWR _21831_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19744__B1 _19743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24550_ _24555_/CLK _24550_/D HRESETn VGND VGND VPWR VPWR _16530_/A sky130_fd_sc_hd__dfrtp_4
X_21762_ _14678_/X _21762_/B VGND VGND VPWR VPWR _21762_/X sky130_fd_sc_hd__or2_4
XANTENNA__16558__B1 _16295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_68_0_HCLK clkbuf_7_69_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_68_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23501_ _23378_/CLK _23501_/D VGND VGND VPWR VPWR _23501_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20713_ _13116_/A _13116_/B _13117_/B VGND VGND VPWR VPWR _20713_/Y sky130_fd_sc_hd__a21boi_4
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24481_ _24594_/CLK _24481_/D HRESETn VGND VGND VPWR VPWR _24481_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21693_ _17704_/C _21649_/X VGND VGND VPWR VPWR _21693_/Y sky130_fd_sc_hd__nor2_4
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23432_ _23441_/CLK _20291_/X VGND VGND VPWR VPWR _20290_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20644_ _17399_/X VGND VGND VPWR VPWR _20661_/C sky130_fd_sc_hd__buf_2
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22673__A _16503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23363_ _23363_/A VGND VGND VPWR VPWR IRQ[19] sky130_fd_sc_hd__buf_2
XANTENNA__17767__A _17555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20575_ _20575_/A VGND VGND VPWR VPWR _20575_/Y sky130_fd_sc_hd__inv_2
X_25102_ _23958_/CLK _14522_/X HRESETn VGND VGND VPWR VPWR _25102_/Q sky130_fd_sc_hd__dfrtp_4
X_22314_ _14362_/Y _14182_/A _14461_/Y _21155_/B VGND VGND VPWR VPWR _22314_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21289__A _21119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23294_ _23235_/A _23294_/B VGND VGND VPWR VPWR _23294_/Y sky130_fd_sc_hd__nor2_4
XFILLER_191_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25033_ _25021_/CLK _25033_/D HRESETn VGND VGND VPWR VPWR _25033_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15287__A _15331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12347__B2 _24835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22245_ _22007_/X _22243_/X _22244_/X VGND VGND VPWR VPWR _22245_/X sky130_fd_sc_hd__and3_4
XFILLER_145_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22176_ _21832_/A _22175_/X VGND VGND VPWR VPWR _22176_/X sky130_fd_sc_hd__and2_4
XANTENNA__24389__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21127_ _15981_/A VGND VGND VPWR VPWR _21127_/X sky130_fd_sc_hd__buf_2
XFILLER_132_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24920__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24318__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21058_ _21111_/A VGND VGND VPWR VPWR _21058_/X sky130_fd_sc_hd__buf_2
XFILLER_101_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12900_ _12838_/A _12838_/B _12741_/X _12892_/B VGND VGND VPWR VPWR _12906_/B sky130_fd_sc_hd__or4_4
XFILLER_59_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20009_ _21206_/B _20003_/X _20008_/X _19990_/Y VGND VGND VPWR VPWR _23539_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13880_ _13922_/A _13914_/A _13879_/X VGND VGND VPWR VPWR _13880_/X sky130_fd_sc_hd__or3_4
XFILLER_219_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16797__B1 _15710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21790__B1 _13772_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12831_ _25378_/Q VGND VGND VPWR VPWR _12834_/C sky130_fd_sc_hd__inv_2
X_24817_ _24819_/CLK _24817_/D HRESETn VGND VGND VPWR VPWR _12968_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_234_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15550_ _15550_/A VGND VGND VPWR VPWR _15550_/Y sky130_fd_sc_hd__inv_2
X_12762_ _12762_/A VGND VGND VPWR VPWR _12762_/Y sky130_fd_sc_hd__inv_2
X_24748_ _24800_/CLK _24748_/D HRESETn VGND VGND VPWR VPWR _21088_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16959__A1_N _16009_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16549__B1 _16459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14490_/B VGND VGND VPWR VPWR _14501_/Y sky130_fd_sc_hd__inv_2
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _25539_/Q VGND VGND VPWR VPWR _11713_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _24069_/Q _15478_/Y _15480_/Y _14542_/Y VGND VGND VPWR VPWR _15482_/B sky130_fd_sc_hd__a211o_4
XFILLER_230_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23953__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12692_/X VGND VGND VPWR VPWR _12693_/X sky130_fd_sc_hd__or2_4
X_24679_ _24679_/CLK _16176_/X HRESETn VGND VGND VPWR VPWR _14755_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_242_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14366__A _14366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14430_/Y _14426_/X _14407_/X _14431_/X VGND VGND VPWR VPWR _14432_/X sky130_fd_sc_hd__a2bb2o_4
X_17220_ _16303_/A _17219_/Y _16308_/Y _24361_/Q VGND VGND VPWR VPWR _17220_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_230_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25106__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17151_ _17041_/C _17124_/X VGND VGND VPWR VPWR _17151_/X sky130_fd_sc_hd__or2_4
XFILLER_168_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _14362_/Y VGND VGND VPWR VPWR _20467_/A sky130_fd_sc_hd__buf_2
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16102_ _16101_/Y _16099_/X _11685_/X _16099_/X VGND VGND VPWR VPWR _16102_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_167_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13314_ _13422_/A VGND VGND VPWR VPWR _13314_/X sky130_fd_sc_hd__buf_2
XFILLER_167_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17082_ _17024_/A _17085_/B VGND VGND VPWR VPWR _17083_/C sky130_fd_sc_hd__or2_4
XFILLER_6_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14294_ _14294_/A VGND VGND VPWR VPWR _14295_/A sky130_fd_sc_hd__inv_2
XFILLER_182_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16033_ _16038_/A VGND VGND VPWR VPWR _16033_/X sky130_fd_sc_hd__buf_2
XANTENNA__12338__B2 _24834_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13245_ _13184_/A VGND VGND VPWR VPWR _13245_/X sky130_fd_sc_hd__buf_2
XFILLER_171_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17277__A1 _17231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13176_ _13172_/A _13176_/B _13176_/C VGND VGND VPWR VPWR _13176_/X sky130_fd_sc_hd__and3_4
XFILLER_124_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12127_ _12126_/X VGND VGND VPWR VPWR _12127_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15925__A _15924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24741__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17984_ _18090_/A VGND VGND VPWR VPWR _17984_/X sky130_fd_sc_hd__buf_2
XFILLER_96_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24059__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19723_ _19723_/A VGND VGND VPWR VPWR _19723_/X sky130_fd_sc_hd__buf_2
X_12058_ _16181_/A _12058_/B _12058_/C _12057_/X VGND VGND VPWR VPWR _12058_/X sky130_fd_sc_hd__or4_4
X_16935_ _16108_/Y _24280_/Q _22564_/A _16895_/X VGND VGND VPWR VPWR _16942_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22573__A2 _22435_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19654_ _13221_/B VGND VGND VPWR VPWR _19654_/Y sky130_fd_sc_hd__inv_2
X_16866_ _16863_/Y _16856_/X _16864_/X _16865_/X VGND VGND VPWR VPWR _24411_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16788__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18605_ _24151_/Q VGND VGND VPWR VPWR _18732_/A sky130_fd_sc_hd__buf_2
X_15817_ _15810_/X _15813_/X _15746_/X _24832_/Q _15811_/X VGND VGND VPWR VPWR _24832_/D
+ sky130_fd_sc_hd__a32o_4
X_19585_ _23686_/Q VGND VGND VPWR VPWR _19585_/X sky130_fd_sc_hd__buf_2
X_16797_ _16796_/Y _16794_/X _15710_/X _16794_/X VGND VGND VPWR VPWR _16797_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19726__B1 _19702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15660__A _15660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18536_ _18407_/Y _18541_/B _18489_/X VGND VGND VPWR VPWR _18536_/Y sky130_fd_sc_hd__a21oi_4
X_15748_ HWDATA[11] VGND VGND VPWR VPWR _15748_/X sky130_fd_sc_hd__buf_2
XFILLER_61_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18467_ _18467_/A _18467_/B _18466_/X VGND VGND VPWR VPWR _18468_/C sky130_fd_sc_hd__or3_4
X_15679_ _15678_/X VGND VGND VPWR VPWR _15679_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17418_ _14403_/A VGND VGND VPWR VPWR _17418_/X sky130_fd_sc_hd__buf_2
XANTENNA__22089__A1 _14710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18398_ _18393_/X _18394_/X _18398_/C _18397_/X VGND VGND VPWR VPWR _18398_/X sky130_fd_sc_hd__or4_4
XANTENNA__22493__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17349_ _24352_/Q _17349_/B VGND VGND VPWR VPWR _17351_/B sky130_fd_sc_hd__or2_4
XFILLER_193_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20360_ _21806_/B _20355_/X _19613_/A _20355_/X VGND VGND VPWR VPWR _23405_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_228_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16712__B1 _16435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19019_ _19017_/Y _19018_/X _18948_/X _19018_/X VGND VGND VPWR VPWR _19019_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24829__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20291_ _22244_/B _20288_/X _19967_/X _20288_/X VGND VGND VPWR VPWR _20291_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_228_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22940__B _22817_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22797__C1 _22520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22030_ _22016_/A _19605_/Y VGND VGND VPWR VPWR _22030_/X sky130_fd_sc_hd__or2_4
XFILLER_103_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24482__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24411__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23981_ _23986_/CLK _23981_/D HRESETn VGND VGND VPWR VPWR _20643_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_229_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12501__B2 _24886_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_31_0_HCLK clkbuf_5_31_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_63_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22932_ _22932_/A VGND VGND VPWR VPWR _23177_/B sky130_fd_sc_hd__buf_2
XFILLER_29_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22863_ _23043_/A _22863_/B VGND VGND VPWR VPWR _22873_/C sky130_fd_sc_hd__and2_4
XFILLER_243_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24602_ _24520_/CLK _24602_/D HRESETn VGND VGND VPWR VPWR _24602_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15570__A _15553_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21814_ _21487_/A _21814_/B VGND VGND VPWR VPWR _21814_/X sky130_fd_sc_hd__or2_4
XFILLER_37_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22794_ _22794_/A VGND VGND VPWR VPWR _22794_/X sky130_fd_sc_hd__buf_2
XFILLER_243_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21524__B1 _25522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24533_ _24573_/CLK _24533_/D HRESETn VGND VGND VPWR VPWR _16574_/A sky130_fd_sc_hd__dfrtp_4
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21745_ _16708_/Y _21745_/B VGND VGND VPWR VPWR _21745_/X sky130_fd_sc_hd__and2_4
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24464_ _24463_/CLK _24464_/D HRESETn VGND VGND VPWR VPWR _24464_/Q sky130_fd_sc_hd__dfrtp_4
X_21676_ _21809_/A _21676_/B VGND VGND VPWR VPWR _21676_/X sky130_fd_sc_hd__or2_4
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23415_ _23415_/CLK _23415_/D VGND VGND VPWR VPWR _20333_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20627_ _20627_/A VGND VGND VPWR VPWR _20627_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_155_0_HCLK clkbuf_7_77_0_HCLK/X VGND VGND VPWR VPWR _25164_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24395_ _24390_/CLK _17086_/Y HRESETn VGND VGND VPWR VPWR _24395_/Q sky130_fd_sc_hd__dfrtp_4
X_23346_ _23346_/A _23346_/B VGND VGND VPWR VPWR _23346_/Y sky130_fd_sc_hd__nor2_4
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20558_ _20558_/A _20553_/A VGND VGND VPWR VPWR _20559_/B sky130_fd_sc_hd__nand2_4
XFILLER_192_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13517__B1 SCLK_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23277_ _23277_/A _23277_/B VGND VGND VPWR VPWR _23277_/X sky130_fd_sc_hd__and2_4
X_20489_ _20496_/A _20489_/B _20503_/C VGND VGND VPWR VPWR _20490_/B sky130_fd_sc_hd__and3_4
XFILLER_106_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13030_ _13087_/A VGND VGND VPWR VPWR _13048_/A sky130_fd_sc_hd__buf_2
X_25016_ _24967_/CLK _25016_/D HRESETn VGND VGND VPWR VPWR _25016_/Q sky130_fd_sc_hd__dfrtp_4
X_22228_ _22228_/A _22228_/B _22228_/C VGND VGND VPWR VPWR _22228_/X sky130_fd_sc_hd__and3_4
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15745__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22159_ _15072_/A _22932_/A VGND VGND VPWR VPWR _22162_/B sky130_fd_sc_hd__or2_4
XANTENNA__24152__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14981_ _14981_/A VGND VGND VPWR VPWR _14982_/A sky130_fd_sc_hd__inv_2
XFILLER_75_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19956__B1 _19620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16720_ _22844_/A VGND VGND VPWR VPWR _22539_/A sky130_fd_sc_hd__buf_2
XFILLER_219_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13932_ _13924_/A _13932_/B _13932_/C _13940_/A VGND VGND VPWR VPWR _13932_/X sky130_fd_sc_hd__or4_4
XFILLER_208_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13863_ _25248_/Q _13850_/X _21723_/A _13852_/X VGND VGND VPWR VPWR _13863_/X sky130_fd_sc_hd__o22a_4
X_16651_ _16650_/Y _16648_/X _16467_/X _16648_/X VGND VGND VPWR VPWR _16651_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16576__A _16576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22307__A2 _22807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25358__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12814_ _25390_/Q _12812_/Y _12813_/Y _24805_/Q VGND VGND VPWR VPWR _12814_/X sky130_fd_sc_hd__a2bb2o_4
X_15602_ _22683_/A _15596_/X _11739_/X _15601_/X VGND VGND VPWR VPWR _15602_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15480__A HTRANS[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19370_ _19369_/Y _19367_/X _19279_/X _19367_/X VGND VGND VPWR VPWR _23761_/D sky130_fd_sc_hd__a2bb2o_4
X_13794_ _25272_/Q VGND VGND VPWR VPWR _13794_/Y sky130_fd_sc_hd__inv_2
X_16582_ _16582_/A VGND VGND VPWR VPWR _16582_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18321_ _17703_/X _17706_/X _18320_/X VGND VGND VPWR VPWR _18322_/A sky130_fd_sc_hd__or3_4
X_12745_ _25378_/Q _12743_/Y _12744_/Y _24811_/Q VGND VGND VPWR VPWR _12745_/X sky130_fd_sc_hd__a2bb2o_4
X_15533_ _15530_/A VGND VGND VPWR VPWR _15533_/X sky130_fd_sc_hd__buf_2
XFILLER_187_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14096__A _14096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_51_0_HCLK clkbuf_7_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15464_ _15462_/Y _15458_/X _14407_/X _15463_/X VGND VGND VPWR VPWR _15464_/X sky130_fd_sc_hd__a2bb2o_4
X_18252_ _18234_/Y VGND VGND VPWR VPWR _18252_/X sky130_fd_sc_hd__buf_2
X_12676_ _12676_/A _12675_/Y VGND VGND VPWR VPWR _12677_/C sky130_fd_sc_hd__or2_4
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _14408_/A VGND VGND VPWR VPWR _14415_/X sky130_fd_sc_hd__buf_2
X_17203_ _17203_/A VGND VGND VPWR VPWR _17203_/X sky130_fd_sc_hd__buf_2
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__B2 _24868_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22744__C _22743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15395_ _15106_/Y _15395_/B VGND VGND VPWR VPWR _15395_/Y sky130_fd_sc_hd__nand2_4
X_18183_ _18151_/A _23876_/Q VGND VGND VPWR VPWR _18183_/X sky130_fd_sc_hd__or2_4
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ MSO_S3 _14345_/X _25160_/Q _14340_/X VGND VGND VPWR VPWR _14346_/Y sky130_fd_sc_hd__a22oi_4
X_17134_ _17038_/C _17132_/X _17133_/Y VGND VGND VPWR VPWR _24384_/D sky130_fd_sc_hd__o21a_4
XANTENNA__24993__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22491__B2 _22490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_195_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17065_ _17022_/A _17063_/X _17064_/X _17058_/Y VGND VGND VPWR VPWR _17066_/A sky130_fd_sc_hd__a211o_4
XFILLER_143_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24922__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14277_ _14289_/A VGND VGND VPWR VPWR _14285_/A sky130_fd_sc_hd__inv_2
XFILLER_171_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16016_ _24738_/Q VGND VGND VPWR VPWR _16016_/Y sky130_fd_sc_hd__inv_2
X_13228_ _13227_/X _13228_/B VGND VGND VPWR VPWR _13228_/X sky130_fd_sc_hd__or2_4
XFILLER_170_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17854__B _17849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12731__B2 _24796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13159_ _13175_/A _23618_/Q VGND VGND VPWR VPWR _13159_/X sky130_fd_sc_hd__or2_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18031__A _17999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17967_ _14628_/A VGND VGND VPWR VPWR _18220_/A sky130_fd_sc_hd__buf_2
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22546__A2 _22542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19706_ _19706_/A VGND VGND VPWR VPWR _19706_/Y sky130_fd_sc_hd__inv_2
X_16918_ _21521_/A _16917_/A _16159_/Y _16917_/Y VGND VGND VPWR VPWR _16918_/X sky130_fd_sc_hd__o22a_4
XFILLER_78_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17898_ _21993_/A _17910_/B VGND VGND VPWR VPWR _17898_/Y sky130_fd_sc_hd__nand2_4
XFILLER_238_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19637_ _19636_/Y _19634_/X _19534_/X _19634_/X VGND VGND VPWR VPWR _23671_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16849_ _19063_/A VGND VGND VPWR VPWR _16849_/X sky130_fd_sc_hd__buf_2
XFILLER_53_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19568_ _23690_/Q VGND VGND VPWR VPWR _19568_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25028__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18519_ _18497_/A _18515_/B _18518_/X VGND VGND VPWR VPWR _24181_/D sky130_fd_sc_hd__and3_4
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13622__B _13586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19499_ _21197_/B _19494_/X _19475_/X _19494_/A VGND VGND VPWR VPWR _23715_/D sky130_fd_sc_hd__a2bb2o_4
X_21530_ _22716_/A _21530_/B VGND VGND VPWR VPWR _21530_/X sky130_fd_sc_hd__and2_4
XFILLER_167_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16933__B1 _16126_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21461_ _21207_/A VGND VGND VPWR VPWR _21462_/A sky130_fd_sc_hd__buf_2
XFILLER_194_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_228_0_HCLK clkbuf_8_229_0_HCLK/A VGND VGND VPWR VPWR _25005_/CLK sky130_fd_sc_hd__clkbuf_1
X_23200_ _16650_/Y _23291_/B VGND VGND VPWR VPWR _23200_/X sky130_fd_sc_hd__and2_4
X_20412_ _20412_/A VGND VGND VPWR VPWR _22217_/B sky130_fd_sc_hd__inv_2
X_24180_ _24675_/CLK _18522_/Y HRESETn VGND VGND VPWR VPWR _24180_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_239_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21392_ _25061_/Q VGND VGND VPWR VPWR _22197_/A sky130_fd_sc_hd__buf_2
XFILLER_146_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23131_ _23169_/A _23131_/B VGND VGND VPWR VPWR _23131_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24663__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20343_ _23411_/Q VGND VGND VPWR VPWR _20343_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14172__B1 _14171_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23062_ _23062_/A _23061_/X VGND VGND VPWR VPWR _23072_/B sky130_fd_sc_hd__nor2_4
XANTENNA__21567__A _21730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20274_ _23438_/Q VGND VGND VPWR VPWR _21921_/B sky130_fd_sc_hd__inv_2
XFILLER_89_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17764__B _16940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22013_ _22024_/A _22010_/X _22012_/X VGND VGND VPWR VPWR _22013_/X sky130_fd_sc_hd__and3_4
XFILLER_161_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21286__B _21224_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13085__A _13085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17780__A _16913_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23964_ _24146_/CLK _20483_/X HRESETn VGND VGND VPWR VPWR _23964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_245_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22915_ _12201_/Y _22499_/X _24277_/Q _22914_/X VGND VGND VPWR VPWR _22915_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23895_ _23844_/CLK _18989_/X VGND VGND VPWR VPWR _23895_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16620__A2_N _16541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22846_ _21868_/X VGND VGND VPWR VPWR _22846_/X sky130_fd_sc_hd__buf_2
XANTENNA__15975__A1 _15784_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15975__B2 _15925_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22777_ _22776_/X VGND VGND VPWR VPWR _22777_/Y sky130_fd_sc_hd__inv_2
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12334__A2_N _12332_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12530_ _24862_/Q VGND VGND VPWR VPWR _12530_/Y sky130_fd_sc_hd__inv_2
X_24516_ _24133_/CLK _24516_/D HRESETn VGND VGND VPWR VPWR _24516_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_38_0_HCLK clkbuf_5_19_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_77_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_21728_ _21721_/Y _21722_/Y _21725_/Y _21728_/D VGND VGND VPWR VPWR _21728_/X sky130_fd_sc_hd__or4_4
XFILLER_158_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25496_ _25499_/CLK _25496_/D HRESETn VGND VGND VPWR VPWR _11932_/B sky130_fd_sc_hd__dfrtp_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23022__A _24602_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12461_ _12461_/A VGND VGND VPWR VPWR _12461_/Y sky130_fd_sc_hd__inv_2
X_24447_ _24477_/CLK _16788_/X HRESETn VGND VGND VPWR VPWR _16786_/A sky130_fd_sc_hd__dfrtp_4
X_21659_ _21472_/A _21657_/X _21658_/X VGND VGND VPWR VPWR _21659_/X sky130_fd_sc_hd__and3_4
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14200_ _14198_/Y _14199_/X _13791_/X _14190_/X VGND VGND VPWR VPWR _25205_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18116__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17020__A _24645_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15180_ _15180_/A VGND VGND VPWR VPWR _15180_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12392_ _12391_/X VGND VGND VPWR VPWR _25461_/D sky130_fd_sc_hd__inv_2
X_24378_ _24725_/CLK _24378_/D HRESETn VGND VGND VPWR VPWR _16991_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_149_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14131_ _14091_/A _14091_/B _14091_/A _14091_/B VGND VGND VPWR VPWR _14131_/X sky130_fd_sc_hd__a2bb2o_4
X_23329_ _23329_/A _23022_/B VGND VGND VPWR VPWR _23329_/X sky130_fd_sc_hd__or2_4
XFILLER_125_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24333__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14062_ _14054_/A _14061_/Y VGND VGND VPWR VPWR _14062_/X sky130_fd_sc_hd__and2_4
XFILLER_153_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13013_ _12987_/X _13005_/D _13005_/A VGND VGND VPWR VPWR _13013_/X sky130_fd_sc_hd__o21a_4
X_18870_ _23950_/Q VGND VGND VPWR VPWR _18871_/A sky130_fd_sc_hd__inv_2
XFILLER_121_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17821_ _17761_/A _16921_/Y _17760_/Y _17813_/B VGND VGND VPWR VPWR _17827_/B sky130_fd_sc_hd__or4_4
XFILLER_0_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12611__B _12681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25539__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17752_ _17752_/A _16917_/Y _17752_/C VGND VGND VPWR VPWR _17753_/D sky130_fd_sc_hd__or3_4
XANTENNA__12477__B1 _12382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14964_ _14964_/A VGND VGND VPWR VPWR _14964_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16703_ _24484_/Q VGND VGND VPWR VPWR _16703_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13915_ _24974_/Q _13913_/X _13922_/A _13914_/X VGND VGND VPWR VPWR _13915_/X sky130_fd_sc_hd__or4_4
XANTENNA__17504__A1_N _25541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17683_ _17574_/D _17668_/B VGND VGND VPWR VPWR _17685_/B sky130_fd_sc_hd__nand2_4
XFILLER_74_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14895_ _24424_/Q VGND VGND VPWR VPWR _14895_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19422_ _19421_/Y _19419_/X _19351_/X _19419_/X VGND VGND VPWR VPWR _23743_/D sky130_fd_sc_hd__a2bb2o_4
X_16634_ _16634_/A VGND VGND VPWR VPWR _24512_/D sky130_fd_sc_hd__inv_2
XFILLER_35_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16130__A1_N _16128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13846_ _13844_/X _13845_/Y _20476_/B VGND VGND VPWR VPWR _13846_/X sky130_fd_sc_hd__a21o_4
XANTENNA__25121__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19353_ _18103_/B VGND VGND VPWR VPWR _19353_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21940__A _21463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13777_ _21138_/A _12081_/A _12084_/A _17436_/B VGND VGND VPWR VPWR _14462_/A sky130_fd_sc_hd__or4_4
X_16565_ _16564_/Y _16560_/X _16391_/X _16560_/X VGND VGND VPWR VPWR _24537_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_62_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18304_ _18301_/X _18306_/A _18298_/X VGND VGND VPWR VPWR _24214_/D sky130_fd_sc_hd__o21a_4
X_15516_ _11673_/B VGND VGND VPWR VPWR _15516_/Y sky130_fd_sc_hd__inv_2
X_12728_ _12728_/A VGND VGND VPWR VPWR _12728_/Y sky130_fd_sc_hd__inv_2
X_19284_ _19281_/Y _19276_/X _19282_/X _19283_/X VGND VGND VPWR VPWR _23792_/D sky130_fd_sc_hd__a2bb2o_4
X_16496_ _16521_/A VGND VGND VPWR VPWR _16496_/X sky130_fd_sc_hd__buf_2
XANTENNA__20556__A _14096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_230_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18235_ _18234_/Y VGND VGND VPWR VPWR _18236_/A sky130_fd_sc_hd__buf_2
XFILLER_176_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12659_ _12677_/A _12659_/B _12658_/X VGND VGND VPWR VPWR _25422_/D sky130_fd_sc_hd__and3_4
X_15447_ _15429_/A VGND VGND VPWR VPWR _15447_/X sky130_fd_sc_hd__buf_2
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18166_ _17966_/X _18165_/X _24244_/Q _18024_/X VGND VGND VPWR VPWR _24244_/D sky130_fd_sc_hd__o22a_4
X_15378_ _15300_/A _15376_/A VGND VGND VPWR VPWR _15378_/X sky130_fd_sc_hd__or2_4
XANTENNA__22771__A _24801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17117_ _17043_/B _17117_/B VGND VGND VPWR VPWR _17120_/B sky130_fd_sc_hd__or2_4
X_14329_ _14329_/A _14334_/A _14329_/C _14332_/B VGND VGND VPWR VPWR _14329_/X sky130_fd_sc_hd__or4_4
XFILLER_117_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18097_ _18097_/A _23823_/Q VGND VGND VPWR VPWR _18098_/C sky130_fd_sc_hd__or2_4
XFILLER_128_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24074__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_58_0_HCLK clkbuf_8_59_0_HCLK/A VGND VGND VPWR VPWR _25272_/CLK sky130_fd_sc_hd__clkbuf_1
X_17048_ _17019_/Y _17047_/X VGND VGND VPWR VPWR _17050_/B sky130_fd_sc_hd__nor2_4
XANTENNA__24003__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24958__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18999_ _18997_/Y _18993_/X _18998_/X _18986_/A VGND VGND VPWR VPWR _23891_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20961_ _25326_/Q _11929_/X _11948_/B VGND VGND VPWR VPWR _20961_/X sky130_fd_sc_hd__a21o_4
X_22700_ _22700_/A VGND VGND VPWR VPWR _22726_/B sky130_fd_sc_hd__inv_2
XFILLER_242_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23680_ _23559_/CLK _19608_/X VGND VGND VPWR VPWR _19605_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_81_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20892_ _20919_/A VGND VGND VPWR VPWR _20892_/X sky130_fd_sc_hd__buf_2
XFILLER_242_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22946__A _22946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22631_ _21109_/A _22630_/X _22296_/X _24867_/Q _21098_/A VGND VGND VPWR VPWR _22631_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_241_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25350_ _25346_/CLK _13055_/X HRESETn VGND VGND VPWR VPWR _25350_/Q sky130_fd_sc_hd__dfrtp_4
X_22562_ _22279_/A _22561_/X _21541_/X _24726_/Q _21708_/X VGND VGND VPWR VPWR _22562_/X
+ sky130_fd_sc_hd__a32o_4
X_24301_ _24297_/CLK _17676_/X HRESETn VGND VGND VPWR VPWR _24301_/Q sky130_fd_sc_hd__dfrtp_4
X_21513_ _18274_/A _21508_/X _21510_/X _21512_/X VGND VGND VPWR VPWR _21513_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24844__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25281_ _24227_/CLK _25281_/D HRESETn VGND VGND VPWR VPWR _11836_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_10_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22493_ _22194_/A VGND VGND VPWR VPWR _22493_/X sky130_fd_sc_hd__buf_2
XFILLER_166_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24232_ _24233_/CLK _18253_/X HRESETn VGND VGND VPWR VPWR _11808_/A sky130_fd_sc_hd__dfrtp_4
X_21444_ _21525_/A _21438_/X _23277_/A _21443_/X VGND VGND VPWR VPWR _21444_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__22455__A1 _16515_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14393__B1 _14392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18659__B1 _16569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22455__B2 _16792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15999__A1_N _15995_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24163_ _24654_/CLK _18584_/X HRESETn VGND VGND VPWR VPWR _24163_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17775__A _16913_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21375_ _19570_/X VGND VGND VPWR VPWR _21959_/B sky130_fd_sc_hd__buf_2
XANTENNA__17331__B1 _17276_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23114_ _23108_/X _23111_/Y _22868_/X _23113_/X VGND VGND VPWR VPWR _23115_/D sky130_fd_sc_hd__a2bb2o_4
X_20326_ _20326_/A VGND VGND VPWR VPWR _22343_/B sky130_fd_sc_hd__inv_2
X_24094_ _23916_/CLK _24094_/D HRESETn VGND VGND VPWR VPWR _11979_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_1_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20218__B1 _19759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15893__B1 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23045_ _24635_/Q _22904_/X VGND VGND VPWR VPWR _23045_/X sky130_fd_sc_hd__or2_4
XFILLER_150_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20257_ _20257_/A VGND VGND VPWR VPWR _21408_/B sky130_fd_sc_hd__inv_2
XFILLER_103_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14630__C _14630_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20188_ _20187_/Y _20185_/X _20099_/X _20185_/X VGND VGND VPWR VPWR _20188_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24996_ _25005_/CLK _24996_/D HRESETn VGND VGND VPWR VPWR _24996_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11961_ _11948_/A _11938_/A _11961_/C VGND VGND VPWR VPWR _11962_/B sky130_fd_sc_hd__or3_4
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23947_ _25134_/CLK _23947_/D HRESETn VGND VGND VPWR VPWR _23947_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_233_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13700_ _13664_/Y VGND VGND VPWR VPWR _13700_/X sky130_fd_sc_hd__buf_2
XFILLER_244_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14680_ _21252_/A VGND VGND VPWR VPWR _14681_/A sky130_fd_sc_hd__buf_2
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11892_ _11888_/X VGND VGND VPWR VPWR _11892_/Y sky130_fd_sc_hd__inv_2
X_23878_ _23844_/CLK _19038_/X VGND VGND VPWR VPWR _19037_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_189_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22856__A _22819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16070__B1 _15976_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13631_ _13631_/A VGND VGND VPWR VPWR _14294_/A sky130_fd_sc_hd__buf_2
X_22829_ _22829_/A VGND VGND VPWR VPWR _22829_/X sky130_fd_sc_hd__buf_2
XFILLER_232_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14620__B2 _14611_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13562_ _13562_/A VGND VGND VPWR VPWR _13562_/Y sky130_fd_sc_hd__inv_2
X_16350_ _16318_/A VGND VGND VPWR VPWR _16350_/X sky130_fd_sc_hd__buf_2
XANTENNA__18898__B1 _17440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25100__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12513_ _25411_/Q _12511_/Y _12512_/Y _24881_/Q VGND VGND VPWR VPWR _12513_/X sky130_fd_sc_hd__a2bb2o_4
X_15301_ _15301_/A _15331_/B VGND VGND VPWR VPWR _15301_/X sky130_fd_sc_hd__or2_4
X_16281_ _24642_/Q VGND VGND VPWR VPWR _16281_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24585__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13493_ _13492_/Y _13488_/X _11770_/X _13488_/X VGND VGND VPWR VPWR _25312_/D sky130_fd_sc_hd__a2bb2o_4
X_25479_ _25479_/CLK _25479_/D HRESETn VGND VGND VPWR VPWR _12078_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_157_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18020_ _18020_/A _18015_/X _18020_/C VGND VGND VPWR VPWR _18021_/C sky130_fd_sc_hd__or3_4
XFILLER_200_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12444_ _12434_/A _12444_/B _12444_/C VGND VGND VPWR VPWR _12444_/X sky130_fd_sc_hd__and3_4
X_15232_ _15231_/X VGND VGND VPWR VPWR _25022_/D sky130_fd_sc_hd__inv_2
XANTENNA__24514__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_211_0_HCLK clkbuf_8_211_0_HCLK/A VGND VGND VPWR VPWR _24427_/CLK sky130_fd_sc_hd__clkbuf_1
X_15163_ _14883_/A _15162_/Y VGND VGND VPWR VPWR _15163_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_3_0_0_HCLK_A clkbuf_3_1_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12375_ _12167_/A _12374_/Y VGND VGND VPWR VPWR _12377_/B sky130_fd_sc_hd__or2_4
XFILLER_176_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14114_ _14113_/X VGND VGND VPWR VPWR _14114_/X sky130_fd_sc_hd__buf_2
X_15094_ _24588_/Q VGND VGND VPWR VPWR _15094_/Y sky130_fd_sc_hd__inv_2
X_19971_ _19962_/Y VGND VGND VPWR VPWR _19971_/X sky130_fd_sc_hd__buf_2
XFILLER_4_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20209__B1 _19702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15884__B1 _22714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14045_ _14044_/X VGND VGND VPWR VPWR _14067_/A sky130_fd_sc_hd__buf_2
X_18922_ _13334_/B VGND VGND VPWR VPWR _18922_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12698__B1 _12641_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21957__B1 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18853_ _16487_/Y _24145_/Q _16487_/Y _24145_/Q VGND VGND VPWR VPWR _18853_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21935__A _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25373__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17804_ _17795_/X VGND VGND VPWR VPWR _17804_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18784_ _18686_/B VGND VGND VPWR VPWR _18788_/B sky130_fd_sc_hd__buf_2
XFILLER_94_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15996_ HWDATA[29] VGND VGND VPWR VPWR _15996_/X sky130_fd_sc_hd__buf_2
XANTENNA__21709__B1 _24719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_208_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17735_ _17731_/X _17734_/X _17731_/X _17734_/X VGND VGND VPWR VPWR _17735_/X sky130_fd_sc_hd__a2bb2o_4
X_14947_ _25021_/Q VGND VGND VPWR VPWR _15063_/A sky130_fd_sc_hd__inv_2
XFILLER_82_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17666_ _17578_/Y _17666_/B VGND VGND VPWR VPWR _17686_/A sky130_fd_sc_hd__or2_4
X_14878_ _14878_/A VGND VGND VPWR VPWR _14878_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22766__A _22733_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19405_ _19405_/A VGND VGND VPWR VPWR _19405_/Y sky130_fd_sc_hd__inv_2
X_16617_ _24516_/Q VGND VGND VPWR VPWR _16617_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13829_ _13829_/A VGND VGND VPWR VPWR _13829_/X sky130_fd_sc_hd__buf_2
X_17597_ _17597_/A _17597_/B VGND VGND VPWR VPWR _17600_/B sky130_fd_sc_hd__or2_4
XFILLER_211_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19336_ _23772_/Q VGND VGND VPWR VPWR _19336_/Y sky130_fd_sc_hd__inv_2
X_16548_ _16548_/A VGND VGND VPWR VPWR _16548_/X sky130_fd_sc_hd__buf_2
XFILLER_210_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22685__A1 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_21_0_HCLK clkbuf_5_10_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19267_ _21614_/B _19266_/X _16882_/X _19266_/X VGND VGND VPWR VPWR _23797_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16479_ _24569_/Q VGND VGND VPWR VPWR _16479_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18218_ _18014_/A _18218_/B VGND VGND VPWR VPWR _18218_/X sky130_fd_sc_hd__or2_4
XANTENNA__24255__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19198_ _18161_/B VGND VGND VPWR VPWR _19198_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12925__A1 _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18149_ _13617_/X _18141_/X _18148_/X VGND VGND VPWR VPWR _18149_/X sky130_fd_sc_hd__and3_4
XANTENNA__21829__B _21751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20999__A1 _14817_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23288__A1_N _12254_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21160_ _14203_/Y _14181_/A _21158_/Y _21159_/X VGND VGND VPWR VPWR _21162_/C sky130_fd_sc_hd__o22a_4
XFILLER_236_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12809__A2_N _24789_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20111_ _23499_/Q VGND VGND VPWR VPWR _20111_/Y sky130_fd_sc_hd__inv_2
X_21091_ _21090_/X VGND VGND VPWR VPWR _21091_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16004__A HWDATA[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20042_ _20041_/Y _20039_/X _19817_/X _20039_/X VGND VGND VPWR VPWR _20042_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24850_ _25390_/CLK _24850_/D HRESETn VGND VGND VPWR VPWR _24850_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25043__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23801_ _24413_/CLK _23801_/D VGND VGND VPWR VPWR _23801_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24781_ _24855_/CLK _15919_/X HRESETn VGND VGND VPWR VPWR _24781_/Q sky130_fd_sc_hd__dfrtp_4
X_21993_ _21993_/A _20324_/Y _21992_/X VGND VGND VPWR VPWR _21993_/X sky130_fd_sc_hd__and3_4
XFILLER_39_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23732_ _23747_/CLK _23732_/D VGND VGND VPWR VPWR _19449_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_227_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20944_ _13653_/X VGND VGND VPWR VPWR _20949_/B sky130_fd_sc_hd__inv_2
XPHY_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_103_0_HCLK clkbuf_6_51_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_206_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ _24209_/CLK _23663_/D VGND VGND VPWR VPWR _13303_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_42_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21566__A2_N _16180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14609__D _13525_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20875_ _20874_/X VGND VGND VPWR VPWR _20875_/X sky130_fd_sc_hd__buf_2
XFILLER_241_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22125__B1 _21556_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22614_ _22581_/X _22614_/B _22614_/C _22613_/Y VGND VGND VPWR VPWR HRDATA[11] sky130_fd_sc_hd__or4_4
X_25402_ _25403_/CLK _25402_/D HRESETn VGND VGND VPWR VPWR _12724_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23594_ _23575_/CLK _19858_/X VGND VGND VPWR VPWR _19854_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25333_ _23391_/CLK _25333_/D HRESETn VGND VGND VPWR VPWR _25333_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22545_ _17347_/C _22543_/X _22544_/Y VGND VGND VPWR VPWR _22545_/X sky130_fd_sc_hd__o21a_4
XFILLER_167_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25264_ _25089_/CLK _13821_/X HRESETn VGND VGND VPWR VPWR _13820_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_167_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22476_ _22476_/A _23278_/B VGND VGND VPWR VPWR _22476_/X sky130_fd_sc_hd__or2_4
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24215_ _23678_/CLK _24215_/D HRESETn VGND VGND VPWR VPWR _18314_/A sky130_fd_sc_hd__dfrtp_4
X_21427_ _21427_/A VGND VGND VPWR VPWR _21427_/X sky130_fd_sc_hd__buf_2
X_25195_ _25043_/CLK _14228_/X HRESETn VGND VGND VPWR VPWR _25195_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21739__B _21579_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12160_ _13462_/C _12058_/B _12160_/C _13483_/A VGND VGND VPWR VPWR _12160_/X sky130_fd_sc_hd__or4_4
X_24146_ _24146_/CLK _24146_/D HRESETn VGND VGND VPWR VPWR _24146_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21358_ _13501_/Y _21570_/A _12029_/Y _21571_/A VGND VGND VPWR VPWR _21358_/X sky130_fd_sc_hd__o22a_4
XFILLER_108_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21651__A2 _21648_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14945__A2_N _24428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23978__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15866__B1 _15564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_41_0_HCLK clkbuf_7_20_0_HCLK/X VGND VGND VPWR VPWR _25499_/CLK sky130_fd_sc_hd__clkbuf_1
X_20309_ _17446_/X _22396_/B VGND VGND VPWR VPWR _20309_/X sky130_fd_sc_hd__or2_4
X_12091_ _12080_/Y _12090_/X _11753_/X _12090_/X VGND VGND VPWR VPWR _25478_/D sky130_fd_sc_hd__a2bb2o_4
X_24077_ _24074_/CLK _24077_/D HRESETn VGND VGND VPWR VPWR _24077_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21289_ _21119_/X VGND VGND VPWR VPWR _21289_/X sky130_fd_sc_hd__buf_2
XFILLER_122_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23028_ _23094_/A _23027_/X VGND VGND VPWR VPWR _23028_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__17952__B _17952_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16849__A _19063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15850_ _15850_/A VGND VGND VPWR VPWR _15850_/X sky130_fd_sc_hd__buf_2
XFILLER_92_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14801_ _14814_/C _14799_/Y _14801_/C VGND VGND VPWR VPWR _14802_/C sky130_fd_sc_hd__and3_4
XFILLER_76_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15781_ _15781_/A VGND VGND VPWR VPWR _15918_/B sky130_fd_sc_hd__buf_2
XANTENNA__21167__A1 _16536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12993_ _12993_/A _12993_/B VGND VGND VPWR VPWR _12994_/C sky130_fd_sc_hd__or2_4
X_24979_ _24980_/CLK _24979_/D HRESETn VGND VGND VPWR VPWR _24979_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_206_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17520_ _25529_/Q _24300_/Q _11752_/Y _17519_/Y VGND VGND VPWR VPWR _17520_/X sky130_fd_sc_hd__o22a_4
X_14732_ _14728_/Y _14731_/Y _14727_/X _14730_/X VGND VGND VPWR VPWR _14732_/X sky130_fd_sc_hd__o22a_4
XFILLER_91_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11944_ _11944_/A VGND VGND VPWR VPWR _11944_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16043__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17451_ _13187_/A _17450_/X VGND VGND VPWR VPWR _17451_/X sky130_fd_sc_hd__and2_4
XFILLER_232_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24766__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11875_ _11801_/Y _11896_/B _11858_/Y _11874_/X VGND VGND VPWR VPWR _11875_/X sky130_fd_sc_hd__a211o_4
X_14663_ _25070_/Q VGND VGND VPWR VPWR _21787_/A sky130_fd_sc_hd__inv_2
XFILLER_233_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16402_ HWDATA[17] VGND VGND VPWR VPWR _16402_/X sky130_fd_sc_hd__buf_2
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13614_ _13614_/A _14787_/A _13610_/Y _13614_/D VGND VGND VPWR VPWR _13620_/C sky130_fd_sc_hd__or4_4
XFILLER_232_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17382_ _17341_/A _17344_/B _17381_/X VGND VGND VPWR VPWR _24341_/D sky130_fd_sc_hd__and3_4
X_14594_ _14553_/B _14593_/Y _14588_/X _14591_/X _13569_/A VGND VGND VPWR VPWR _25087_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_220_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19121_ _18012_/B VGND VGND VPWR VPWR _19121_/Y sky130_fd_sc_hd__inv_2
X_16333_ _16331_/Y _16332_/X _16240_/X _16332_/X VGND VGND VPWR VPWR _24623_/D sky130_fd_sc_hd__a2bb2o_4
X_13545_ _13544_/Y _14548_/A _13544_/Y _14548_/A VGND VGND VPWR VPWR _13545_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12617__A _12681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19052_ _19051_/Y _19049_/X _18981_/X _19049_/X VGND VGND VPWR VPWR _23873_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13476_ _13464_/A VGND VGND VPWR VPWR _13476_/X sky130_fd_sc_hd__buf_2
X_16264_ _16263_/Y _16184_/X _15901_/X _16184_/X VGND VGND VPWR VPWR _16264_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14440__A1_N _14171_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18003_ _18085_/A _18000_/X _18003_/C VGND VGND VPWR VPWR _18009_/B sky130_fd_sc_hd__and3_4
X_12427_ _12426_/X VGND VGND VPWR VPWR _25453_/D sky130_fd_sc_hd__inv_2
X_15215_ _14921_/X _15214_/X _15169_/X VGND VGND VPWR VPWR _15215_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__19296__B1 _19295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16195_ _23206_/A VGND VGND VPWR VPWR _16195_/Y sky130_fd_sc_hd__inv_2
X_12358_ _25357_/Q _12356_/Y _12357_/Y _24840_/Q VGND VGND VPWR VPWR _12358_/X sky130_fd_sc_hd__a2bb2o_4
X_15146_ _24998_/Q _15144_/Y _15293_/B _24600_/Q VGND VGND VPWR VPWR _15147_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15077_ _15077_/A _15077_/B _15074_/X _15077_/D VGND VGND VPWR VPWR _15116_/A sky130_fd_sc_hd__or4_4
X_19954_ _19952_/Y _19953_/X _19617_/X _19953_/X VGND VGND VPWR VPWR _23557_/D sky130_fd_sc_hd__a2bb2o_4
X_12289_ _12281_/X _12283_/X _12289_/C _12288_/X VGND VGND VPWR VPWR _12289_/X sky130_fd_sc_hd__or4_4
XFILLER_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14028_ _14028_/A _14028_/B VGND VGND VPWR VPWR _14029_/B sky130_fd_sc_hd__nand2_4
X_18905_ _11699_/A _11707_/X HWDATA[30] _24113_/Q _11708_/X VGND VGND VPWR VPWR _24113_/D
+ sky130_fd_sc_hd__a32o_4
X_19885_ _19883_/Y _19879_/X _19606_/X _19884_/X VGND VGND VPWR VPWR _23584_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15609__B1 _13818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16759__A _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18836_ _16494_/A _24142_/Q _16494_/Y _18692_/Y VGND VGND VPWR VPWR _18836_/X sky130_fd_sc_hd__o22a_4
XFILLER_110_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18271__A1 _13783_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16282__B1 _15554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18767_ _18691_/B _18767_/B VGND VGND VPWR VPWR _18770_/B sky130_fd_sc_hd__or2_4
XFILLER_209_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15979_ _15784_/X _15850_/A _15920_/X _21088_/A _15925_/X VGND VGND VPWR VPWR _24748_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17718_ _21208_/A VGND VGND VPWR VPWR _21924_/A sky130_fd_sc_hd__buf_2
X_18698_ _18698_/A _18697_/X VGND VGND VPWR VPWR _18706_/A sky130_fd_sc_hd__or2_4
XANTENNA__16034__B1 _11726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17649_ _17647_/A _17643_/B _17648_/Y VGND VGND VPWR VPWR _17649_/X sky130_fd_sc_hd__and3_4
XANTENNA__16494__A _16494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24436__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20660_ _17394_/A _17394_/B VGND VGND VPWR VPWR _20660_/Y sky130_fd_sc_hd__nand2_4
XFILLER_195_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19319_ _23778_/Q VGND VGND VPWR VPWR _19319_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20591_ _20591_/A VGND VGND VPWR VPWR _23947_/D sky130_fd_sc_hd__inv_2
X_22330_ _20628_/A _21722_/B _20673_/A _22181_/B VGND VGND VPWR VPWR _22330_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23120__A _22468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22261_ _22261_/A _19859_/Y VGND VGND VPWR VPWR _22263_/B sky130_fd_sc_hd__or2_4
XFILLER_118_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15838__A _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23083__A1 _12194_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13020__B1 _13019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24000_ _25226_/CLK _20523_/X HRESETn VGND VGND VPWR VPWR _20522_/A sky130_fd_sc_hd__dfrtp_4
X_21212_ _18314_/Y _21203_/X _21212_/C VGND VGND VPWR VPWR _21212_/X sky130_fd_sc_hd__or3_4
XFILLER_133_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22192_ _21124_/B _22191_/X _21298_/X VGND VGND VPWR VPWR _22192_/X sky130_fd_sc_hd__and3_4
XANTENNA__22830__B2 _22290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_0_0_HCLK clkbuf_7_0_0_HCLK/X VGND VGND VPWR VPWR _23378_/CLK sky130_fd_sc_hd__clkbuf_1
X_21143_ _18896_/Y _21132_/Y _21343_/A _21142_/X VGND VGND VPWR VPWR _21224_/A sky130_fd_sc_hd__a211o_4
Xclkbuf_7_28_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_28_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21074_ _21056_/X _21059_/X _21073_/X VGND VGND VPWR VPWR _21074_/X sky130_fd_sc_hd__and3_4
XFILLER_113_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20025_ _20012_/Y VGND VGND VPWR VPWR _20025_/X sky130_fd_sc_hd__buf_2
X_24902_ _24903_/CLK _15611_/X HRESETn VGND VGND VPWR VPWR _24902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24833_ _24855_/CLK _15816_/X HRESETn VGND VGND VPWR VPWR _24833_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21149__A1 _13503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _21278_/X _21974_/X _21975_/X _23346_/A _21643_/X VGND VGND VPWR VPWR _21977_/B
+ sky130_fd_sc_hd__a32o_4
X_24764_ _25375_/CLK _24764_/D HRESETn VGND VGND VPWR VPWR _24764_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20927_ _20919_/X _20926_/Y _24501_/Q _20923_/X VGND VGND VPWR VPWR _24057_/D sky130_fd_sc_hd__a2bb2o_4
X_23715_ _23691_/CLK _23715_/D VGND VGND VPWR VPWR _23715_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24695_ _24696_/CLK _16130_/X HRESETn VGND VGND VPWR VPWR _24695_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14917__A _14917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24177__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11660_/A VGND VGND VPWR VPWR _14365_/C sky130_fd_sc_hd__buf_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _20862_/A _20862_/B _20857_/X VGND VGND VPWR VPWR _20858_/X sky130_fd_sc_hd__o21a_4
X_23646_ _23665_/CLK _23646_/D VGND VGND VPWR VPWR _13346_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_187_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24106__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23577_ _24199_/CLK _19903_/X VGND VGND VPWR VPWR _19902_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20789_ _20789_/A VGND VGND VPWR VPWR _20789_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21321__A1 _21289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _13394_/A _13330_/B _13329_/X VGND VGND VPWR VPWR _13338_/B sky130_fd_sc_hd__or3_4
XFILLER_167_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22528_ _22528_/A _22528_/B _22521_/Y _22528_/D VGND VGND VPWR VPWR _22528_/X sky130_fd_sc_hd__or4_4
X_25316_ _25474_/CLK _13486_/X HRESETn VGND VGND VPWR VPWR _12009_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13300_/A _13259_/X _13260_/X VGND VGND VPWR VPWR _13261_/X sky130_fd_sc_hd__and3_4
XANTENNA__15748__A HWDATA[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22459_ _16272_/X _22459_/B VGND VGND VPWR VPWR _22472_/A sky130_fd_sc_hd__nor2_4
X_25247_ _25249_/CLK _13866_/X HRESETn VGND VGND VPWR VPWR _21723_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14884__A2_N _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12212_ _21534_/A VGND VGND VPWR VPWR _12212_/Y sky130_fd_sc_hd__inv_2
X_15000_ _24475_/Q VGND VGND VPWR VPWR _15000_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13192_ _13396_/A _23857_/Q VGND VGND VPWR VPWR _13193_/C sky130_fd_sc_hd__or2_4
X_25178_ _23887_/CLK _25178_/D HRESETn VGND VGND VPWR VPWR MSO_S2 sky130_fd_sc_hd__dfrtp_4
XFILLER_157_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12143_ _12139_/A _12135_/X _12141_/Y VGND VGND VPWR VPWR _12143_/X sky130_fd_sc_hd__o21a_4
X_24129_ _24133_/CLK _24129_/D HRESETn VGND VGND VPWR VPWR _18683_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13268__A _13397_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20832__B1 _20828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12074_ _12074_/A VGND VGND VPWR VPWR _12074_/Y sky130_fd_sc_hd__inv_2
X_16951_ _16950_/X VGND VGND VPWR VPWR _17791_/A sky130_fd_sc_hd__inv_2
XFILLER_104_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22585__B1 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15902_ _12783_/Y _15896_/X _15901_/X _15861_/X VGND VGND VPWR VPWR _15902_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_238_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19670_ _13141_/B VGND VGND VPWR VPWR _19670_/Y sky130_fd_sc_hd__inv_2
X_16882_ _19824_/A VGND VGND VPWR VPWR _16882_/X sky130_fd_sc_hd__buf_2
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12900__A _12838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19450__B1 _19360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16264__B1 _15901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18621_ _24134_/Q VGND VGND VPWR VPWR _18783_/A sky130_fd_sc_hd__inv_2
X_15833_ _12322_/Y _15827_/X _15472_/X _15827_/X VGND VGND VPWR VPWR _24822_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24947__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18552_ _16441_/X _18478_/X VGND VGND VPWR VPWR _18553_/B sky130_fd_sc_hd__or2_4
X_15764_ _11780_/A VGND VGND VPWR VPWR _15764_/X sky130_fd_sc_hd__buf_2
X_12976_ _12302_/Y _12291_/X _12976_/C _12976_/D VGND VGND VPWR VPWR _12976_/X sky130_fd_sc_hd__or4_4
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17503_ _24110_/Q VGND VGND VPWR VPWR _17503_/Y sky130_fd_sc_hd__inv_2
X_14715_ _14715_/A VGND VGND VPWR VPWR _14715_/Y sky130_fd_sc_hd__inv_2
X_11927_ _19620_/A VGND VGND VPWR VPWR _11927_/X sky130_fd_sc_hd__buf_2
X_18483_ _16441_/X _18416_/Y _18493_/A _18483_/D VGND VGND VPWR VPWR _18483_/X sky130_fd_sc_hd__or4_4
XFILLER_205_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15695_ _24887_/Q _15694_/X _15687_/A VGND VGND VPWR VPWR _24887_/D sky130_fd_sc_hd__o21a_4
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17434_ _17433_/Y _17429_/X _16716_/X _17429_/A VGND VGND VPWR VPWR _17434_/X sky130_fd_sc_hd__a2bb2o_4
X_14646_ _19387_/A VGND VGND VPWR VPWR _19341_/A sky130_fd_sc_hd__buf_2
X_11858_ _11857_/X VGND VGND VPWR VPWR _11858_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17365_ _17346_/A _17367_/B _17364_/Y VGND VGND VPWR VPWR _17365_/X sky130_fd_sc_hd__o21a_4
X_11789_ _11699_/X _11707_/X _11788_/X _25521_/Q _11708_/X VGND VGND VPWR VPWR _25521_/D
+ sky130_fd_sc_hd__a32o_4
X_14577_ _14562_/A _14575_/X _14576_/X _13758_/X _25094_/Q VGND VGND VPWR VPWR _14577_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15790__A2 _15789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19104_ _19103_/Y _19101_/X _19057_/X _19101_/X VGND VGND VPWR VPWR _23855_/D sky130_fd_sc_hd__a2bb2o_4
X_16316_ _16315_/Y _16311_/X _15953_/X _16311_/X VGND VGND VPWR VPWR _16316_/X sky130_fd_sc_hd__a2bb2o_4
X_13528_ _24251_/Q _24250_/Q _13528_/C VGND VGND VPWR VPWR _13528_/X sky130_fd_sc_hd__and3_4
XFILLER_186_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17296_ _17295_/X VGND VGND VPWR VPWR _24365_/D sky130_fd_sc_hd__inv_2
XFILLER_9_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19035_ _23879_/Q VGND VGND VPWR VPWR _19035_/Y sky130_fd_sc_hd__inv_2
X_16247_ _24655_/Q VGND VGND VPWR VPWR _16247_/Y sky130_fd_sc_hd__inv_2
X_13459_ _13459_/A VGND VGND VPWR VPWR _13459_/X sky130_fd_sc_hd__buf_2
X_16178_ _16364_/A _14178_/B _15636_/C _14365_/D VGND VGND VPWR VPWR _16179_/A sky130_fd_sc_hd__or4_4
XFILLER_126_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15129_ _15300_/A _24593_/Q _15300_/A _24593_/Q VGND VGND VPWR VPWR _15129_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19937_ _21209_/B _19932_/X _19874_/X _19932_/A VGND VGND VPWR VPWR _23563_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19868_ _19868_/A VGND VGND VPWR VPWR _19868_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19441__B1 _19395_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16255__B1 _16062_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20051__B2 _20034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24688__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18819_ _18819_/A _18815_/X VGND VGND VPWR VPWR _18819_/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19799_ _19798_/Y _19796_/X _19711_/X _19796_/X VGND VGND VPWR VPWR _19799_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21830_ _24039_/Q VGND VGND VPWR VPWR _21830_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24617__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21761_ _21757_/A _21759_/X _21761_/C VGND VGND VPWR VPWR _21761_/X sky130_fd_sc_hd__and3_4
XFILLER_212_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12292__B2 _24836_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20712_ _20712_/A VGND VGND VPWR VPWR _20712_/Y sky130_fd_sc_hd__inv_2
X_23500_ _23378_/CLK _23500_/D VGND VGND VPWR VPWR _23500_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24270__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24480_ _24035_/CLK _24480_/D HRESETn VGND VGND VPWR VPWR _24480_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_212_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21692_ _21503_/X _21691_/X _11841_/Y _21503_/X VGND VGND VPWR VPWR _21692_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_212_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23431_ _23441_/CLK _23431_/D VGND VGND VPWR VPWR _23431_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20643_ _20643_/A _20640_/A VGND VGND VPWR VPWR _20643_/Y sky130_fd_sc_hd__nand2_4
XFILLER_177_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18648__A1_N _16587_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12257__A _25439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22673__B _22816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22500__B1 _16915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23362_ _23349_/X VGND VGND VPWR VPWR IRQ[18] sky130_fd_sc_hd__buf_2
X_20574_ _14419_/Y _20566_/X _20557_/X _20573_/X VGND VGND VPWR VPWR _20575_/A sky130_fd_sc_hd__a211o_4
XFILLER_177_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22313_ _14421_/Y _22327_/B VGND VGND VPWR VPWR _22313_/Y sky130_fd_sc_hd__nor2_4
X_25101_ _25238_/CLK _25101_/D HRESETn VGND VGND VPWR VPWR scl_oen_o_S4 sky130_fd_sc_hd__dfstp_4
XANTENNA__25476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23293_ _23120_/X _23291_/X _23123_/X _23292_/X VGND VGND VPWR VPWR _23294_/B sky130_fd_sc_hd__o22a_4
X_25032_ _25021_/CLK _25032_/D HRESETn VGND VGND VPWR VPWR _14913_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22244_ _22015_/A _22244_/B VGND VGND VPWR VPWR _22244_/X sky130_fd_sc_hd__or2_4
XFILLER_3_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22173__A2_N _14245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22175_ _17366_/A _22429_/A _25439_/Q _21075_/Y VGND VGND VPWR VPWR _22175_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21126_ _21041_/X _21125_/X _13129_/Y _15661_/A VGND VGND VPWR VPWR _21126_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21057_ _21024_/X VGND VGND VPWR VPWR _21111_/A sky130_fd_sc_hd__buf_2
XFILLER_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23009__B _23075_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_115_0_HCLK clkbuf_7_57_0_HCLK/X VGND VGND VPWR VPWR _24886_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__16246__B1 _16141_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20008_ _19874_/A VGND VGND VPWR VPWR _20008_/X sky130_fd_sc_hd__buf_2
XFILLER_219_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16926__A2_N _17880_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_178_0_HCLK clkbuf_7_89_0_HCLK/X VGND VGND VPWR VPWR _23938_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_246_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12830_ _12830_/A _12781_/Y _12830_/C _12749_/Y VGND VGND VPWR VPWR _12835_/C sky130_fd_sc_hd__or4_4
X_24816_ _24886_/CLK _15858_/X HRESETn VGND VGND VPWR VPWR _24816_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24358__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12761_ _25392_/Q _24809_/Q _12759_/Y _12760_/Y VGND VGND VPWR VPWR _12761_/X sky130_fd_sc_hd__o22a_4
X_24747_ _24639_/CLK _24747_/D HRESETn VGND VGND VPWR VPWR _15980_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _19583_/Y _21959_/B VGND VGND VPWR VPWR _21959_/X sky130_fd_sc_hd__or2_4
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14499_/X VGND VGND VPWR VPWR _14500_/X sky130_fd_sc_hd__buf_2
XFILLER_243_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11712_ _11710_/Y _11692_/X _11711_/X _11692_/X VGND VGND VPWR VPWR _25540_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12692_/A _12711_/A VGND VGND VPWR VPWR _12692_/X sky130_fd_sc_hd__or2_4
X_15480_ HTRANS[1] VGND VGND VPWR VPWR _15480_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24678_ _24678_/CLK _16186_/X HRESETn VGND VGND VPWR VPWR _23329_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14366__B _21343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14431_/A VGND VGND VPWR VPWR _14431_/X sky130_fd_sc_hd__buf_2
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23629_ _23627_/CLK _23629_/D VGND VGND VPWR VPWR _19753_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12167__A _12167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _17149_/X VGND VGND VPWR VPWR _24377_/D sky130_fd_sc_hd__inv_2
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14362_ _20469_/A VGND VGND VPWR VPWR _14362_/Y sky130_fd_sc_hd__inv_2
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16101_ _23112_/A VGND VGND VPWR VPWR _16101_/Y sky130_fd_sc_hd__inv_2
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _13231_/X _13311_/X _13312_/X VGND VGND VPWR VPWR _13313_/X sky130_fd_sc_hd__and3_4
XFILLER_128_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14293_ _14293_/A VGND VGND VPWR VPWR _25179_/D sky130_fd_sc_hd__inv_2
X_17081_ _17074_/X VGND VGND VPWR VPWR _17085_/B sky130_fd_sc_hd__inv_2
XFILLER_7_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13244_ _11951_/X _13217_/X _13242_/X _25333_/Q _13243_/X VGND VGND VPWR VPWR _13244_/X
+ sky130_fd_sc_hd__o32a_4
X_16032_ _15988_/X VGND VGND VPWR VPWR _16038_/A sky130_fd_sc_hd__buf_2
XFILLER_164_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_14_0_HCLK_A clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13175_ _13175_/A _23914_/Q VGND VGND VPWR VPWR _13176_/C sky130_fd_sc_hd__or2_4
XFILLER_184_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22270__A2 _22250_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12126_ _24103_/Q _12120_/A _12125_/Y VGND VGND VPWR VPWR _12126_/X sky130_fd_sc_hd__o21a_4
X_17983_ _17983_/A VGND VGND VPWR VPWR _18227_/A sky130_fd_sc_hd__buf_2
XFILLER_112_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_11_0_HCLK clkbuf_6_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_22_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19722_ _13275_/B VGND VGND VPWR VPWR _19722_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_74_0_HCLK clkbuf_7_75_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_74_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12057_ _12057_/A VGND VGND VPWR VPWR _12057_/X sky130_fd_sc_hd__buf_2
X_16934_ _16930_/X _16934_/B _16934_/C _16934_/D VGND VGND VPWR VPWR _16934_/X sky130_fd_sc_hd__or4_4
XANTENNA__13726__A _13726_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12630__A _12681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16237__B1 _16236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21230__B1 _20822_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19653_ _19648_/Y _19651_/X _19652_/X _19651_/X VGND VGND VPWR VPWR _19653_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24781__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16865_ _14777_/X VGND VGND VPWR VPWR _16865_/X sky130_fd_sc_hd__buf_2
X_18604_ _16605_/A _18686_/B _16552_/Y _24153_/Q VGND VGND VPWR VPWR _18607_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23974__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15816_ _15810_/X _15813_/X _16233_/A _24833_/Q _15811_/X VGND VGND VPWR VPWR _15816_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24099__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24710__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19584_ _19583_/Y _19581_/X _19534_/X _19581_/X VGND VGND VPWR VPWR _23687_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_225_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16796_ _16796_/A VGND VGND VPWR VPWR _16796_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18535_ _18467_/A _18467_/B _18466_/B _18538_/B VGND VGND VPWR VPWR _18541_/B sky130_fd_sc_hd__or4_4
XANTENNA__24028__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15747_ _15745_/X _15738_/X _15746_/X _24867_/Q _15736_/X VGND VGND VPWR VPWR _15747_/X
+ sky130_fd_sc_hd__a32o_4
X_12959_ _12775_/Y _12959_/B VGND VGND VPWR VPWR _12963_/B sky130_fd_sc_hd__or2_4
XFILLER_61_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18466_ _18407_/Y _18466_/B _18466_/C _18465_/Y VGND VGND VPWR VPWR _18466_/X sky130_fd_sc_hd__or4_4
XFILLER_178_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15678_ _15676_/Y _15686_/A _15675_/Y VGND VGND VPWR VPWR _15678_/X sky130_fd_sc_hd__or3_4
XFILLER_233_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22774__A _22429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17417_ _24332_/Q VGND VGND VPWR VPWR _17417_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14629_ _18044_/A VGND VGND VPWR VPWR _18009_/A sky130_fd_sc_hd__buf_2
XFILLER_60_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18397_ _16200_/Y _18461_/A _16200_/Y _18461_/A VGND VGND VPWR VPWR _18397_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16772__A _24453_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17348_ _17348_/A VGND VGND VPWR VPWR _17349_/B sky130_fd_sc_hd__inv_2
XFILLER_158_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17279_ _17333_/A _17256_/B VGND VGND VPWR VPWR _17280_/A sky130_fd_sc_hd__or2_4
XFILLER_134_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19018_ _19011_/A VGND VGND VPWR VPWR _19018_/X sky130_fd_sc_hd__buf_2
X_20290_ _20290_/A VGND VGND VPWR VPWR _22244_/B sky130_fd_sc_hd__inv_2
XFILLER_173_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18699__A _18745_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22940__C _23075_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19662__B1 _19587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16476__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24869__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23980_ _23986_/CLK _23980_/D HRESETn VGND VGND VPWR VPWR _23980_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12540__A _24857_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22931_ _16444_/X _22927_/X _22930_/X VGND VGND VPWR VPWR _22931_/X sky130_fd_sc_hd__and3_4
XFILLER_217_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15851__A _15845_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24451__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22862_ _21424_/X _22861_/X _21427_/X _24873_/Q _21428_/X VGND VGND VPWR VPWR _22863_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24601_ _24597_/CLK _24601_/D HRESETn VGND VGND VPWR VPWR _15084_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_71_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21813_ _21809_/A _21813_/B VGND VGND VPWR VPWR _21813_/X sky130_fd_sc_hd__or2_4
X_22793_ _23060_/A _22793_/B VGND VGND VPWR VPWR _22793_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__21524__B2 _22522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21744_ _21738_/X _21744_/B VGND VGND VPWR VPWR _21751_/C sky130_fd_sc_hd__nor2_4
X_24532_ _24573_/CLK _16577_/X HRESETn VGND VGND VPWR VPWR _16576_/A sky130_fd_sc_hd__dfrtp_4
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21675_ _21674_/X VGND VGND VPWR VPWR _22021_/A sky130_fd_sc_hd__buf_2
X_24463_ _24463_/CLK _24463_/D HRESETn VGND VGND VPWR VPWR _15025_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20626_ _15465_/Y _20615_/X _20672_/A _20625_/X VGND VGND VPWR VPWR _20627_/A sky130_fd_sc_hd__a211o_4
X_23414_ _23415_/CLK _20337_/X VGND VGND VPWR VPWR _23414_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24394_ _24390_/CLK _24394_/D HRESETn VGND VGND VPWR VPWR _16964_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11776__B1 _11775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23345_ _18268_/Y _21822_/A _17478_/Y _21504_/A VGND VGND VPWR VPWR _23345_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20557_ _20556_/X VGND VGND VPWR VPWR _20557_/X sky130_fd_sc_hd__buf_2
XANTENNA__23029__B2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23011__C _23010_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23276_ _22129_/X _23275_/X _23145_/X _24850_/Q _22838_/X VGND VGND VPWR VPWR _23277_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_153_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20488_ _24076_/Q _20488_/B VGND VGND VPWR VPWR _20503_/C sky130_fd_sc_hd__and2_4
XFILLER_138_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22227_ _22212_/A _22227_/B _22227_/C VGND VGND VPWR VPWR _22228_/C sky130_fd_sc_hd__or3_4
X_25015_ _25015_/CLK _25015_/D HRESETn VGND VGND VPWR VPWR _25015_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20263__A1 _23442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22158_ _22041_/X _22127_/X _22158_/C _22158_/D VGND VGND VPWR VPWR HRDATA[5] sky130_fd_sc_hd__or4_4
XFILLER_160_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21109_ _21109_/A _21102_/X _21109_/C VGND VGND VPWR VPWR _21109_/X sky130_fd_sc_hd__and3_4
XFILLER_248_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24539__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14980_ _14935_/X _14979_/X VGND VGND VPWR VPWR _14981_/A sky130_fd_sc_hd__or2_4
X_22089_ _14710_/A _22065_/Y _22074_/Y _22082_/Y _22088_/Y VGND VGND VPWR VPWR _22089_/X
+ sky130_fd_sc_hd__a32o_4
X_13931_ _13931_/A _13931_/B _13915_/X _13947_/C VGND VGND VPWR VPWR _13940_/A sky130_fd_sc_hd__or4_4
XFILLER_75_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24192__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16650_ _24506_/Q VGND VGND VPWR VPWR _16650_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13862_ _13860_/X _13861_/X _14251_/A _13856_/X VGND VGND VPWR VPWR _13862_/X sky130_fd_sc_hd__o22a_4
XFILLER_19_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12579__A2_N _24858_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15601_ _15576_/A VGND VGND VPWR VPWR _15601_/X sky130_fd_sc_hd__buf_2
X_12813_ _25388_/Q VGND VGND VPWR VPWR _12813_/Y sky130_fd_sc_hd__inv_2
X_16581_ _16578_/Y _16580_/X _16320_/X _16580_/X VGND VGND VPWR VPWR _24531_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_216_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13793_ _13790_/Y _13784_/X _13791_/X _13792_/X VGND VGND VPWR VPWR _25273_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12256__B2 _24752_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18320_ _18320_/A _17736_/B _18317_/X _18319_/X VGND VGND VPWR VPWR _18320_/X sky130_fd_sc_hd__or4_4
X_15532_ _12086_/X _15530_/X HADDR[3] _15530_/X VGND VGND VPWR VPWR _15532_/X sky130_fd_sc_hd__a2bb2o_4
X_12744_ _25394_/Q VGND VGND VPWR VPWR _12744_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17195__B2 _17358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22594__A _24796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25398__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18251_ _18238_/X _18240_/X _18250_/X _24233_/Q _18241_/X VGND VGND VPWR VPWR _18251_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15463_ _15458_/A VGND VGND VPWR VPWR _15463_/X sky130_fd_sc_hd__buf_2
X_12675_ _12675_/A VGND VGND VPWR VPWR _12675_/Y sky130_fd_sc_hd__inv_2
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _17202_/A VGND VGND VPWR VPWR _17203_/A sky130_fd_sc_hd__inv_2
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25327__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14414_ _14414_/A VGND VGND VPWR VPWR _14414_/Y sky130_fd_sc_hd__inv_2
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18182_ _18182_/A _19020_/A VGND VGND VPWR VPWR _18184_/B sky130_fd_sc_hd__or2_4
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ _15379_/A _15394_/B _15393_/Y VGND VGND VPWR VPWR _15394_/X sky130_fd_sc_hd__and3_4
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11767__B1 _11765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _17038_/C _17132_/X _17053_/X VGND VGND VPWR VPWR _17133_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_128_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ _14345_/A VGND VGND VPWR VPWR _14345_/X sky130_fd_sc_hd__buf_2
XFILLER_128_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19892__B1 _19617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17064_ _17381_/B VGND VGND VPWR VPWR _17064_/X sky130_fd_sc_hd__buf_2
X_14276_ _25181_/Q VGND VGND VPWR VPWR _14280_/A sky130_fd_sc_hd__inv_2
XFILLER_183_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16015_ _16014_/Y _16012_/X _11691_/X _16012_/X VGND VGND VPWR VPWR _16015_/X sky130_fd_sc_hd__a2bb2o_4
X_13227_ _13421_/A VGND VGND VPWR VPWR _13227_/X sky130_fd_sc_hd__buf_2
XFILLER_171_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19644__B1 _19543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17854__C _16895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24962__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13158_ _13157_/X _23634_/Q VGND VGND VPWR VPWR _13158_/X sky130_fd_sc_hd__or2_4
XFILLER_98_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12109_ _12109_/A VGND VGND VPWR VPWR _12154_/A sky130_fd_sc_hd__inv_2
XFILLER_100_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13089_ _13089_/A VGND VGND VPWR VPWR _13090_/B sky130_fd_sc_hd__inv_2
X_17966_ _17966_/A VGND VGND VPWR VPWR _17966_/X sky130_fd_sc_hd__buf_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16917_ _16917_/A VGND VGND VPWR VPWR _16917_/Y sky130_fd_sc_hd__inv_2
X_19705_ _19704_/Y _19699_/X _19587_/X _19699_/X VGND VGND VPWR VPWR _23646_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24209__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17897_ _17896_/Y _17906_/B _21991_/A _17894_/Y VGND VGND VPWR VPWR _17910_/B sky130_fd_sc_hd__o22a_4
XFILLER_66_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16848_ _16847_/Y _16845_/X _16783_/X _16845_/X VGND VGND VPWR VPWR _16848_/X sky130_fd_sc_hd__a2bb2o_4
X_19636_ _13307_/B VGND VGND VPWR VPWR _19636_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_161_0_HCLK clkbuf_7_80_0_HCLK/X VGND VGND VPWR VPWR _25073_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_4_0_HCLK clkbuf_7_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19567_ _21192_/B _19562_/X _19475_/X _19549_/Y VGND VGND VPWR VPWR _23691_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_18_0_HCLK clkbuf_7_9_0_HCLK/X VGND VGND VPWR VPWR _23534_/CLK sky130_fd_sc_hd__clkbuf_1
X_16779_ _16725_/A VGND VGND VPWR VPWR _16779_/X sky130_fd_sc_hd__buf_2
XFILLER_240_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18518_ _24181_/Q _18521_/B VGND VGND VPWR VPWR _18518_/X sky130_fd_sc_hd__or2_4
X_19498_ _23715_/Q VGND VGND VPWR VPWR _21197_/B sky130_fd_sc_hd__inv_2
XFILLER_221_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18449_ _23238_/A _18440_/Y _16256_/Y _24162_/Q VGND VGND VPWR VPWR _18449_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25068__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21460_ _21803_/A _21457_/X _21459_/X VGND VGND VPWR VPWR _21460_/X sky130_fd_sc_hd__and3_4
XFILLER_178_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11758__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20411_ _20407_/Y _20410_/X _16854_/X _20410_/X VGND VGND VPWR VPWR _20411_/X sky130_fd_sc_hd__a2bb2o_4
X_21391_ _21387_/X _21390_/X _21247_/X VGND VGND VPWR VPWR _21391_/X sky130_fd_sc_hd__o21a_4
XFILLER_174_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23130_ _20796_/Y _22992_/X _20935_/Y _22794_/X VGND VGND VPWR VPWR _23131_/B sky130_fd_sc_hd__o22a_4
X_20342_ _20340_/Y _20341_/X _19617_/A _20341_/X VGND VGND VPWR VPWR _20342_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23061_ _20789_/Y _22992_/X _20928_/Y _21227_/X VGND VGND VPWR VPWR _23061_/X sky130_fd_sc_hd__o22a_4
X_20273_ _20271_/Y _20267_/X _19970_/X _20272_/X VGND VGND VPWR VPWR _20273_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16958__A1_N _24722_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22012_ _22020_/A _20271_/Y VGND VGND VPWR VPWR _22012_/X sky130_fd_sc_hd__or2_4
XANTENNA__16449__B1 _16361_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24632__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23963_ _23972_/CLK _25184_/Q HRESETn VGND VGND VPWR VPWR _22331_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_245_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15581__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22914_ _22194_/A VGND VGND VPWR VPWR _22914_/X sky130_fd_sc_hd__buf_2
X_23894_ _23844_/CLK _23894_/D VGND VGND VPWR VPWR _18122_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_72_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16621__B1 _13577_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22845_ _22824_/X _22828_/Y _22835_/Y _22844_/X VGND VGND VPWR VPWR _22845_/X sky130_fd_sc_hd__a211o_4
XANTENNA__12238__B2 _24763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22776_ _22486_/X _22775_/X _22489_/X _16031_/A _22490_/X VGND VGND VPWR VPWR _22776_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17177__B2 _17239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25491__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24515_ _24133_/CLK _16620_/X HRESETn VGND VGND VPWR VPWR _24515_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18907__A2_N _11794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21727_ _21727_/A VGND VGND VPWR VPWR _21728_/D sky130_fd_sc_hd__inv_2
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25495_ _25474_/CLK _25495_/D HRESETn VGND VGND VPWR VPWR _25495_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14925__A _24443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12460_ _12208_/X _12191_/X _12267_/Y _12459_/X VGND VGND VPWR VPWR _12461_/A sky130_fd_sc_hd__or4_4
X_21658_ _21662_/A _21658_/B VGND VGND VPWR VPWR _21658_/X sky130_fd_sc_hd__or2_4
X_24446_ _24477_/CLK _24446_/D HRESETn VGND VGND VPWR VPWR _24446_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_184_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11749__B1 _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12391_ _12264_/Y _12379_/X _12390_/X _12386_/Y VGND VGND VPWR VPWR _12391_/X sky130_fd_sc_hd__a211o_4
X_20609_ _20457_/X _20465_/B _20541_/B VGND VGND VPWR VPWR _23958_/D sky130_fd_sc_hd__o21a_4
X_21589_ _22758_/A VGND VGND VPWR VPWR _21748_/A sky130_fd_sc_hd__buf_2
X_24377_ _24377_/CLK _24377_/D HRESETn VGND VGND VPWR VPWR _17039_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_137_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14130_ _23955_/D _14129_/Y _25141_/Q _23955_/D VGND VGND VPWR VPWR _25221_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16688__B1 _15746_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23328_ _23328_/A _23327_/Y VGND VGND VPWR VPWR _23337_/B sky130_fd_sc_hd__nor2_4
XFILLER_165_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17955__B _17955_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14061_ _14024_/Y _14060_/X VGND VGND VPWR VPWR _14061_/Y sky130_fd_sc_hd__nor2_4
X_23259_ _16645_/Y _22829_/X _15556_/Y _22832_/X VGND VGND VPWR VPWR _23259_/X sky130_fd_sc_hd__o22a_4
X_13012_ _12970_/X _13010_/X _13011_/X VGND VGND VPWR VPWR _13012_/X sky130_fd_sc_hd__and3_4
XFILLER_79_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_5_6_0_HCLK_A clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17820_ _17819_/X VGND VGND VPWR VPWR _17820_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24373__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17751_ _24261_/Q VGND VGND VPWR VPWR _17752_/A sky130_fd_sc_hd__inv_2
XANTENNA__21493__A _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24302__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14963_ _15244_/A _24418_/Q _25036_/Q _14962_/Y VGND VGND VPWR VPWR _14969_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16702_ _16701_/Y _16697_/X _16522_/X _16697_/X VGND VGND VPWR VPWR _24485_/D sky130_fd_sc_hd__a2bb2o_4
X_13914_ _13914_/A VGND VGND VPWR VPWR _13914_/X sky130_fd_sc_hd__buf_2
XFILLER_236_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17682_ _17682_/A _17670_/B _17681_/Y VGND VGND VPWR VPWR _17682_/X sky130_fd_sc_hd__and3_4
X_14894_ _15214_/C _16820_/A _15062_/D _16820_/A VGND VGND VPWR VPWR _14894_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19421_ _23743_/Q VGND VGND VPWR VPWR _19421_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16612__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16633_ _16628_/A _16631_/X _16629_/Y _16632_/Y VGND VGND VPWR VPWR _16634_/A sky130_fd_sc_hd__a211o_4
XFILLER_223_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_234_0_HCLK clkbuf_8_234_0_HCLK/A VGND VGND VPWR VPWR _23976_/CLK sky130_fd_sc_hd__clkbuf_1
X_13845_ _23995_/Q VGND VGND VPWR VPWR _13845_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25508__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19352_ _19350_/Y _19348_/X _19351_/X _19348_/X VGND VGND VPWR VPWR _23767_/D sky130_fd_sc_hd__a2bb2o_4
X_16564_ _16564_/A VGND VGND VPWR VPWR _16564_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13776_ _11667_/B VGND VGND VPWR VPWR _17436_/B sky130_fd_sc_hd__buf_2
XFILLER_200_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22161__A1 _14885_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18303_ _18302_/Y _18303_/B VGND VGND VPWR VPWR _18306_/A sky130_fd_sc_hd__and2_4
XFILLER_188_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15515_ _15514_/Y _15512_/X HADDR[11] _15512_/X VGND VGND VPWR VPWR _15515_/X sky130_fd_sc_hd__a2bb2o_4
X_12727_ _12726_/X VGND VGND VPWR VPWR _12727_/Y sky130_fd_sc_hd__inv_2
X_19283_ _19290_/A VGND VGND VPWR VPWR _19283_/X sky130_fd_sc_hd__buf_2
XFILLER_231_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16495_ _16453_/A VGND VGND VPWR VPWR _16521_/A sky130_fd_sc_hd__buf_2
XFILLER_231_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18234_ _18241_/A VGND VGND VPWR VPWR _18234_/Y sky130_fd_sc_hd__inv_2
X_15446_ _13934_/C _15444_/X _15441_/X _13943_/A _15439_/X VGND VGND VPWR VPWR _15446_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_175_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12658_ _12596_/Y _12656_/A VGND VGND VPWR VPWR _12658_/X sky130_fd_sc_hd__or2_4
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18165_ _15691_/A _18149_/X _18164_/X _24245_/Q _18022_/X VGND VGND VPWR VPWR _18165_/X
+ sky130_fd_sc_hd__o32a_4
X_15377_ _24989_/Q _15376_/Y VGND VGND VPWR VPWR _15377_/X sky130_fd_sc_hd__or2_4
X_12589_ _12588_/X VGND VGND VPWR VPWR _12617_/B sky130_fd_sc_hd__buf_2
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17116_ _17062_/A _17042_/X VGND VGND VPWR VPWR _17117_/B sky130_fd_sc_hd__or2_4
XFILLER_117_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14328_ _12148_/C VGND VGND VPWR VPWR _14329_/C sky130_fd_sc_hd__inv_2
XFILLER_144_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18096_ _18128_/A _23831_/Q VGND VGND VPWR VPWR _18098_/B sky130_fd_sc_hd__or2_4
XFILLER_171_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17047_ _17062_/A _16978_/Y _17047_/C _17056_/B VGND VGND VPWR VPWR _17047_/X sky130_fd_sc_hd__or4_4
XANTENNA__15666__A _15666_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14259_ _14247_/A VGND VGND VPWR VPWR _14259_/X sky130_fd_sc_hd__buf_2
XFILLER_98_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18042__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17881__A _16917_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18998_ _17440_/A VGND VGND VPWR VPWR _18998_/X sky130_fd_sc_hd__buf_2
XANTENNA__16851__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24043__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_44_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_89_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_17949_ _17949_/A _17949_/B VGND VGND VPWR VPWR _17950_/C sky130_fd_sc_hd__or2_4
XFILLER_94_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20960_ _20822_/A _13655_/A _13655_/B _23323_/A _20874_/X VGND VGND VPWR VPWR _24066_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_226_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19619_ _19619_/A VGND VGND VPWR VPWR _21496_/B sky130_fd_sc_hd__inv_2
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20891_ _20870_/X _20890_/X _16682_/A _20875_/X VGND VGND VPWR VPWR _24049_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15957__A2 _15928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22630_ _24797_/Q _22630_/B VGND VGND VPWR VPWR _22630_/X sky130_fd_sc_hd__or2_4
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22561_ _24622_/Q _21337_/X VGND VGND VPWR VPWR _22561_/X sky130_fd_sc_hd__or2_4
XANTENNA__23123__A _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21512_ _18900_/A _21511_/X VGND VGND VPWR VPWR _21512_/X sky130_fd_sc_hd__and2_4
X_24300_ _24947_/CLK _17678_/X HRESETn VGND VGND VPWR VPWR _24300_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22492_ _22492_/A VGND VGND VPWR VPWR _22492_/Y sky130_fd_sc_hd__inv_2
X_25280_ _23528_/CLK _13742_/Y HRESETn VGND VGND VPWR VPWR _25280_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21443_ _21305_/B _21442_/X _21312_/X _24821_/Q _22523_/B VGND VGND VPWR VPWR _21443_/X
+ sky130_fd_sc_hd__a32o_4
X_24231_ _25292_/CLK _24231_/D HRESETn VGND VGND VPWR VPWR _24231_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15590__B1 _11718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22455__A2 _22282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18659__B2 _18658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24162_ _24654_/CLK _24162_/D HRESETn VGND VGND VPWR VPWR _24162_/Q sky130_fd_sc_hd__dfrtp_4
X_21374_ _21345_/Y _21356_/X _21362_/Y _21373_/Y VGND VGND VPWR VPWR _21419_/C sky130_fd_sc_hd__a211o_4
XFILLER_162_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24884__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20325_ _20324_/Y _20315_/Y _19759_/X _20315_/Y VGND VGND VPWR VPWR _20325_/X sky130_fd_sc_hd__a2bb2o_4
X_23113_ _22908_/X _23112_/X _23050_/X _11650_/A _22910_/X VGND VGND VPWR VPWR _23113_/X
+ sky130_fd_sc_hd__a32o_4
X_24093_ _23916_/CLK _20965_/X HRESETn VGND VGND VPWR VPWR _24093_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19048__A _19047_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24813__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23044_ _21864_/B VGND VGND VPWR VPWR _23044_/X sky130_fd_sc_hd__buf_2
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_126_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_126_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20256_ _21633_/B _20255_/X _19824_/A _20255_/X VGND VGND VPWR VPWR _20256_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20187_ _23471_/Q VGND VGND VPWR VPWR _20187_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16842__B1 _16522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24995_ _24551_/CLK _24995_/D HRESETn VGND VGND VPWR VPWR _15090_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22202__A _22202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21718__A1 _14391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22915__B1 _24277_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13824__A _11760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11960_ _11934_/A _11934_/B _11852_/Y VGND VGND VPWR VPWR _11961_/C sky130_fd_sc_hd__o21a_4
X_23946_ _25134_/CLK _23946_/D HRESETn VGND VGND VPWR VPWR _23946_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22391__A1 _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11891_ _11873_/X _11883_/A VGND VGND VPWR VPWR _11891_/Y sky130_fd_sc_hd__nor2_4
X_23877_ _23884_/CLK _19041_/X VGND VGND VPWR VPWR _23877_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_204_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13630_ _13630_/A _14290_/A VGND VGND VPWR VPWR _13631_/A sky130_fd_sc_hd__or2_4
X_22828_ _12428_/B _23268_/A _22827_/X VGND VGND VPWR VPWR _22828_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_64_0_HCLK clkbuf_7_32_0_HCLK/X VGND VGND VPWR VPWR _24725_/CLK sky130_fd_sc_hd__clkbuf_1
X_13561_ _13559_/A _13560_/A _13559_/Y _13560_/Y VGND VGND VPWR VPWR _13561_/X sky130_fd_sc_hd__o22a_4
X_22759_ _21431_/X _22754_/X _21832_/X _22758_/Y VGND VGND VPWR VPWR _22759_/X sky130_fd_sc_hd__a211o_4
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15300_ _15300_/A _15123_/Y _15300_/C VGND VGND VPWR VPWR _15331_/B sky130_fd_sc_hd__or3_4
X_12512_ _25427_/Q VGND VGND VPWR VPWR _12512_/Y sky130_fd_sc_hd__inv_2
X_16280_ _16275_/Y _16279_/X _15991_/X _16279_/X VGND VGND VPWR VPWR _24643_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_197_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13492_ _13492_/A VGND VGND VPWR VPWR _13492_/Y sky130_fd_sc_hd__inv_2
X_25478_ _25474_/CLK _25478_/D HRESETn VGND VGND VPWR VPWR _25478_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15476__A1_N _14876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15231_ _15039_/X _15205_/C _15194_/X _15228_/B VGND VGND VPWR VPWR _15231_/X sky130_fd_sc_hd__a211o_4
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12443_ _12443_/A _12443_/B VGND VGND VPWR VPWR _12444_/C sky130_fd_sc_hd__or2_4
X_24429_ _24462_/CLK _16825_/X HRESETn VGND VGND VPWR VPWR _24429_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15162_ _15162_/A VGND VGND VPWR VPWR _15162_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21488__A _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12374_ _12374_/A VGND VGND VPWR VPWR _12374_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14113_ _14113_/A VGND VGND VPWR VPWR _14113_/X sky130_fd_sc_hd__buf_2
XFILLER_125_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15486__A _15489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24554__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15093_ _15093_/A VGND VGND VPWR VPWR _15294_/B sky130_fd_sc_hd__inv_2
X_19970_ _19970_/A VGND VGND VPWR VPWR _19970_/X sky130_fd_sc_hd__buf_2
XANTENNA__12903__A _12741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14044_ _14523_/A _13965_/X _14049_/A _14043_/Y VGND VGND VPWR VPWR _14044_/X sky130_fd_sc_hd__o22a_4
X_18921_ _18920_/Y _18918_/X _16778_/X _18918_/X VGND VGND VPWR VPWR _23919_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21957__A1 _21939_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18852_ _16477_/Y _18739_/A _16477_/Y _18739_/A VGND VGND VPWR VPWR _18852_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17803_ _17803_/A VGND VGND VPWR VPWR _17803_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18783_ _18783_/A VGND VGND VPWR VPWR _18797_/A sky130_fd_sc_hd__buf_2
X_15995_ _24745_/Q VGND VGND VPWR VPWR _15995_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22906__B1 _24735_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17734_ _18285_/A _17726_/X _24219_/Q _17727_/Y VGND VGND VPWR VPWR _17734_/X sky130_fd_sc_hd__o22a_4
X_14946_ _14946_/A _14946_/B _14943_/X _14945_/X VGND VGND VPWR VPWR _14946_/X sky130_fd_sc_hd__or4_4
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21951__A _21936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17665_ _17575_/Y _17521_/Y _17580_/C _17665_/D VGND VGND VPWR VPWR _17666_/B sky130_fd_sc_hd__or4_4
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14877_ _14866_/X _14875_/Y _14823_/X _14876_/Y _14826_/A VGND VGND VPWR VPWR _14878_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_223_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11758__A1_N _11755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25342__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16616_ _16615_/Y _16611_/X _16435_/X _16611_/X VGND VGND VPWR VPWR _16616_/X sky130_fd_sc_hd__a2bb2o_4
X_19404_ _19402_/Y _19403_/X _19357_/X _19403_/X VGND VGND VPWR VPWR _19404_/X sky130_fd_sc_hd__a2bb2o_4
X_13828_ _13832_/A VGND VGND VPWR VPWR _13828_/X sky130_fd_sc_hd__buf_2
X_17596_ _17614_/A _17585_/X VGND VGND VPWR VPWR _17597_/B sky130_fd_sc_hd__or2_4
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23331__B1 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16547_ _16547_/A VGND VGND VPWR VPWR _16548_/A sky130_fd_sc_hd__buf_2
X_19335_ _19333_/Y _19334_/X _19200_/X _19334_/X VGND VGND VPWR VPWR _23773_/D sky130_fd_sc_hd__a2bb2o_4
X_13759_ _14664_/A VGND VGND VPWR VPWR _13807_/A sky130_fd_sc_hd__buf_2
XFILLER_204_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17010__B1 _15993_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19266_ _19253_/Y VGND VGND VPWR VPWR _19266_/X sky130_fd_sc_hd__buf_2
X_16478_ _16477_/Y _16475_/X _16301_/X _16475_/X VGND VGND VPWR VPWR _16478_/X sky130_fd_sc_hd__a2bb2o_4
X_18217_ _18053_/A _23771_/Q VGND VGND VPWR VPWR _18219_/B sky130_fd_sc_hd__or2_4
X_15429_ _15429_/A VGND VGND VPWR VPWR _15436_/B sky130_fd_sc_hd__buf_2
X_19197_ _19196_/Y _19191_/X _19106_/X _19191_/X VGND VGND VPWR VPWR _19197_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18148_ _18052_/A _18144_/X _18147_/X VGND VGND VPWR VPWR _18148_/X sky130_fd_sc_hd__or3_4
XFILLER_8_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24295__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18079_ _17990_/X _18076_/X _18079_/C VGND VGND VPWR VPWR _18079_/X sky130_fd_sc_hd__and3_4
XANTENNA__12813__A _25388_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_236_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20110_ _21397_/B _20105_/X _20109_/X _20105_/X VGND VGND VPWR VPWR _23500_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24224__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21090_ _24781_/Q _15649_/Y _21042_/X _21089_/X VGND VGND VPWR VPWR _21090_/X sky130_fd_sc_hd__a211o_4
XFILLER_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17077__B1 _17053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20041_ _20041_/A VGND VGND VPWR VPWR _20041_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18500__A _18823_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23118__A _23118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23800_ _23610_/CLK _19260_/X VGND VGND VPWR VPWR _23800_/Q sky130_fd_sc_hd__dfxtp_4
X_24780_ _24819_/CLK _24780_/D HRESETn VGND VGND VPWR VPWR _12728_/A sky130_fd_sc_hd__dfrtp_4
X_21992_ _21991_/A _20322_/Y VGND VGND VPWR VPWR _21992_/X sky130_fd_sc_hd__or2_4
XANTENNA__16020__A HWDATA[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23731_ _23747_/CLK _19452_/X VGND VGND VPWR VPWR _18209_/B sky130_fd_sc_hd__dfxtp_4
XPHY_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ _20919_/X _20942_/X _24505_/Q _20923_/X VGND VGND VPWR VPWR _24061_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25083__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _23665_/CLK _23662_/D VGND VGND VPWR VPWR _13339_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_26_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _20923_/A VGND VGND VPWR VPWR _20874_/X sky130_fd_sc_hd__buf_2
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25012__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25401_ _25403_/CLK _12727_/Y HRESETn VGND VGND VPWR VPWR _25401_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22613_ _22612_/X VGND VGND VPWR VPWR _22613_/Y sky130_fd_sc_hd__inv_2
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23593_ _23559_/CLK _19860_/X VGND VGND VPWR VPWR _19859_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_34_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14475__A _14468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17001__B1 _24726_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25332_ _23391_/CLK _25332_/D HRESETn VGND VGND VPWR VPWR _25332_/Q sky130_fd_sc_hd__dfrtp_4
X_22544_ _24045_/Q _21303_/X _13118_/A _21317_/X VGND VGND VPWR VPWR _22544_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_210_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25263_ _25089_/CLK _13823_/X HRESETn VGND VGND VPWR VPWR _13562_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17786__A _17602_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22475_ _21087_/A VGND VGND VPWR VPWR _23278_/B sky130_fd_sc_hd__buf_2
X_24214_ _23678_/CLK _24214_/D HRESETn VGND VGND VPWR VPWR _24214_/Q sky130_fd_sc_hd__dfrtp_4
X_21426_ _21298_/X VGND VGND VPWR VPWR _21427_/A sky130_fd_sc_hd__buf_2
X_25194_ _24953_/CLK _14230_/X HRESETn VGND VGND VPWR VPWR _25194_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_135_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21357_ SSn_S3 _12087_/B SSn_S2 _13482_/B VGND VGND VPWR VPWR _21357_/X sky130_fd_sc_hd__o22a_4
X_24145_ _24139_/CLK _18757_/X HRESETn VGND VGND VPWR VPWR _24145_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20308_ _20307_/X VGND VGND VPWR VPWR _22396_/B sky130_fd_sc_hd__buf_2
X_12090_ _12102_/A VGND VGND VPWR VPWR _12090_/X sky130_fd_sc_hd__buf_2
XFILLER_190_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21288_ _21288_/A _21074_/X _21288_/C _21287_/Y VGND VGND VPWR VPWR HRDATA[0] sky130_fd_sc_hd__or4_4
X_24076_ _24074_/CLK _20514_/X HRESETn VGND VGND VPWR VPWR _24076_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_150_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20239_ _20238_/Y _20234_/X _19759_/X _20227_/A VGND VGND VPWR VPWR _23451_/D sky130_fd_sc_hd__a2bb2o_4
X_23027_ _12247_/Y _22718_/X _22719_/X _12356_/Y _22846_/X VGND VGND VPWR VPWR _23027_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_131_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16815__B1 HWDATA[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23947__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14800_ _25056_/Q VGND VGND VPWR VPWR _14801_/C sky130_fd_sc_hd__inv_2
XFILLER_92_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15780_ _14366_/A _15780_/B VGND VGND VPWR VPWR _15781_/A sky130_fd_sc_hd__or2_4
X_12992_ _12282_/A _12998_/B VGND VGND VPWR VPWR _12992_/X sky130_fd_sc_hd__or2_4
X_24978_ _24980_/CLK _24978_/D HRESETn VGND VGND VPWR VPWR _24978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14731_ _14730_/X VGND VGND VPWR VPWR _14731_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11943_ _18902_/B _11942_/X VGND VGND VPWR VPWR _11944_/A sky130_fd_sc_hd__or2_4
X_23929_ _25100_/CLK _23929_/D HRESETn VGND VGND VPWR VPWR _23929_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_206_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16865__A _14777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17450_ _13247_/A _13388_/A VGND VGND VPWR VPWR _17450_/X sky130_fd_sc_hd__and2_4
X_14662_ _19116_/B _13588_/X _19141_/B VGND VGND VPWR VPWR _14662_/X sky130_fd_sc_hd__o21a_4
XFILLER_189_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11874_ RsRx_S1 _11873_/X VGND VGND VPWR VPWR _11874_/X sky130_fd_sc_hd__and2_4
XFILLER_221_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16401_ _15113_/Y _16398_/X _16400_/X _16398_/X VGND VGND VPWR VPWR _16401_/X sky130_fd_sc_hd__a2bb2o_4
X_13613_ _13613_/A _13594_/X VGND VGND VPWR VPWR _13614_/D sky130_fd_sc_hd__and2_4
X_17381_ _17239_/A _17381_/B VGND VGND VPWR VPWR _17381_/X sky130_fd_sc_hd__or2_4
X_14593_ _14552_/A _14551_/X VGND VGND VPWR VPWR _14593_/Y sky130_fd_sc_hd__nand2_4
XFILLER_198_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19120_ _19115_/Y _19119_/X _19006_/X _19119_/X VGND VGND VPWR VPWR _23850_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_213_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16332_ _16344_/A VGND VGND VPWR VPWR _16332_/X sky130_fd_sc_hd__buf_2
X_13544_ _13544_/A VGND VGND VPWR VPWR _13544_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21875__B1 _11772_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12617__B _12617_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19051_ _23873_/Q VGND VGND VPWR VPWR _19051_/Y sky130_fd_sc_hd__inv_2
X_16263_ _21335_/A VGND VGND VPWR VPWR _16263_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24735__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13475_ _13475_/A VGND VGND VPWR VPWR _13475_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_8_0_HCLK clkbuf_5_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_8_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18002_ _18222_/A _18002_/B VGND VGND VPWR VPWR _18003_/C sky130_fd_sc_hd__or2_4
XFILLER_200_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15214_ _15219_/A _15214_/B _15214_/C _15214_/D VGND VGND VPWR VPWR _15214_/X sky130_fd_sc_hd__or4_4
X_12426_ _12248_/Y _12420_/X _12390_/X _12422_/Y VGND VGND VPWR VPWR _12426_/X sky130_fd_sc_hd__a211o_4
X_16194_ _16193_/Y _16191_/X _16001_/X _16191_/X VGND VGND VPWR VPWR _16194_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23092__A2 _23083_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15145_ _24996_/Q VGND VGND VPWR VPWR _15293_/B sky130_fd_sc_hd__inv_2
XFILLER_126_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12357_ _25355_/Q VGND VGND VPWR VPWR _12357_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15076_ _15075_/Y _24605_/Q _15075_/Y _24605_/Q VGND VGND VPWR VPWR _15077_/D sky130_fd_sc_hd__a2bb2o_4
X_19953_ _19946_/A VGND VGND VPWR VPWR _19953_/X sky130_fd_sc_hd__buf_2
X_12288_ _12287_/Y _24845_/Q _12287_/Y _24845_/Q VGND VGND VPWR VPWR _12288_/X sky130_fd_sc_hd__a2bb2o_4
X_14027_ _14026_/X VGND VGND VPWR VPWR _14040_/C sky130_fd_sc_hd__inv_2
X_18904_ _11699_/A _11707_/X HWDATA[31] _24114_/Q _11708_/X VGND VGND VPWR VPWR _18904_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_68_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19884_ _19878_/Y VGND VGND VPWR VPWR _19884_/X sky130_fd_sc_hd__buf_2
XFILLER_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18835_ _18835_/A _18832_/X _18833_/X _18835_/D VGND VGND VPWR VPWR _18835_/X sky130_fd_sc_hd__or4_4
XFILLER_68_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25523__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15978_ _12219_/Y _15972_/X _15901_/X _15931_/X VGND VGND VPWR VPWR _24749_/D sky130_fd_sc_hd__a2bb2o_4
X_18766_ _18765_/X VGND VGND VPWR VPWR _24142_/D sky130_fd_sc_hd__inv_2
XFILLER_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14929_ _24423_/Q VGND VGND VPWR VPWR _14929_/Y sky130_fd_sc_hd__inv_2
X_17717_ _24212_/Q VGND VGND VPWR VPWR _21208_/A sky130_fd_sc_hd__buf_2
XFILLER_224_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18697_ _18697_/A _18696_/X VGND VGND VPWR VPWR _18697_/X sky130_fd_sc_hd__or2_4
XANTENNA__18693__C _18693_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17648_ _17648_/A _17648_/B VGND VGND VPWR VPWR _17648_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__20381__A3 _14262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17579_ _24291_/Q VGND VGND VPWR VPWR _17580_/D sky130_fd_sc_hd__inv_2
XANTENNA__20669__A1 _14215_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19318_ _19317_/Y _19313_/X _19295_/X _19299_/Y VGND VGND VPWR VPWR _19318_/X sky130_fd_sc_hd__a2bb2o_4
X_20590_ _14410_/Y _20543_/A _20556_/X _20589_/X VGND VGND VPWR VPWR _20591_/A sky130_fd_sc_hd__a211o_4
XFILLER_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24476__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19249_ _19249_/A VGND VGND VPWR VPWR _21240_/B sky130_fd_sc_hd__inv_2
X_22260_ _22007_/X _22258_/X _22260_/C VGND VGND VPWR VPWR _22260_/X sky130_fd_sc_hd__and3_4
XANTENNA__24405__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21211_ _21207_/X _21210_/X _24214_/Q VGND VGND VPWR VPWR _21212_/C sky130_fd_sc_hd__o21a_4
X_22191_ _22191_/A _21309_/A VGND VGND VPWR VPWR _22191_/X sky130_fd_sc_hd__or2_4
XFILLER_133_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21142_ _21343_/B _21141_/X _17438_/B VGND VGND VPWR VPWR _21142_/X sky130_fd_sc_hd__o21a_4
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21856__A _21856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14180__D _13765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21073_ _25520_/Q _21061_/X _21062_/X _21072_/X VGND VGND VPWR VPWR _21073_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15854__A _21064_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20024_ _20024_/A VGND VGND VPWR VPWR _21658_/B sky130_fd_sc_hd__inv_2
X_24901_ _24900_/CLK _15614_/X HRESETn VGND VGND VPWR VPWR _24901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24832_ _24866_/CLK _24832_/D HRESETn VGND VGND VPWR VPWR _24832_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_5_14_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24763_ _24763_/CLK _24763_/D HRESETn VGND VGND VPWR VPWR _24763_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21975_ _20377_/Y _21960_/B VGND VGND VPWR VPWR _21975_/X sky130_fd_sc_hd__or2_4
XFILLER_27_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23714_ _23406_/CLK _23714_/D VGND VGND VPWR VPWR _23714_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _24057_/Q _20921_/X _20925_/Y VGND VGND VPWR VPWR _20926_/Y sky130_fd_sc_hd__a21oi_4
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24694_ _24762_/CLK _24694_/D HRESETn VGND VGND VPWR VPWR _22662_/A sky130_fd_sc_hd__dfrtp_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _23644_/CLK _19709_/X VGND VGND VPWR VPWR _19706_/A sky130_fd_sc_hd__dfxtp_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ _24042_/Q _20857_/B VGND VGND VPWR VPWR _20857_/X sky130_fd_sc_hd__or2_4
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23576_ _23528_/CLK _19906_/X VGND VGND VPWR VPWR _19904_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20788_ _20780_/X _20787_/Y _15578_/A _20784_/X VGND VGND VPWR VPWR _20788_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25315_ _25474_/CLK _13487_/X HRESETn VGND VGND VPWR VPWR _25315_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22527_ _22527_/A _22686_/A VGND VGND VPWR VPWR _22528_/D sky130_fd_sc_hd__nor2_4
XFILLER_195_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15536__B1 HADDR[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21872__A3 _23075_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_138_0_HCLK clkbuf_7_69_0_HCLK/X VGND VGND VPWR VPWR _24252_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13260_ _13260_/A _13260_/B VGND VGND VPWR VPWR _13260_/X sky130_fd_sc_hd__or2_4
X_25246_ _25204_/CLK _13868_/X HRESETn VGND VGND VPWR VPWR _21559_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24146__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22458_ _16247_/Y _22454_/X _15094_/Y _22450_/X VGND VGND VPWR VPWR _22459_/B sky130_fd_sc_hd__o22a_4
XFILLER_194_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12211_ _25435_/Q VGND VGND VPWR VPWR _12211_/Y sky130_fd_sc_hd__inv_2
X_21409_ _22202_/A _20048_/Y VGND VGND VPWR VPWR _21409_/X sky130_fd_sc_hd__or2_4
X_13191_ _13249_/A VGND VGND VPWR VPWR _13396_/A sky130_fd_sc_hd__buf_2
X_25177_ _23884_/CLK _25177_/D HRESETn VGND VGND VPWR VPWR _25177_/Q sky130_fd_sc_hd__dfrtp_4
X_22389_ _21896_/X _22385_/X _22386_/X _22387_/X _22388_/X VGND VGND VPWR VPWR _22389_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_124_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12142_ _12140_/A _12141_/A _12140_/Y _12141_/Y VGND VGND VPWR VPWR _12145_/C sky130_fd_sc_hd__o22a_4
X_24128_ _25056_/CLK _18820_/X HRESETn VGND VGND VPWR VPWR _24128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15764__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12073_ _12071_/Y _12072_/X _11786_/X _12072_/X VGND VGND VPWR VPWR _25481_/D sky130_fd_sc_hd__a2bb2o_4
X_16950_ _16950_/A _16950_/B VGND VGND VPWR VPWR _16950_/X sky130_fd_sc_hd__or2_4
X_24059_ _24060_/CLK _20934_/X HRESETn VGND VGND VPWR VPWR _24059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21485__B _19893_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15901_ _18951_/A VGND VGND VPWR VPWR _15901_/X sky130_fd_sc_hd__buf_2
XFILLER_238_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16881_ _19827_/A VGND VGND VPWR VPWR _16881_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12900__B _12838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15832_ _15818_/X _15829_/X _15764_/X _24823_/Q _15786_/X VGND VGND VPWR VPWR _24823_/D
+ sky130_fd_sc_hd__a32o_4
X_18620_ _16574_/A _24144_/Q _16574_/Y _18760_/A VGND VGND VPWR VPWR _18627_/A sky130_fd_sc_hd__o22a_4
XFILLER_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22597__A _22597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15763_ _15745_/X _15761_/X _15762_/X _24859_/Q _15706_/X VGND VGND VPWR VPWR _24859_/D
+ sky130_fd_sc_hd__a32o_4
X_18551_ _18580_/A VGND VGND VPWR VPWR _18572_/A sky130_fd_sc_hd__buf_2
X_12975_ _25356_/Q VGND VGND VPWR VPWR _12975_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14714_ _14714_/A _14704_/Y _14708_/X _14713_/X VGND VGND VPWR VPWR _14715_/A sky130_fd_sc_hd__or4_4
X_17502_ _17502_/A VGND VGND VPWR VPWR _17502_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11926_ _19874_/A VGND VGND VPWR VPWR _11926_/Y sky130_fd_sc_hd__inv_2
X_18482_ _18499_/A _18499_/B VGND VGND VPWR VPWR _18483_/D sky130_fd_sc_hd__or2_4
X_15694_ _15694_/A _15691_/A VGND VGND VPWR VPWR _15694_/X sky130_fd_sc_hd__and2_4
XFILLER_61_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24987__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18961__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17433_ _17433_/A VGND VGND VPWR VPWR _17433_/Y sky130_fd_sc_hd__inv_2
X_14645_ _13615_/A VGND VGND VPWR VPWR _19387_/A sky130_fd_sc_hd__inv_2
XFILLER_32_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11857_ _11853_/X _11856_/X _11797_/A _11799_/X VGND VGND VPWR VPWR _11857_/X sky130_fd_sc_hd__a211o_4
XFILLER_220_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24916__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17364_ _17346_/A _17367_/B _17268_/X VGND VGND VPWR VPWR _17364_/Y sky130_fd_sc_hd__a21oi_4
XPHY_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14576_ _25094_/Q _14576_/B VGND VGND VPWR VPWR _14576_/X sky130_fd_sc_hd__or2_4
XANTENNA__16651__A1_N _16650_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ HWDATA[1] VGND VGND VPWR VPWR _11788_/X sky130_fd_sc_hd__buf_2
XFILLER_159_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_7_34_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_34_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15790__A3 _15710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16315_ _22821_/A VGND VGND VPWR VPWR _16315_/Y sky130_fd_sc_hd__inv_2
X_19103_ _23855_/Q VGND VGND VPWR VPWR _19103_/Y sky130_fd_sc_hd__inv_2
X_13527_ _15688_/A _13527_/B VGND VGND VPWR VPWR _14608_/A sky130_fd_sc_hd__or2_4
XFILLER_158_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15939__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15527__B1 HADDR[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_97_0_HCLK clkbuf_7_97_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_97_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17295_ _17183_/Y _17299_/B _17276_/X _17292_/B VGND VGND VPWR VPWR _17295_/X sky130_fd_sc_hd__a211o_4
XFILLER_174_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19034_ _19032_/Y _19028_/X _18985_/X _19033_/X VGND VGND VPWR VPWR _19034_/X sky130_fd_sc_hd__a2bb2o_4
X_16246_ _16244_/Y _16239_/X _16141_/X _16245_/X VGND VGND VPWR VPWR _24656_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13458_ _13458_/A VGND VGND VPWR VPWR _13458_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16036__A1_N _16035_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23934__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12409_ _12194_/Y _12413_/B _12390_/X _12405_/Y VGND VGND VPWR VPWR _12410_/A sky130_fd_sc_hd__a211o_4
XANTENNA__16666__A1_N _16665_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13459__A _13459_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16177_ _23329_/A VGND VGND VPWR VPWR _16177_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13389_ _13389_/A _23852_/Q VGND VGND VPWR VPWR _13390_/C sky130_fd_sc_hd__or2_4
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12761__B1 _12759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15128_ _24989_/Q VGND VGND VPWR VPWR _15300_/A sky130_fd_sc_hd__inv_2
XFILLER_115_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_HCLK clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_6_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_141_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15059_ _15059_/A _15265_/A _15056_/X _15058_/X VGND VGND VPWR VPWR _15059_/X sky130_fd_sc_hd__or4_4
X_19936_ _19936_/A VGND VGND VPWR VPWR _21209_/B sky130_fd_sc_hd__inv_2
XFILLER_101_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19867_ _19866_/Y _19862_/X _19613_/X _19862_/X VGND VGND VPWR VPWR _19867_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18985__A _18985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11707__A _11706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18818_ _18683_/Y _18820_/B _18817_/Y VGND VGND VPWR VPWR _24129_/D sky130_fd_sc_hd__o21a_4
XFILLER_96_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19798_ _13414_/B VGND VGND VPWR VPWR _19798_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22328__B2 _14245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18749_ _18749_/A VGND VGND VPWR VPWR _18749_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20339__B1 _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21760_ _14753_/X _21760_/B VGND VGND VPWR VPWR _21761_/C sky130_fd_sc_hd__or2_4
XANTENNA__18615__A2_N _18613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18952__B1 _18951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20711_ _15621_/Y _20708_/X _20696_/X _20710_/X VGND VGND VPWR VPWR _20712_/A sky130_fd_sc_hd__o22a_4
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15766__B1 _15472_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24657__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21691_ _13783_/D _21690_/X _18268_/A _18263_/X VGND VGND VPWR VPWR _21691_/X sky130_fd_sc_hd__o22a_4
XFILLER_168_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23430_ _23534_/CLK _23430_/D VGND VGND VPWR VPWR _23430_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_149_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20642_ _20641_/X VGND VGND VPWR VPWR _23980_/D sky130_fd_sc_hd__inv_2
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22500__B2 _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20573_ _18877_/X _20571_/Y _20572_/X VGND VGND VPWR VPWR _20573_/X sky130_fd_sc_hd__and3_4
X_23361_ _23348_/X VGND VGND VPWR VPWR IRQ[17] sky130_fd_sc_hd__buf_2
XANTENNA__14753__A _22225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25100_ _25100_/CLK _25100_/D HRESETn VGND VGND VPWR VPWR sda_oen_o_S4 sky130_fd_sc_hd__dfstp_4
X_22312_ _23176_/A _22309_/X _22311_/X VGND VGND VPWR VPWR _22394_/B sky130_fd_sc_hd__and3_4
X_23292_ _15549_/Y _23292_/B VGND VGND VPWR VPWR _23292_/X sky130_fd_sc_hd__and2_4
XFILLER_118_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21067__A1 _24714_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25031_ _25021_/CLK _25031_/D HRESETn VGND VGND VPWR VPWR _25031_/Q sky130_fd_sc_hd__dfrtp_4
X_22243_ _22251_/A _22243_/B VGND VGND VPWR VPWR _22243_/X sky130_fd_sc_hd__or2_4
XFILLER_145_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22803__A2 _22661_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22174_ _22174_/A _22174_/B _22174_/C _22173_/X VGND VGND VPWR VPWR _22174_/X sky130_fd_sc_hd__or4_4
XANTENNA__25445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21125_ _21017_/B _16268_/A _15651_/A _20684_/A _16270_/A VGND VGND VPWR VPWR _21125_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_132_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21056_ _21055_/X VGND VGND VPWR VPWR _21056_/X sky130_fd_sc_hd__buf_2
XFILLER_247_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23009__C _23075_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20007_ _20007_/A VGND VGND VPWR VPWR _21206_/B sky130_fd_sc_hd__inv_2
XFILLER_143_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14257__B1 _13788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23951__D scl_i_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24815_ _24886_/CLK _24815_/D HRESETn VGND VGND VPWR VPWR _24815_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_246_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12760_ _24809_/Q VGND VGND VPWR VPWR _12760_/Y sky130_fd_sc_hd__inv_2
X_24746_ _24639_/CLK _15994_/X HRESETn VGND VGND VPWR VPWR _15993_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _13536_/A _21958_/B VGND VGND VPWR VPWR _21958_/X sky130_fd_sc_hd__or2_4
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18943__B1 _18942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ HWDATA[20] VGND VGND VPWR VPWR _11711_/X sky130_fd_sc_hd__buf_2
XFILLER_203_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _20892_/X _20908_/X _24497_/Q _20896_/X VGND VGND VPWR VPWR _20909_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15757__B1 _15616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24398__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12569_/Y _12690_/X VGND VGND VPWR VPWR _12711_/A sky130_fd_sc_hd__or2_4
X_24677_ _24678_/CLK _16188_/X HRESETn VGND VGND VPWR VPWR _23297_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _21913_/A _20187_/Y VGND VGND VPWR VPWR _21889_/X sky130_fd_sc_hd__or2_4
XFILLER_187_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _25135_/Q VGND VGND VPWR VPWR _14430_/Y sky130_fd_sc_hd__inv_2
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628_ _23627_/CLK _19757_/X VGND VGND VPWR VPWR _19756_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24327__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23295__A2 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _25154_/Q _14349_/A _14345_/X _12078_/A _14344_/A VGND VGND VPWR VPWR _14361_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__15509__B1 HADDR[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23559_ _23559_/CLK _19949_/X VGND VGND VPWR VPWR _19948_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14663__A _25070_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16100_ _16098_/Y _16099_/X _15567_/X _16099_/X VGND VGND VPWR VPWR _16100_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _13312_/A _19725_/A VGND VGND VPWR VPWR _13312_/X sky130_fd_sc_hd__or2_4
XFILLER_11_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17080_ _17070_/A _17076_/X _17080_/C VGND VGND VPWR VPWR _17080_/X sky130_fd_sc_hd__and3_4
XFILLER_168_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14292_ _14283_/A _14283_/B _13627_/X _14291_/X VGND VGND VPWR VPWR _14293_/A sky130_fd_sc_hd__a211o_4
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16031_ _16031_/A VGND VGND VPWR VPWR _16031_/Y sky130_fd_sc_hd__inv_2
X_13243_ _11950_/A VGND VGND VPWR VPWR _13243_/X sky130_fd_sc_hd__buf_2
X_25229_ _25230_/CLK _25229_/D HRESETn VGND VGND VPWR VPWR _14005_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_182_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17974__A _18090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19120__B1 _19006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13174_ _13170_/A _20386_/A VGND VGND VPWR VPWR _13176_/B sky130_fd_sc_hd__or2_4
XFILLER_170_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22270__A3 _22265_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23962__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25186__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12125_ _12125_/A VGND VGND VPWR VPWR _12125_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15494__A _15489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17982_ _18220_/A _17973_/X _17981_/X VGND VGND VPWR VPWR _17997_/B sky130_fd_sc_hd__or3_4
XFILLER_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19721_ _19720_/Y _19718_/X _19630_/X _19718_/X VGND VGND VPWR VPWR _23641_/D sky130_fd_sc_hd__a2bb2o_4
X_12056_ _21571_/A VGND VGND VPWR VPWR _12057_/A sky130_fd_sc_hd__buf_2
X_16933_ _16126_/Y _17757_/A _16126_/Y _17757_/A VGND VGND VPWR VPWR _16934_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17434__B1 _16716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19652_ _19006_/A VGND VGND VPWR VPWR _19652_/X sky130_fd_sc_hd__buf_2
XFILLER_78_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16864_ _16858_/X VGND VGND VPWR VPWR _16864_/X sky130_fd_sc_hd__buf_2
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14248__B1 _13824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18603_ _24132_/Q VGND VGND VPWR VPWR _18686_/B sky130_fd_sc_hd__inv_2
XFILLER_237_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15815_ _15810_/X _15813_/X _15741_/X _24834_/Q _15811_/X VGND VGND VPWR VPWR _24834_/D
+ sky130_fd_sc_hd__a32o_4
X_16795_ _16791_/Y _16794_/X _15545_/X _16794_/X VGND VGND VPWR VPWR _16795_/X sky130_fd_sc_hd__a2bb2o_4
X_19583_ _21969_/D VGND VGND VPWR VPWR _19583_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19187__B1 _19144_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15746_ HWDATA[12] VGND VGND VPWR VPWR _15746_/X sky130_fd_sc_hd__buf_2
X_18534_ _18466_/C _18533_/X VGND VGND VPWR VPWR _18538_/B sky130_fd_sc_hd__or2_4
X_12958_ _12833_/C _12958_/B VGND VGND VPWR VPWR _12959_/B sky130_fd_sc_hd__or2_4
XFILLER_46_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15044__A2_N _24477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11909_ _19974_/A VGND VGND VPWR VPWR _19610_/A sky130_fd_sc_hd__buf_2
XANTENNA__24750__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15677_ _24887_/Q VGND VGND VPWR VPWR _15686_/A sky130_fd_sc_hd__inv_2
X_18465_ _18465_/A VGND VGND VPWR VPWR _18465_/Y sky130_fd_sc_hd__inv_2
X_12889_ _12967_/A VGND VGND VPWR VPWR _12889_/X sky130_fd_sc_hd__buf_2
XANTENNA__16590__A1_N _16589_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14628_ _14628_/A VGND VGND VPWR VPWR _18044_/A sky130_fd_sc_hd__buf_2
X_17416_ _20672_/A _17414_/X _17415_/X _17414_/X VGND VGND VPWR VPWR _17416_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24068__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18396_ _22163_/A _18471_/D _16195_/Y _24185_/Q VGND VGND VPWR VPWR _18398_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14420__B1 _14389_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15763__A3 _15762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17347_ _17358_/A _17352_/B _17347_/C _17352_/C VGND VGND VPWR VPWR _17348_/A sky130_fd_sc_hd__or4_4
X_14559_ _25093_/Q _14559_/B VGND VGND VPWR VPWR _14576_/B sky130_fd_sc_hd__and2_4
XFILLER_159_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17278_ _17277_/X VGND VGND VPWR VPWR _17278_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22790__A _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_121_0_HCLK clkbuf_7_60_0_HCLK/X VGND VGND VPWR VPWR _24855_/CLK sky130_fd_sc_hd__clkbuf_1
X_16229_ _16229_/A VGND VGND VPWR VPWR _16229_/X sky130_fd_sc_hd__buf_2
X_19017_ _18150_/B VGND VGND VPWR VPWR _19017_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17884__A _16917_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_184_0_HCLK clkbuf_7_92_0_HCLK/X VGND VGND VPWR VPWR _25211_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_155_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22797__A1 _21283_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17122__C1 _17053_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17673__B1 _17593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12821__A _25374_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22549__A1 _16510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19919_ _18285_/X VGND VGND VPWR VPWR _19932_/A sky130_fd_sc_hd__inv_2
XFILLER_102_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17425__B1 _16778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22930_ _16571_/A _22884_/X _22928_/X _22929_/X VGND VGND VPWR VPWR _22930_/X sky130_fd_sc_hd__a211o_4
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22861_ _22861_/A _22901_/B VGND VGND VPWR VPWR _22861_/X sky130_fd_sc_hd__or2_4
XANTENNA__24838__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19178__B1 _19063_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24600_ _24520_/CLK _16396_/X HRESETn VGND VGND VPWR VPWR _24600_/Q sky130_fd_sc_hd__dfrtp_4
X_21812_ _21808_/X _21811_/X _21489_/X VGND VGND VPWR VPWR _21812_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17124__A _17020_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22792_ _22786_/X _22788_/X _22789_/X _22791_/X VGND VGND VPWR VPWR _22793_/B sky130_fd_sc_hd__o22a_4
XFILLER_225_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22965__A _22942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24531_ _24540_/CLK _24531_/D HRESETn VGND VGND VPWR VPWR _16578_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__23117__A1_N _17236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21743_ _16366_/B _21740_/X _16180_/X _21742_/X VGND VGND VPWR VPWR _21744_/B sky130_fd_sc_hd__o22a_4
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24491__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22684__B _22684_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24462_ _24462_/CLK _24462_/D HRESETn VGND VGND VPWR VPWR _14998_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24420__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21674_ _21207_/A VGND VGND VPWR VPWR _21674_/X sky130_fd_sc_hd__buf_2
XFILLER_197_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14411__B1 _14380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23413_ _23678_/CLK _23413_/D VGND VGND VPWR VPWR _20338_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20625_ _17386_/X _20624_/Y _20621_/C VGND VGND VPWR VPWR _20625_/X sky130_fd_sc_hd__and3_4
XANTENNA__12418__D _12370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24393_ _24390_/CLK _24393_/D HRESETn VGND VGND VPWR VPWR _24393_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23344_ _25271_/Q _23343_/X VGND VGND VPWR VPWR _23344_/X sky130_fd_sc_hd__and2_4
X_20556_ _14096_/A VGND VGND VPWR VPWR _20556_/X sky130_fd_sc_hd__buf_2
XANTENNA__16164__B1 _15475_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23029__A2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_80_0_HCLK clkbuf_7_81_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_80_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23275_ _23275_/A _22658_/B VGND VGND VPWR VPWR _23275_/X sky130_fd_sc_hd__or2_4
X_20487_ _20516_/A _20483_/X _20486_/Y VGND VGND VPWR VPWR _20488_/B sky130_fd_sc_hd__o21a_4
XFILLER_3_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19102__B1 _18985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25014_ _24967_/CLK _25014_/D HRESETn VGND VGND VPWR VPWR _25014_/Q sky130_fd_sc_hd__dfrtp_4
X_22226_ _22226_/A _22224_/X _22225_/X VGND VGND VPWR VPWR _22227_/C sky130_fd_sc_hd__and3_4
XFILLER_105_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22205__A _22205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22157_ _22157_/A _22157_/B VGND VGND VPWR VPWR _22158_/D sky130_fd_sc_hd__and2_4
XFILLER_105_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21108_ _21040_/X _21106_/X _21047_/X _21107_/X VGND VGND VPWR VPWR _21109_/C sky130_fd_sc_hd__a211o_4
X_22088_ _21773_/X _22087_/X _14710_/A VGND VGND VPWR VPWR _22088_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_154_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17416__B1 _17415_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13930_ _13930_/A VGND VGND VPWR VPWR _13932_/B sky130_fd_sc_hd__inv_2
XFILLER_59_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21039_ _21038_/X VGND VGND VPWR VPWR _21128_/B sky130_fd_sc_hd__buf_2
XFILLER_87_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22960__B2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13861_ _25249_/Q _13850_/X _25248_/Q _13852_/X VGND VGND VPWR VPWR _13861_/X sky130_fd_sc_hd__o22a_4
XFILLER_219_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24579__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15978__B1 _15901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15600_ _15600_/A VGND VGND VPWR VPWR _22683_/A sky130_fd_sc_hd__inv_2
X_12812_ _24807_/Q VGND VGND VPWR VPWR _12812_/Y sky130_fd_sc_hd__inv_2
X_16580_ _16598_/A VGND VGND VPWR VPWR _16580_/X sky130_fd_sc_hd__buf_2
XANTENNA__24508__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13792_ _13792_/A VGND VGND VPWR VPWR _13792_/X sky130_fd_sc_hd__buf_2
XFILLER_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14393__A1_N _14391_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18916__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15531_ _13457_/D _15530_/X HADDR[4] _15530_/X VGND VGND VPWR VPWR _15531_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_215_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12743_ _22553_/A VGND VGND VPWR VPWR _12743_/Y sky130_fd_sc_hd__inv_2
X_24729_ _24357_/CLK _24729_/D HRESETn VGND VGND VPWR VPWR _16040_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12178__A _22558_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18250_ HWDATA[7] VGND VGND VPWR VPWR _18250_/X sky130_fd_sc_hd__buf_2
XFILLER_242_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15462_ _24956_/Q VGND VGND VPWR VPWR _15462_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24161__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12674_ _12677_/A _12668_/B _12673_/Y VGND VGND VPWR VPWR _12674_/X sky130_fd_sc_hd__and3_4
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _22821_/A _17200_/Y _16346_/Y _24346_/Q VGND VGND VPWR VPWR _17201_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14412_/Y _14408_/X _14392_/X _14408_/X VGND VGND VPWR VPWR _14413_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18181_ _13617_/X _18173_/X _18180_/X VGND VGND VPWR VPWR _18181_/X sky130_fd_sc_hd__and3_4
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15489__A _15489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _15390_/A _15390_/B VGND VGND VPWR VPWR _15393_/Y sky130_fd_sc_hd__nand2_4
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17132_ _17038_/D _17131_/X VGND VGND VPWR VPWR _17132_/X sky130_fd_sc_hd__or2_4
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ _14344_/A VGND VGND VPWR VPWR _14344_/X sky130_fd_sc_hd__buf_2
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17063_ _17023_/Y _17045_/X _16965_/Y _17062_/X VGND VGND VPWR VPWR _17063_/X sky130_fd_sc_hd__or4_4
XFILLER_195_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25367__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14275_ _13509_/A _14290_/A VGND VGND VPWR VPWR _25183_/D sky130_fd_sc_hd__and2_4
XFILLER_183_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15902__B1 _15901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22779__A1 _11681_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16014_ _16014_/A VGND VGND VPWR VPWR _16014_/Y sky130_fd_sc_hd__inv_2
X_13226_ _13374_/A _23793_/Q VGND VGND VPWR VPWR _13229_/B sky130_fd_sc_hd__or2_4
XFILLER_98_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21451__A1 _23328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13157_ _13167_/A VGND VGND VPWR VPWR _13157_/X sky130_fd_sc_hd__buf_2
XANTENNA__12641__A _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14469__B1 _14407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12108_ _12106_/Y _12102_/X _11786_/X _12107_/X VGND VGND VPWR VPWR _25471_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21954__A _21954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13088_ _13072_/B _13088_/B _13091_/C VGND VGND VPWR VPWR _25341_/D sky130_fd_sc_hd__and3_4
X_17965_ _17947_/X _17962_/X _18024_/A _24249_/Q _17966_/A VGND VGND VPWR VPWR _24249_/D
+ sky130_fd_sc_hd__a32o_4
X_19704_ _13346_/B VGND VGND VPWR VPWR _19704_/Y sky130_fd_sc_hd__inv_2
X_12039_ _16364_/A _15636_/B _15636_/C _12039_/D VGND VGND VPWR VPWR _21574_/B sky130_fd_sc_hd__or4_4
X_16916_ _22494_/A _16915_/A _16140_/Y _16915_/Y VGND VGND VPWR VPWR _16919_/C sky130_fd_sc_hd__o22a_4
X_17896_ _21991_/A VGND VGND VPWR VPWR _17896_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19635_ _19632_/Y _19627_/X _19633_/X _19634_/X VGND VGND VPWR VPWR _23672_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15671__B _15670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16847_ _16847_/A VGND VGND VPWR VPWR _16847_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15969__B1 _15754_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24931__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24249__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19566_ _19566_/A VGND VGND VPWR VPWR _21192_/B sky130_fd_sc_hd__inv_2
XFILLER_241_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16778_ _18942_/A VGND VGND VPWR VPWR _16778_/X sky130_fd_sc_hd__buf_2
XFILLER_92_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_5_23_0_HCLK_A clkbuf_5_23_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22785__A _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22703__A1 _24428_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18907__B1 HWDATA[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18517_ _18510_/X VGND VGND VPWR VPWR _18521_/B sky130_fd_sc_hd__inv_2
XFILLER_240_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15729_ _12514_/Y _15728_/X _15581_/X _15728_/X VGND VGND VPWR VPWR _24876_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19497_ _19496_/Y _19494_/X _11927_/X _19494_/X VGND VGND VPWR VPWR _19497_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20714__B1 _20696_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18448_ _16187_/Y _24188_/Q _16187_/Y _24188_/Q VGND VGND VPWR VPWR _18448_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16394__B1 _16020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18379_ _18373_/Y VGND VGND VPWR VPWR _18379_/X sky130_fd_sc_hd__buf_2
XFILLER_119_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__19332__B1 _19221_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20410_ _20409_/Y VGND VGND VPWR VPWR _20410_/X sky130_fd_sc_hd__buf_2
XFILLER_175_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21390_ _22196_/A _21388_/X _21389_/X VGND VGND VPWR VPWR _21390_/X sky130_fd_sc_hd__and3_4
XANTENNA__16146__B1 _16145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13540__A1_N _13538_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20341_ _20328_/Y VGND VGND VPWR VPWR _20341_/X sky130_fd_sc_hd__buf_2
XFILLER_128_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25037__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20272_ _20266_/Y VGND VGND VPWR VPWR _20272_/X sky130_fd_sc_hd__buf_2
X_23060_ _23060_/A _23060_/B VGND VGND VPWR VPWR _23060_/Y sky130_fd_sc_hd__nor2_4
XFILLER_162_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22011_ _22015_/A VGND VGND VPWR VPWR _22020_/A sky130_fd_sc_hd__buf_2
XFILLER_103_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12551__A _12551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21286__D _21285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21864__A _15022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19399__B1 _19351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15862__A _15861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23962_ _24146_/CLK _23962_/D HRESETn VGND VGND VPWR VPWR _23962_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22913_ _22781_/A _22900_/X _22913_/C _22912_/X VGND VGND VPWR VPWR _22913_/X sky130_fd_sc_hd__or4_4
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24672__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23893_ _23887_/CLK _23893_/D VGND VGND VPWR VPWR _18154_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__14478__A HWDATA[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22844_ _22844_/A _22837_/X _22844_/C VGND VGND VPWR VPWR _22844_/X sky130_fd_sc_hd__and3_4
XANTENNA__24601__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15975__A3 _15764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22775_ _24628_/Q _22487_/X VGND VGND VPWR VPWR _22775_/X sky130_fd_sc_hd__or2_4
XFILLER_13_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24514_ _24679_/CLK _24514_/D HRESETn VGND VGND VPWR VPWR _13727_/A sky130_fd_sc_hd__dfrtp_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21726_ _14205_/Y _14182_/X _14222_/Y _21351_/X VGND VGND VPWR VPWR _21727_/A sky130_fd_sc_hd__o22a_4
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25494_ _25474_/CLK _25494_/D HRESETn VGND VGND VPWR VPWR _25494_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16385__B1 _16295_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20181__B2 _20180_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24445_ _24477_/CLK _16795_/X HRESETn VGND VGND VPWR VPWR _24445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21657_ _21657_/A _19868_/Y VGND VGND VPWR VPWR _21657_/X sky130_fd_sc_hd__or2_4
XFILLER_200_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19323__B1 _19301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20608_ _20603_/X _20607_/X _20541_/B VGND VGND VPWR VPWR _20608_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16137__B1 _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12390_ _12415_/A VGND VGND VPWR VPWR _12390_/X sky130_fd_sc_hd__buf_2
X_24376_ _24725_/CLK _24376_/D HRESETn VGND VGND VPWR VPWR _17036_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_177_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21588_ _21588_/A VGND VGND VPWR VPWR _22758_/A sky130_fd_sc_hd__buf_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23327_ _13126_/A _21292_/X _13655_/A _21315_/X VGND VGND VPWR VPWR _23327_/Y sky130_fd_sc_hd__a22oi_4
X_20539_ _20539_/A _23927_/Q VGND VGND VPWR VPWR _23923_/D sky130_fd_sc_hd__and2_4
XFILLER_192_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14060_ _14043_/Y _14060_/B _14039_/X _14004_/X VGND VGND VPWR VPWR _14060_/X sky130_fd_sc_hd__or4_4
X_23258_ _20952_/Y _21597_/A _20813_/Y _22290_/A VGND VGND VPWR VPWR _23258_/X sky130_fd_sc_hd__o22a_4
XFILLER_152_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13011_ _12285_/Y _13008_/X VGND VGND VPWR VPWR _13011_/X sky130_fd_sc_hd__or2_4
X_22209_ _22209_/A _22209_/B VGND VGND VPWR VPWR _22211_/B sky130_fd_sc_hd__or2_4
XFILLER_106_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23189_ _23280_/A _23189_/B VGND VGND VPWR VPWR _23196_/C sky130_fd_sc_hd__and2_4
Xclkbuf_8_24_0_HCLK clkbuf_7_12_0_HCLK/X VGND VGND VPWR VPWR _23678_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_87_0_HCLK clkbuf_8_87_0_HCLK/A VGND VGND VPWR VPWR _25341_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14962_ _14962_/A VGND VGND VPWR VPWR _14962_/Y sky130_fd_sc_hd__inv_2
X_17750_ _17747_/Y _16925_/Y _17748_/Y _17750_/D VGND VGND VPWR VPWR _17750_/X sky130_fd_sc_hd__or4_4
XFILLER_121_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16701_ _16701_/A VGND VGND VPWR VPWR _16701_/Y sky130_fd_sc_hd__inv_2
X_13913_ _24973_/Q VGND VGND VPWR VPWR _13913_/X sky130_fd_sc_hd__buf_2
XFILLER_207_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14893_ _15062_/D VGND VGND VPWR VPWR _15214_/C sky130_fd_sc_hd__buf_2
X_17681_ _17513_/Y _17669_/B VGND VGND VPWR VPWR _17681_/Y sky130_fd_sc_hd__nand2_4
XFILLER_235_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19420_ _19418_/Y _19413_/X _19395_/X _19419_/X VGND VGND VPWR VPWR _23744_/D sky130_fd_sc_hd__a2bb2o_4
X_13844_ _13840_/C VGND VGND VPWR VPWR _13844_/X sky130_fd_sc_hd__buf_2
X_16632_ _16170_/B _16632_/B VGND VGND VPWR VPWR _16632_/Y sky130_fd_sc_hd__nor2_4
XFILLER_235_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24342__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19351_ _18942_/A VGND VGND VPWR VPWR _19351_/X sky130_fd_sc_hd__buf_2
X_13775_ _14180_/A VGND VGND VPWR VPWR _21138_/A sky130_fd_sc_hd__buf_2
X_16563_ _16562_/Y _16560_/X _16301_/X _16560_/X VGND VGND VPWR VPWR _16563_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22161__A2 _22807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17010__A2_N _24403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18302_ _18292_/X VGND VGND VPWR VPWR _18302_/Y sky130_fd_sc_hd__inv_2
X_12726_ _12689_/A _12626_/D _12627_/X _12724_/B VGND VGND VPWR VPWR _12726_/X sky130_fd_sc_hd__a211o_4
X_15514_ _11673_/A VGND VGND VPWR VPWR _15514_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18904__A3 HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16494_ _16494_/A VGND VGND VPWR VPWR _16494_/Y sky130_fd_sc_hd__inv_2
X_19282_ _18985_/A VGND VGND VPWR VPWR _19282_/X sky130_fd_sc_hd__buf_2
XFILLER_130_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15445_ _13943_/A _15444_/X _15441_/X _13932_/C _15439_/X VGND VGND VPWR VPWR _15445_/X
+ sky130_fd_sc_hd__a32o_4
X_18233_ _21962_/A _20369_/A VGND VGND VPWR VPWR _18241_/A sky130_fd_sc_hd__or2_4
X_12657_ _12657_/A _12657_/B VGND VGND VPWR VPWR _12659_/B sky130_fd_sc_hd__or2_4
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12636__A _12627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__19314__B1 _19200_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15012__A _24476_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15376_ _15376_/A VGND VGND VPWR VPWR _15376_/Y sky130_fd_sc_hd__inv_2
X_18164_ _18132_/A _18156_/X _18164_/C VGND VGND VPWR VPWR _18164_/X sky130_fd_sc_hd__and3_4
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ _12588_/A _12588_/B VGND VGND VPWR VPWR _12588_/X sky130_fd_sc_hd__or2_4
XFILLER_184_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ _14338_/A VGND VGND VPWR VPWR _14334_/A sky130_fd_sc_hd__inv_2
X_17115_ _17087_/A VGND VGND VPWR VPWR _17142_/A sky130_fd_sc_hd__buf_2
XFILLER_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18095_ _18095_/A VGND VGND VPWR VPWR _18098_/A sky130_fd_sc_hd__buf_2
XFILLER_171_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17046_ _17023_/Y _17045_/X VGND VGND VPWR VPWR _17056_/B sky130_fd_sc_hd__or2_4
X_14258_ _25187_/Q VGND VGND VPWR VPWR _21557_/A sky130_fd_sc_hd__inv_2
XFILLER_171_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13209_ _13365_/A _13209_/B _13209_/C VGND VGND VPWR VPWR _13209_/X sky130_fd_sc_hd__and3_4
XFILLER_171_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22621__B1 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14189_ _14189_/A VGND VGND VPWR VPWR _14190_/A sky130_fd_sc_hd__buf_2
XFILLER_171_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12371__A _12370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18997_ _18218_/B VGND VGND VPWR VPWR _18997_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17948_ _18016_/A _17948_/B VGND VGND VPWR VPWR _17950_/B sky130_fd_sc_hd__or2_4
XFILLER_239_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17879_ _17878_/X VGND VGND VPWR VPWR _17879_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19618_ _21684_/B _19616_/X _19617_/X _19616_/X VGND VGND VPWR VPWR _23677_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11715__A HWDATA[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24083__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20890_ _20887_/Y _20888_/Y _20889_/X VGND VGND VPWR VPWR _20890_/X sky130_fd_sc_hd__o21a_4
XANTENNA__15957__A3 HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24012__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19549_ _19548_/X VGND VGND VPWR VPWR _19549_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22688__B1 _22687_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22560_ _21294_/X _22558_/X _21300_/A _24830_/Q _22559_/X VGND VGND VPWR VPWR _22560_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_179_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14745__B _14739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21511_ _13771_/A VGND VGND VPWR VPWR _21511_/X sky130_fd_sc_hd__buf_2
XANTENNA__25289__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22491_ _22486_/X _22488_/X _22489_/X _24725_/Q _22490_/X VGND VGND VPWR VPWR _22492_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_167_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16018__A _24737_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24230_ _24233_/CLK _18255_/X HRESETn VGND VGND VPWR VPWR _24230_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21442_ _21442_/A _21441_/X VGND VGND VPWR VPWR _21442_/X sky130_fd_sc_hd__or2_4
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16119__B1 _15951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22455__A3 _16724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12265__B _12194_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24161_ _24325_/CLK _18591_/X HRESETn VGND VGND VPWR VPWR _24161_/Q sky130_fd_sc_hd__dfrtp_4
X_21373_ _21556_/A _21372_/X VGND VGND VPWR VPWR _21373_/Y sky130_fd_sc_hd__nor2_4
XFILLER_175_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23112_ _23112_/A _22909_/B VGND VGND VPWR VPWR _23112_/X sky130_fd_sc_hd__or2_4
X_20324_ _21214_/A VGND VGND VPWR VPWR _20324_/Y sky130_fd_sc_hd__inv_2
X_24092_ _25308_/CLK _20964_/X HRESETn VGND VGND VPWR VPWR _11977_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_190_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23043_ _23043_/A _23043_/B VGND VGND VPWR VPWR _23053_/C sky130_fd_sc_hd__and2_4
XFILLER_150_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20255_ _20243_/A VGND VGND VPWR VPWR _20255_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_240_0_HCLK clkbuf_8_241_0_HCLK/A VGND VGND VPWR VPWR _24539_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_103_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20186_ _22063_/B _20180_/X _20095_/X _20185_/X VGND VGND VPWR VPWR _20186_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24853__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12501__A2_N _24886_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24994_ _24551_/CLK _24994_/D HRESETn VGND VGND VPWR VPWR _24994_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_130_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23945_ _25140_/CLK _20583_/Y HRESETn VGND VGND VPWR VPWR _23945_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19792__B1 _19702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11890_ _11848_/A _11888_/X _11883_/A _11889_/Y VGND VGND VPWR VPWR _25512_/D sky130_fd_sc_hd__o22a_4
X_23876_ _23884_/CLK _19043_/X VGND VGND VPWR VPWR _23876_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22827_ _12838_/B _21446_/X _16921_/Y _22826_/X VGND VGND VPWR VPWR _22827_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22856__C _22845_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19544__B1 _19543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23340__B2 _25057_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13560_ _13560_/A VGND VGND VPWR VPWR _13560_/Y sky130_fd_sc_hd__inv_2
X_25546_ _24626_/CLK _25546_/D HRESETn VGND VGND VPWR VPWR _25546_/Q sky130_fd_sc_hd__dfrtp_4
X_22758_ _22758_/A _22758_/B VGND VGND VPWR VPWR _22758_/Y sky130_fd_sc_hd__nor2_4
XFILLER_240_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12511_ _12511_/A VGND VGND VPWR VPWR _12511_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21709_ _22279_/A _21707_/X _21541_/X _24719_/Q _21708_/X VGND VGND VPWR VPWR _21709_/X
+ sky130_fd_sc_hd__a32o_4
X_13491_ _13490_/Y _13488_/X _11765_/X _13488_/X VGND VGND VPWR VPWR _25313_/D sky130_fd_sc_hd__a2bb2o_4
X_25477_ _25474_/CLK _25477_/D HRESETn VGND VGND VPWR VPWR _25477_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_212_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22689_ _20748_/Y _23129_/A _15598_/Y _22279_/X VGND VGND VPWR VPWR _22689_/X sky130_fd_sc_hd__o22a_4
X_15230_ _15203_/X _15230_/B _15230_/C VGND VGND VPWR VPWR _25023_/D sky130_fd_sc_hd__and3_4
X_12442_ _12236_/A _12442_/B VGND VGND VPWR VPWR _12444_/B sky130_fd_sc_hd__or2_4
X_24428_ _24462_/CLK _16828_/X HRESETn VGND VGND VPWR VPWR _24428_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20673__A _20673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15161_ _15168_/A _15168_/B _14972_/Y _15161_/D VGND VGND VPWR VPWR _15162_/A sky130_fd_sc_hd__or4_4
XFILLER_172_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12373_ _12204_/Y _12264_/Y _12254_/Y _12385_/B VGND VGND VPWR VPWR _12374_/A sky130_fd_sc_hd__or4_4
X_24359_ _24629_/CLK _17320_/X HRESETn VGND VGND VPWR VPWR _17179_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22851__B1 _11720_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14671__A _22069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_50_0_HCLK clkbuf_6_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_50_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14112_ _14111_/X _14099_/A VGND VGND VPWR VPWR _14113_/A sky130_fd_sc_hd__and2_4
XFILLER_153_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15092_ _15090_/A _15091_/A _15291_/A _15091_/Y VGND VGND VPWR VPWR _15102_/A sky130_fd_sc_hd__o22a_4
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14043_ _14042_/X VGND VGND VPWR VPWR _14043_/Y sky130_fd_sc_hd__inv_2
X_18920_ _18920_/A VGND VGND VPWR VPWR _18920_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22603__B1 _25531_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21957__A2 _21954_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18851_ _18847_/X _18848_/X _18849_/X _18850_/X VGND VGND VPWR VPWR _18851_/X sky130_fd_sc_hd__or4_4
XANTENNA__24594__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17802_ _16906_/Y _17796_/X _17783_/X _17798_/Y VGND VGND VPWR VPWR _17803_/A sky130_fd_sc_hd__a211o_4
XFILLER_121_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24523__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18782_ _18744_/A VGND VGND VPWR VPWR _18793_/A sky130_fd_sc_hd__buf_2
X_15994_ _15993_/Y _15990_/X _15554_/X _15990_/X VGND VGND VPWR VPWR _15994_/X sky130_fd_sc_hd__a2bb2o_4
X_17733_ _17732_/Y VGND VGND VPWR VPWR _18285_/A sky130_fd_sc_hd__buf_2
X_14945_ _14944_/Y _24428_/Q _14944_/Y _24428_/Q VGND VGND VPWR VPWR _14945_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12855__C1 _12854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19702__A _11774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17664_ _17559_/Y _17580_/D VGND VGND VPWR VPWR _17665_/D sky130_fd_sc_hd__or2_4
XFILLER_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14876_ _24951_/Q VGND VGND VPWR VPWR _14876_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19403_ _19388_/Y VGND VGND VPWR VPWR _19403_/X sky130_fd_sc_hd__buf_2
X_16615_ _16615_/A VGND VGND VPWR VPWR _16615_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13827_ _13538_/Y _13822_/X _13826_/X _13822_/X VGND VGND VPWR VPWR _13827_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17595_ _17595_/A VGND VGND VPWR VPWR _17595_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23331__A1 _24546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19535__B1 _19534_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19334_ _19327_/A VGND VGND VPWR VPWR _19334_/X sky130_fd_sc_hd__buf_2
XFILLER_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13758_ _13757_/Y VGND VGND VPWR VPWR _13758_/X sky130_fd_sc_hd__buf_2
X_16546_ _24544_/Q VGND VGND VPWR VPWR _16546_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12709_ _12680_/A VGND VGND VPWR VPWR _12722_/C sky130_fd_sc_hd__buf_2
XANTENNA__17010__B2 _24403_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25382__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19265_ _23797_/Q VGND VGND VPWR VPWR _21614_/B sky130_fd_sc_hd__inv_2
X_13689_ _13686_/A _13686_/B VGND VGND VPWR VPWR _13689_/Y sky130_fd_sc_hd__nand2_4
X_16477_ _16477_/A VGND VGND VPWR VPWR _16477_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25406__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18216_ _17990_/X _18214_/X _18215_/X VGND VGND VPWR VPWR _18216_/X sky130_fd_sc_hd__and3_4
XANTENNA__25311__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15428_ _15425_/X VGND VGND VPWR VPWR _15429_/A sky130_fd_sc_hd__inv_2
X_19196_ _23822_/Q VGND VGND VPWR VPWR _19196_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15359_ _15291_/A _15357_/X _15358_/Y VGND VGND VPWR VPWR _24995_/D sky130_fd_sc_hd__o21a_4
X_18147_ _17968_/X _18145_/X _18147_/C VGND VGND VPWR VPWR _18147_/X sky130_fd_sc_hd__and3_4
XFILLER_129_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18078_ _18146_/A _18078_/B VGND VGND VPWR VPWR _18079_/C sky130_fd_sc_hd__or2_4
XFILLER_172_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17029_ _17029_/A VGND VGND VPWR VPWR _17030_/D sky130_fd_sc_hd__inv_2
X_20040_ _20038_/Y _20034_/X _19813_/X _20039_/X VGND VGND VPWR VPWR _20040_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18906__A2_N _11794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24264__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16301__A HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_70_0_HCLK clkbuf_8_70_0_HCLK/A VGND VGND VPWR VPWR _24278_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_67_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22022__B _19945_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21991_ _21991_/A _20322_/Y VGND VGND VPWR VPWR _21991_/X sky130_fd_sc_hd__and2_4
X_23730_ _23406_/CLK _23730_/D VGND VGND VPWR VPWR _23730_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12310__B2 _12309_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _20939_/Y _20940_/Y _20941_/X VGND VGND VPWR VPWR _20942_/X sky130_fd_sc_hd__o21a_4
XFILLER_215_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16588__B1 _16233_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23661_ _24209_/CLK _23661_/D VGND VGND VPWR VPWR _13371_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _20824_/A VGND VGND VPWR VPWR _20923_/A sky130_fd_sc_hd__inv_2
XFILLER_242_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25400_ _24819_/CLK _25400_/D HRESETn VGND VGND VPWR VPWR _21015_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_242_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23322__A1 _12167_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22612_ _22596_/Y _22601_/Y _22609_/Y _21445_/X _22611_/X VGND VGND VPWR VPWR _22612_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23592_ _23559_/CLK _23592_/D VGND VGND VPWR VPWR _19861_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22973__A _21427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25331_ _23456_/CLK _13283_/X HRESETn VGND VGND VPWR VPWR _25331_/Q sky130_fd_sc_hd__dfrtp_4
X_22543_ _22543_/A VGND VGND VPWR VPWR _22543_/X sky130_fd_sc_hd__buf_2
XFILLER_194_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25052__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25262_ _25260_/CLK _25262_/D HRESETn VGND VGND VPWR VPWR _13544_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_195_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22474_ _21537_/X VGND VGND VPWR VPWR _22474_/X sky130_fd_sc_hd__buf_2
X_24213_ _24302_/CLK _24213_/D HRESETn VGND VGND VPWR VPWR _24213_/Q sky130_fd_sc_hd__dfrtp_4
X_21425_ _21425_/A _22420_/B VGND VGND VPWR VPWR _21425_/X sky130_fd_sc_hd__or2_4
X_25193_ _24973_/CLK _14241_/X HRESETn VGND VGND VPWR VPWR sda_oen_o_S5 sky130_fd_sc_hd__dfstp_4
XANTENNA__23300__C _23299_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24144_ _24139_/CLK _18761_/X HRESETn VGND VGND VPWR VPWR _24144_/Q sky130_fd_sc_hd__dfrtp_4
X_21356_ _21347_/X _21356_/B _21356_/C _21355_/Y VGND VGND VPWR VPWR _21356_/X sky130_fd_sc_hd__or4_4
XFILLER_107_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20307_ _19570_/X VGND VGND VPWR VPWR _20307_/X sky130_fd_sc_hd__buf_2
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24075_ _24074_/CLK _20531_/X HRESETn VGND VGND VPWR VPWR _24075_/Q sky130_fd_sc_hd__dfrtp_4
X_21287_ _21287_/A VGND VGND VPWR VPWR _21287_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23026_ _22824_/X _23017_/Y _23021_/Y _23025_/X VGND VGND VPWR VPWR _23034_/C sky130_fd_sc_hd__a211o_4
X_20238_ _13424_/B VGND VGND VPWR VPWR _20238_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22213__A _22213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22600__A3 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20169_ _20168_/Y _20164_/X _20102_/X _20164_/X VGND VGND VPWR VPWR _23478_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12991_ _12993_/B VGND VGND VPWR VPWR _12998_/B sky130_fd_sc_hd__inv_2
X_24977_ _24976_/CLK _15418_/X HRESETn VGND VGND VPWR VPWR _15417_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_18_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11942_ _11935_/X _11942_/B VGND VGND VPWR VPWR _11942_/X sky130_fd_sc_hd__or2_4
X_14730_ _22048_/A _14702_/X _14729_/A _14701_/A VGND VGND VPWR VPWR _14730_/X sky130_fd_sc_hd__o22a_4
XFILLER_18_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19522__A _19522_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23928_ _25100_/CLK _23928_/D HRESETn VGND VGND VPWR VPWR _23928_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23987__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14661_ _19411_/A _19141_/B _19411_/A _19141_/B VGND VGND VPWR VPWR _25072_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23044__A _21864_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11873_ _11872_/X VGND VGND VPWR VPWR _11873_/X sky130_fd_sc_hd__buf_2
X_23859_ _23859_/CLK _23859_/D VGND VGND VPWR VPWR _23859_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14666__A _14672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13612_ _13612_/A VGND VGND VPWR VPWR _13613_/A sky130_fd_sc_hd__buf_2
X_16400_ HWDATA[18] VGND VGND VPWR VPWR _16400_/X sky130_fd_sc_hd__buf_2
XFILLER_232_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14592_ _14554_/B _14590_/Y _14588_/X _14591_/X _25088_/Q VGND VGND VPWR VPWR _14592_/X
+ sky130_fd_sc_hd__a32o_4
X_17380_ _17341_/A _17374_/B _17379_/Y VGND VGND VPWR VPWR _17380_/X sky130_fd_sc_hd__and3_4
XANTENNA__22883__A _22883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13543_ _22734_/A _25098_/Q _22734_/A _25098_/Q VGND VGND VPWR VPWR _13543_/X sky130_fd_sc_hd__a2bb2o_4
X_16331_ _24623_/Q VGND VGND VPWR VPWR _16331_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21875__A1 _16154_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25529_ _25524_/CLK _11754_/X HRESETn VGND VGND VPWR VPWR _25529_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21875__B2 _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16262_ _16261_/Y _16257_/X _15976_/X _16257_/X VGND VGND VPWR VPWR _24649_/D sky130_fd_sc_hd__a2bb2o_4
X_19050_ _19046_/Y _19049_/X _19006_/X _19049_/X VGND VGND VPWR VPWR _23874_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21499__A _17731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13474_ _13473_/Y _13469_/X _11781_/X _13469_/X VGND VGND VPWR VPWR _25320_/D sky130_fd_sc_hd__a2bb2o_4
X_15213_ _15212_/X VGND VGND VPWR VPWR _15213_/Y sky130_fd_sc_hd__inv_2
X_18001_ _18054_/A VGND VGND VPWR VPWR _18222_/A sky130_fd_sc_hd__buf_2
X_12425_ _12434_/A _12425_/B _12424_/X VGND VGND VPWR VPWR _12425_/X sky130_fd_sc_hd__and3_4
X_16193_ _23238_/A VGND VGND VPWR VPWR _16193_/Y sky130_fd_sc_hd__inv_2
X_15144_ _24602_/Q VGND VGND VPWR VPWR _15144_/Y sky130_fd_sc_hd__inv_2
X_12356_ _24842_/Q VGND VGND VPWR VPWR _12356_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24775__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15075_ _15075_/A VGND VGND VPWR VPWR _15075_/Y sky130_fd_sc_hd__inv_2
X_19952_ _23557_/Q VGND VGND VPWR VPWR _19952_/Y sky130_fd_sc_hd__inv_2
X_12287_ _25360_/Q VGND VGND VPWR VPWR _12287_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24704__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14026_ _14001_/A _13990_/C _13999_/C VGND VGND VPWR VPWR _14026_/X sky130_fd_sc_hd__or3_4
X_18903_ _11938_/A _18900_/X _18902_/X VGND VGND VPWR VPWR _24115_/D sky130_fd_sc_hd__o21a_4
X_19883_ _19883_/A VGND VGND VPWR VPWR _19883_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18834_ _16479_/Y _24148_/Q _16479_/Y _24148_/Q VGND VGND VPWR VPWR _18835_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18271__A3 _16267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_57_0_HCLK clkbuf_7_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_57_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18765_ _18692_/Y _18746_/X _18735_/X _18763_/B VGND VGND VPWR VPWR _18765_/X sky130_fd_sc_hd__a211o_4
X_15977_ _12212_/Y _15972_/X _15976_/X _15972_/X VGND VGND VPWR VPWR _24750_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15490__B1 HADDR[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17716_ _19455_/B VGND VGND VPWR VPWR _18280_/C sky130_fd_sc_hd__buf_2
X_14928_ _15058_/A VGND VGND VPWR VPWR _15251_/A sky130_fd_sc_hd__buf_2
X_18696_ _18729_/A _18728_/A _18696_/C _18695_/X VGND VGND VPWR VPWR _18696_/X sky130_fd_sc_hd__or4_4
XFILLER_224_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17647_ _17647_/A _17647_/B _17646_/Y VGND VGND VPWR VPWR _17647_/X sky130_fd_sc_hd__and3_4
XANTENNA__18693__D _18692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16896__A1_N _22564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14859_ _14859_/A _14859_/B _14859_/C _14817_/X VGND VGND VPWR VPWR _14859_/X sky130_fd_sc_hd__or4_4
XFILLER_63_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17578_ _24295_/Q VGND VGND VPWR VPWR _17578_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19317_ _18202_/B VGND VGND VPWR VPWR _19317_/Y sky130_fd_sc_hd__inv_2
X_16529_ _16527_/Y _16521_/X _16349_/X _16528_/X VGND VGND VPWR VPWR _16529_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16791__A _24445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19248_ _21386_/B _19245_/X _16885_/X _19245_/X VGND VGND VPWR VPWR _23804_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__14348__A2 _14340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16742__B1 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19179_ _23828_/Q VGND VGND VPWR VPWR _19179_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21210_ _17707_/X _21210_/B _21210_/C VGND VGND VPWR VPWR _21210_/X sky130_fd_sc_hd__and3_4
X_22190_ _22190_/A _21235_/A VGND VGND VPWR VPWR _22190_/X sky130_fd_sc_hd__or2_4
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21141_ _21135_/Y _21141_/B _21139_/X _21141_/D VGND VGND VPWR VPWR _21141_/X sky130_fd_sc_hd__and4_4
XANTENNA__19607__A _19598_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24445__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18247__B1 _15965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21072_ _21109_/A _21064_/X _21072_/C VGND VGND VPWR VPWR _21072_/X sky130_fd_sc_hd__and3_4
XANTENNA__23240__B1 _22839_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20023_ _20022_/Y _20018_/X _19977_/X _20018_/X VGND VGND VPWR VPWR _23534_/D sky130_fd_sc_hd__a2bb2o_4
X_24900_ _24900_/CLK _15617_/X HRESETn VGND VGND VPWR VPWR _24900_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24831_ _24855_/CLK _15819_/X HRESETn VGND VGND VPWR VPWR _24831_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22664__A1_N _22572_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24762_ _24762_/CLK _24762_/D HRESETn VGND VGND VPWR VPWR _24762_/Q sky130_fd_sc_hd__dfrtp_4
X_21974_ _21974_/A _20307_/X VGND VGND VPWR VPWR _21974_/X sky130_fd_sc_hd__or2_4
XFILLER_132_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23713_ _23406_/CLK _23713_/D VGND VGND VPWR VPWR _23713_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ _20921_/C _13637_/X VGND VGND VPWR VPWR _20925_/Y sky130_fd_sc_hd__nor2_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17222__B2 _17203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24693_ _24762_/CLK _16134_/X HRESETn VGND VGND VPWR VPWR _22638_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23644_ _23644_/CLK _19712_/X VGND VGND VPWR VPWR _13410_/B sky130_fd_sc_hd__dfxtp_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20856_ _24042_/Q VGND VGND VPWR VPWR _20862_/A sky130_fd_sc_hd__inv_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17797__A _16906_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13795__B1 _13521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23575_ _23575_/CLK _23575_/D VGND VGND VPWR VPWR _23575_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20787_ _13108_/C _20782_/X _20786_/Y VGND VGND VPWR VPWR _20787_/Y sky130_fd_sc_hd__a21oi_4
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25314_ _25492_/CLK _25314_/D HRESETn VGND VGND VPWR VPWR _11976_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_22_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22526_ _22525_/X VGND VGND VPWR VPWR _22686_/A sky130_fd_sc_hd__buf_2
XFILLER_194_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16733__B1 _16464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15536__B2 _15533_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22208__A _22223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25245_ _25204_/CLK _13870_/X HRESETn VGND VGND VPWR VPWR _25245_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22457_ _21587_/A _22457_/B VGND VGND VPWR VPWR _22457_/Y sky130_fd_sc_hd__nor2_4
XFILLER_155_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _12207_/A _22476_/A _12208_/X _12209_/Y VGND VGND VPWR VPWR _12214_/C sky130_fd_sc_hd__o22a_4
X_21408_ _22197_/A _21408_/B VGND VGND VPWR VPWR _21408_/X sky130_fd_sc_hd__or2_4
X_13190_ _13285_/A _23873_/Q VGND VGND VPWR VPWR _13193_/B sky130_fd_sc_hd__or2_4
X_25176_ _23884_/CLK _14303_/X HRESETn VGND VGND VPWR VPWR _25176_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22388_ _22378_/A _19831_/Y _22226_/A VGND VGND VPWR VPWR _22388_/X sky130_fd_sc_hd__o21a_4
XFILLER_163_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12141_ _12141_/A VGND VGND VPWR VPWR _12141_/Y sky130_fd_sc_hd__inv_2
X_24127_ _24133_/CLK _24127_/D HRESETn VGND VGND VPWR VPWR _18641_/A sky130_fd_sc_hd__dfrtp_4
X_21339_ _23178_/A VGND VGND VPWR VPWR _21339_/X sky130_fd_sc_hd__buf_2
XFILLER_123_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24186__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12072_ _12060_/A VGND VGND VPWR VPWR _12072_/X sky130_fd_sc_hd__buf_2
X_24058_ _24501_/CLK _20931_/Y HRESETn VGND VGND VPWR VPWR _13651_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24115__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15900_ _12776_/Y _15896_/X _15472_/X _15896_/X VGND VGND VPWR VPWR _24787_/D sky130_fd_sc_hd__a2bb2o_4
X_23009_ _24569_/Q _23075_/B _23075_/C VGND VGND VPWR VPWR _23009_/X sky130_fd_sc_hd__and3_4
X_16880_ _16880_/A VGND VGND VPWR VPWR _19827_/A sky130_fd_sc_hd__buf_2
XFILLER_103_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12900__C _12741_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15831_ _15818_/X _15829_/X _15830_/X _24824_/Q _15786_/X VGND VGND VPWR VPWR _24824_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21782__A _22228_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20060__A3 _18257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15780__A _14366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22597__B _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18550_ _18549_/X VGND VGND VPWR VPWR _24172_/D sky130_fd_sc_hd__inv_2
X_12974_ _12287_/Y _12308_/Y VGND VGND VPWR VPWR _12987_/C sky130_fd_sc_hd__or2_4
X_15762_ _11774_/A VGND VGND VPWR VPWR _15762_/X sky130_fd_sc_hd__buf_2
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21545__B1 _16917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17501_ _25530_/Q _17499_/Y _17585_/A _25546_/Q VGND VGND VPWR VPWR _17501_/X sky130_fd_sc_hd__a2bb2o_4
X_14713_ _14711_/X _14712_/X _14711_/X _14712_/X VGND VGND VPWR VPWR _14713_/X sky130_fd_sc_hd__a2bb2o_4
X_11925_ _11923_/Y _11919_/X _11924_/X _11919_/X VGND VGND VPWR VPWR _11925_/X sky130_fd_sc_hd__a2bb2o_4
X_18481_ _18481_/A _18510_/C _18481_/C _18480_/X VGND VGND VPWR VPWR _18499_/B sky130_fd_sc_hd__or4_4
XFILLER_61_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15693_ _24888_/Q _15687_/Y _15686_/B _15692_/X VGND VGND VPWR VPWR _15693_/X sky130_fd_sc_hd__o22a_4
XFILLER_205_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17432_ _17431_/Y _17429_/X _16787_/X _17429_/X VGND VGND VPWR VPWR _24327_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11856_ _11856_/A _11856_/B VGND VGND VPWR VPWR _11856_/X sky130_fd_sc_hd__and2_4
X_14644_ _17943_/A _14630_/C _14642_/X VGND VGND VPWR VPWR _25075_/D sky130_fd_sc_hd__o21a_4
XANTENNA__23298__B1 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16972__B1 _16052_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13786__B1 _13785_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14575_ _14566_/D VGND VGND VPWR VPWR _14575_/X sky130_fd_sc_hd__buf_2
X_17363_ _17366_/A _17366_/B VGND VGND VPWR VPWR _17367_/B sky130_fd_sc_hd__or2_4
XFILLER_60_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21848__B2 _22327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11787_ _11783_/Y _11778_/X _11786_/X _11778_/X VGND VGND VPWR VPWR _25522_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19102_ _19100_/Y _19096_/X _18985_/X _19101_/X VGND VGND VPWR VPWR _19102_/X sky130_fd_sc_hd__a2bb2o_4
X_16314_ _16313_/Y _16311_/X _15951_/X _16311_/X VGND VGND VPWR VPWR _16314_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13526_ _24784_/Q VGND VGND VPWR VPWR _15688_/A sky130_fd_sc_hd__inv_2
X_17294_ _17230_/X _17292_/X _17294_/C VGND VGND VPWR VPWR _24366_/D sky130_fd_sc_hd__and3_4
XANTENNA__15527__B2 _15524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19033_ _19028_/A VGND VGND VPWR VPWR _19033_/X sky130_fd_sc_hd__buf_2
X_13457_ _13462_/C _13456_/X _12160_/C _13457_/D VGND VGND VPWR VPWR _13458_/A sky130_fd_sc_hd__or4_4
X_16245_ _16239_/A VGND VGND VPWR VPWR _16245_/X sky130_fd_sc_hd__buf_2
X_12408_ _12413_/A _12406_/X _12408_/C VGND VGND VPWR VPWR _12408_/X sky130_fd_sc_hd__and3_4
X_13388_ _13388_/A _23868_/Q VGND VGND VPWR VPWR _13390_/B sky130_fd_sc_hd__or2_4
X_16176_ _14758_/B _16174_/Y _14758_/A _16174_/Y VGND VGND VPWR VPWR _16176_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12347__A2_N _24835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_20_0_HCLK clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_41_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12339_ _12339_/A _12334_/X _12336_/X _12339_/D VGND VGND VPWR VPWR _12369_/A sky130_fd_sc_hd__or4_4
X_15127_ _15127_/A _15127_/B _15127_/C _15127_/D VGND VGND VPWR VPWR _15127_/X sky130_fd_sc_hd__or4_4
XANTENNA__15955__A _15783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15058_ _15058_/A _15002_/A _15246_/C _15243_/A VGND VGND VPWR VPWR _15058_/X sky130_fd_sc_hd__or4_4
X_19935_ _21474_/B _19932_/X _19620_/X _19932_/X VGND VGND VPWR VPWR _23564_/D sky130_fd_sc_hd__a2bb2o_4
X_14009_ _14525_/A _14008_/X VGND VGND VPWR VPWR _14009_/Y sky130_fd_sc_hd__nand2_4
XFILLER_96_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19866_ _19866_/A VGND VGND VPWR VPWR _19866_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18244__A3 _16236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22788__A _16677_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18817_ _18683_/Y _18820_/B _18709_/X VGND VGND VPWR VPWR _18817_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19797_ _19795_/Y _19796_/X _19708_/X _19796_/X VGND VGND VPWR VPWR _23613_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16786__A _16786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22328__A2 _14182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19729__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18748_ _18658_/Y _18748_/B VGND VGND VPWR VPWR _18749_/A sky130_fd_sc_hd__or2_4
XFILLER_36_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_144_0_HCLK clkbuf_7_72_0_HCLK/X VGND VGND VPWR VPWR _23388_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_64_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18679_ _24137_/Q VGND VGND VPWR VPWR _18679_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20710_ _20709_/Y _20704_/Y _13116_/B VGND VGND VPWR VPWR _20710_/X sky130_fd_sc_hd__o21a_4
XFILLER_197_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21690_ _23420_/Q _22396_/B _23396_/Q _22397_/B VGND VGND VPWR VPWR _21690_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16963__B1 _16006_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20641_ _15456_/Y _20638_/X _20629_/X _20640_/X VGND VGND VPWR VPWR _20641_/X sky130_fd_sc_hd__a211o_4
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23360_ _23344_/X VGND VGND VPWR VPWR IRQ[16] sky130_fd_sc_hd__buf_2
XFILLER_149_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17410__A _17410_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20572_ _18886_/X VGND VGND VPWR VPWR _20572_/X sky130_fd_sc_hd__buf_2
XANTENNA__24697__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22311_ _14917_/A _21325_/X _15663_/A _22310_/X VGND VGND VPWR VPWR _22311_/X sky130_fd_sc_hd__a211o_4
XFILLER_164_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23291_ _16639_/Y _23291_/B VGND VGND VPWR VPWR _23291_/X sky130_fd_sc_hd__and2_4
XANTENNA__24626__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25030_ _25028_/CLK _25030_/D HRESETn VGND VGND VPWR VPWR _25030_/Q sky130_fd_sc_hd__dfrtp_4
X_22242_ _22257_/A _22237_/X _22241_/X VGND VGND VPWR VPWR _22242_/X sky130_fd_sc_hd__or3_4
XFILLER_180_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15865__A _15861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22173_ _14465_/Y _14245_/A _25108_/Q _22181_/B VGND VGND VPWR VPWR _22173_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21124_ _21124_/A _21124_/B VGND VGND VPWR VPWR _21130_/B sky130_fd_sc_hd__or2_4
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21055_ _22189_/A VGND VGND VPWR VPWR _21055_/X sky130_fd_sc_hd__buf_2
XFILLER_219_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20006_ _21471_/B _20003_/X _19984_/X _20003_/X VGND VGND VPWR VPWR _20006_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25485__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_40_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_40_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_24814_ _25373_/CLK _24814_/D HRESETn VGND VGND VPWR VPWR _12770_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21957_ _21939_/X _21954_/X _21956_/X VGND VGND VPWR VPWR _21957_/X sky130_fd_sc_hd__a21o_4
X_24745_ _24744_/CLK _24745_/D HRESETn VGND VGND VPWR VPWR _24745_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__23025__C _23024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A VGND VGND VPWR VPWR _11710_/Y sky130_fd_sc_hd__inv_2
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20906_/Y _20903_/X _20907_/X VGND VGND VPWR VPWR _20908_/X sky130_fd_sc_hd__o21a_4
XFILLER_188_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12690_ _12584_/X _12717_/A _12716_/A _12716_/B VGND VGND VPWR VPWR _12690_/X sky130_fd_sc_hd__or4_4
X_24676_ _24678_/CLK _24676_/D HRESETn VGND VGND VPWR VPWR _23248_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _22083_/A _21888_/B VGND VGND VPWR VPWR _21890_/B sky130_fd_sc_hd__or2_4
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23627_ _23627_/CLK _23627_/D VGND VGND VPWR VPWR _19758_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _20838_/Y _13640_/X _13642_/X VGND VGND VPWR VPWR _20839_/X sky130_fd_sc_hd__o21a_4
XFILLER_168_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14344_/A _14359_/X _12074_/A _14349_/A VGND VGND VPWR VPWR _14360_/X sky130_fd_sc_hd__o22a_4
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23558_ _23555_/CLK _23558_/D VGND VGND VPWR VPWR _23558_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13438_/A _13311_/B VGND VGND VPWR VPWR _13311_/X sky130_fd_sc_hd__or2_4
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22509_ _16244_/Y _16180_/X _15107_/Y _16366_/B VGND VGND VPWR VPWR _22509_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14291_ _14288_/Y VGND VGND VPWR VPWR _14291_/X sky130_fd_sc_hd__buf_2
XANTENNA__24367__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23489_ _23497_/CLK _20141_/X VGND VGND VPWR VPWR _20140_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13242_ _13353_/A _13230_/X _13241_/X VGND VGND VPWR VPWR _13242_/X sky130_fd_sc_hd__and3_4
X_16030_ _16029_/Y _16025_/X _15953_/X _16025_/X VGND VGND VPWR VPWR _16030_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_182_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14193__B1 _13826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25228_ _25230_/CLK _25228_/D HRESETn VGND VGND VPWR VPWR _14005_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__21777__A _22380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11696__A1_N _11694_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13173_ _13169_/X _13172_/X _13150_/X VGND VGND VPWR VPWR _13173_/X sky130_fd_sc_hd__o21a_4
X_25159_ _23938_/CLK _14352_/X HRESETn VGND VGND VPWR VPWR _25159_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12124_ _25472_/Q _24101_/Q _25472_/Q _24101_/Q VGND VGND VPWR VPWR _12133_/B sky130_fd_sc_hd__a2bb2o_4
X_17981_ _17981_/A _17981_/B _17981_/C VGND VGND VPWR VPWR _17981_/X sky130_fd_sc_hd__and3_4
XFILLER_124_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19720_ _13235_/B VGND VGND VPWR VPWR _19720_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12055_ _12081_/A _12083_/A VGND VGND VPWR VPWR _21571_/A sky130_fd_sc_hd__or2_4
X_16932_ _16120_/Y _16921_/A _22980_/A _17817_/A VGND VGND VPWR VPWR _16934_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17990__A _18095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19651_ _19650_/Y VGND VGND VPWR VPWR _19651_/X sky130_fd_sc_hd__buf_2
XFILLER_78_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16863_ _16863_/A VGND VGND VPWR VPWR _16863_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23931__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18602_ _16538_/Y _18703_/A _16538_/Y _24157_/Q VGND VGND VPWR VPWR _18607_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15814_ _15810_/X _15813_/X _16226_/A _24835_/Q _15811_/X VGND VGND VPWR VPWR _15814_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19582_ _19580_/Y _19576_/X _19395_/X _19581_/X VGND VGND VPWR VPWR _19582_/X sky130_fd_sc_hd__a2bb2o_4
X_16794_ _16793_/X VGND VGND VPWR VPWR _16794_/X sky130_fd_sc_hd__buf_2
XFILLER_237_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23216__B _22658_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18533_ _18465_/Y _18524_/X VGND VGND VPWR VPWR _18533_/X sky130_fd_sc_hd__or2_4
XFILLER_18_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15745_ _15724_/A VGND VGND VPWR VPWR _15745_/X sky130_fd_sc_hd__buf_2
XFILLER_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12957_ _12956_/X VGND VGND VPWR VPWR _12957_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_217_0_HCLK clkbuf_7_108_0_HCLK/X VGND VGND VPWR VPWR _24463_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11908_ _11905_/Y _11898_/X _11906_/X _11907_/X VGND VGND VPWR VPWR _11908_/X sky130_fd_sc_hd__a2bb2o_4
X_18464_ _24173_/Q VGND VGND VPWR VPWR _18466_/C sky130_fd_sc_hd__inv_2
X_15676_ _24888_/Q VGND VGND VPWR VPWR _15676_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18862__A1_N _16507_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12888_ _12888_/A VGND VGND VPWR VPWR _25390_/D sky130_fd_sc_hd__inv_2
XPHY_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _14400_/A VGND VGND VPWR VPWR _17415_/X sky130_fd_sc_hd__buf_2
XFILLER_61_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14627_ _13525_/Y _13588_/X _13621_/Y VGND VGND VPWR VPWR _14630_/C sky130_fd_sc_hd__o21a_4
X_11839_ _13676_/A _22517_/A _13676_/A _22517_/A VGND VGND VPWR VPWR _11846_/B sky130_fd_sc_hd__a2bb2o_4
X_18395_ _18395_/A VGND VGND VPWR VPWR _18471_/D sky130_fd_sc_hd__inv_2
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14420__B2 _14408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _17346_/A _17366_/A _17346_/C _17346_/D VGND VGND VPWR VPWR _17352_/C sky130_fd_sc_hd__or4_4
X_14558_ _14557_/X VGND VGND VPWR VPWR _14559_/B sky130_fd_sc_hd__inv_2
XANTENNA__24790__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13509_ _13509_/A _13509_/B VGND VGND VPWR VPWR _13509_/X sky130_fd_sc_hd__or2_4
XFILLER_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17277_ _17231_/X _17265_/X _17276_/X _17273_/B VGND VGND VPWR VPWR _17277_/X sky130_fd_sc_hd__a211o_4
XFILLER_158_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14489_ _23958_/Q VGND VGND VPWR VPWR _14490_/C sky130_fd_sc_hd__inv_2
X_19016_ _19015_/Y _19011_/X _18965_/X _19011_/X VGND VGND VPWR VPWR _23886_/D sky130_fd_sc_hd__a2bb2o_4
X_16228_ _22705_/A VGND VGND VPWR VPWR _16228_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24037__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16159_ _21521_/A VGND VGND VPWR VPWR _16159_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22549__A2 _22432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11718__A HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19918_ _23570_/Q VGND VGND VPWR VPWR _19918_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19849_ _23596_/Q VGND VGND VPWR VPWR _19849_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18622__B1 _16600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12224__A2_N _24760_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_27_0_HCLK clkbuf_6_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_55_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_22860_ _22769_/A _22859_/X VGND VGND VPWR VPWR _22860_/X sky130_fd_sc_hd__and2_4
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21811_ _22021_/A _21811_/B _21811_/C VGND VGND VPWR VPWR _21811_/X sky130_fd_sc_hd__and3_4
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22791_ _15593_/Y _22989_/B VGND VGND VPWR VPWR _22791_/X sky130_fd_sc_hd__and2_4
XANTENNA__22182__B1 _14215_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24530_ _24540_/CLK _24530_/D HRESETn VGND VGND VPWR VPWR _16582_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_225_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21742_ _16613_/Y _21581_/X _21582_/A _21741_/X VGND VGND VPWR VPWR _21742_/X sky130_fd_sc_hd__o22a_4
XANTENNA__19620__A _19620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24878__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24461_ _24462_/CLK _24461_/D HRESETn VGND VGND VPWR VPWR _24461_/Q sky130_fd_sc_hd__dfrtp_4
X_21673_ _21656_/A _21671_/X _21673_/C VGND VGND VPWR VPWR _21673_/X sky130_fd_sc_hd__and3_4
XFILLER_212_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24807__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14764__A _14764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23412_ _24302_/CLK _20342_/X VGND VGND VPWR VPWR _20340_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20624_ _23977_/Q _17385_/X VGND VGND VPWR VPWR _20624_/Y sky130_fd_sc_hd__nand2_4
X_24392_ _24315_/CLK _17101_/X HRESETn VGND VGND VPWR VPWR _24392_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23343_ _25274_/Q _21970_/X _23341_/Y _23342_/Y VGND VGND VPWR VPWR _23343_/X sky130_fd_sc_hd__a211o_4
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20555_ _20555_/A VGND VGND VPWR VPWR _20555_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24460__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23029__A3 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12284__A _24826_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21597__A _21597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23274_ _23251_/X _23274_/B _23266_/X _23273_/X VGND VGND VPWR VPWR HRDATA[29] sky130_fd_sc_hd__or4_4
XANTENNA__15911__A1 _14764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20486_ _23998_/Q VGND VGND VPWR VPWR _20486_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25013_ _24967_/CLK _15269_/X HRESETn VGND VGND VPWR VPWR _25013_/Q sky130_fd_sc_hd__dfrtp_4
X_22225_ _22225_/A _22225_/B VGND VGND VPWR VPWR _22225_/X sky130_fd_sc_hd__or2_4
XANTENNA__19067__A _19360_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22156_ _21114_/X _22148_/X _22152_/X _22155_/X VGND VGND VPWR VPWR _22157_/B sky130_fd_sc_hd__a211o_4
XFILLER_161_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_7_109_0_HCLK clkbuf_6_54_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_219_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21107_ _21013_/B _21048_/Y VGND VGND VPWR VPWR _21107_/X sky130_fd_sc_hd__and2_4
XFILLER_248_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22087_ _21896_/X _22083_/X _22084_/X _22085_/X _22086_/X VGND VGND VPWR VPWR _22087_/X
+ sky130_fd_sc_hd__a32o_4
X_21038_ _11676_/B _14462_/A VGND VGND VPWR VPWR _21038_/X sky130_fd_sc_hd__or2_4
XANTENNA__17416__B2 _17414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22221__A _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14939__A _24415_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22960__A2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13860_ _23995_/Q VGND VGND VPWR VPWR _13860_/X sky130_fd_sc_hd__buf_2
XFILLER_247_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14990__A2_N _24474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12811_ _12744_/Y _24811_/Q _25388_/Q _12810_/Y VGND VGND VPWR VPWR _12811_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13791_ _15472_/A VGND VGND VPWR VPWR _13791_/X sky130_fd_sc_hd__buf_2
X_22989_ _15580_/Y _22989_/B VGND VGND VPWR VPWR _22989_/X sky130_fd_sc_hd__and2_4
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15530_ _15530_/A VGND VGND VPWR VPWR _15530_/X sky130_fd_sc_hd__buf_2
X_12742_ _12741_/X _24801_/Q _12741_/X _24801_/Q VGND VGND VPWR VPWR _12742_/X sky130_fd_sc_hd__a2bb2o_4
X_24728_ _24357_/CLK _24728_/D HRESETn VGND VGND VPWR VPWR _16042_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16927__B1 _16133_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18392__A2 _17268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_190_0_HCLK clkbuf_7_95_0_HCLK/X VGND VGND VPWR VPWR _25100_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_43_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12673_ _12664_/C _12663_/X VGND VGND VPWR VPWR _12673_/Y sky130_fd_sc_hd__nand2_4
X_15461_ _15460_/Y _15458_/X _14403_/X _15458_/X VGND VGND VPWR VPWR _15461_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24659_ _24592_/CLK _24659_/D HRESETn VGND VGND VPWR VPWR _24659_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24548__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17200_/A VGND VGND VPWR VPWR _17200_/Y sky130_fd_sc_hd__inv_2
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_8_47_0_HCLK clkbuf_8_47_0_HCLK/A VGND VGND VPWR VPWR _23706_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _25141_/Q VGND VGND VPWR VPWR _14412_/Y sky130_fd_sc_hd__inv_2
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18180_ _18052_/A _18180_/B _18179_/X VGND VGND VPWR VPWR _18180_/X sky130_fd_sc_hd__or3_4
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _15068_/Y _15394_/B _15391_/Y VGND VGND VPWR VPWR _15392_/X sky130_fd_sc_hd__o21a_4
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ _17035_/A _17140_/B VGND VGND VPWR VPWR _17131_/X sky130_fd_sc_hd__or2_4
XFILLER_128_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14343_ _14349_/A VGND VGND VPWR VPWR _14344_/A sky130_fd_sc_hd__inv_2
XANTENNA__17985__A _17999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14274_ _23442_/Q _14269_/X _14273_/A _25184_/Q _14273_/Y VGND VGND VPWR VPWR _14274_/X
+ sky130_fd_sc_hd__a32o_4
X_17062_ _17062_/A _17333_/A VGND VGND VPWR VPWR _17062_/X sky130_fd_sc_hd__and2_4
XANTENNA__24130__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15902__B2 _15861_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20239__B1 _19759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13225_ _13225_/A VGND VGND VPWR VPWR _13374_/A sky130_fd_sc_hd__buf_2
X_16013_ _16011_/Y _16007_/X _15939_/X _16012_/X VGND VGND VPWR VPWR _16013_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13156_ _13169_/A VGND VGND VPWR VPWR _13179_/A sky130_fd_sc_hd__buf_2
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12107_ _12102_/A VGND VGND VPWR VPWR _12107_/X sky130_fd_sc_hd__buf_2
XFILLER_239_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25336__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13087_ _13087_/A VGND VGND VPWR VPWR _13091_/C sky130_fd_sc_hd__buf_2
X_17964_ _17966_/A VGND VGND VPWR VPWR _18024_/A sky130_fd_sc_hd__inv_2
XFILLER_111_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19703_ _19701_/Y _19699_/X _19702_/X _19699_/X VGND VGND VPWR VPWR _23647_/D sky130_fd_sc_hd__a2bb2o_4
X_12038_ _14177_/A _12038_/B VGND VGND VPWR VPWR _12039_/D sky130_fd_sc_hd__or2_4
X_16915_ _16915_/A VGND VGND VPWR VPWR _16915_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17895_ _17893_/Y _17906_/B _17893_/A _17894_/Y VGND VGND VPWR VPWR _17907_/A sky130_fd_sc_hd__o22a_4
X_19634_ _19641_/A VGND VGND VPWR VPWR _19634_/X sky130_fd_sc_hd__buf_2
X_16846_ _16844_/Y _16841_/X _16778_/X _16845_/X VGND VGND VPWR VPWR _24418_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19565_ _21495_/B _19562_/X _11927_/X _19562_/X VGND VGND VPWR VPWR _19565_/X sky130_fd_sc_hd__a2bb2o_4
X_16777_ HWDATA[4] VGND VGND VPWR VPWR _18942_/A sky130_fd_sc_hd__buf_2
X_13989_ _25240_/Q VGND VGND VPWR VPWR _13989_/X sky130_fd_sc_hd__buf_2
XANTENNA__22164__B1 _21339_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22703__A2 _21336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18516_ _18497_/A _18516_/B _18516_/C VGND VGND VPWR VPWR _18516_/X sky130_fd_sc_hd__and3_4
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18907__B2 _11794_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15728_ _15713_/X VGND VGND VPWR VPWR _15728_/X sky130_fd_sc_hd__buf_2
X_19496_ _23716_/Q VGND VGND VPWR VPWR _19496_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24971__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12088__B _12086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18447_ _16259_/Y _24161_/Q _21335_/A _18561_/C VGND VGND VPWR VPWR _18451_/A sky130_fd_sc_hd__a2bb2o_4
X_15659_ _15666_/A VGND VGND VPWR VPWR _15660_/A sky130_fd_sc_hd__inv_2
XANTENNA__24289__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24900__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18056__A _18056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18378_ _24196_/Q VGND VGND VPWR VPWR _18378_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22467__B2 _22279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24218__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17329_ _17329_/A _17329_/B VGND VGND VPWR VPWR _17330_/C sky130_fd_sc_hd__or2_4
X_20340_ _20340_/A VGND VGND VPWR VPWR _20340_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20271_ _20271_/A VGND VGND VPWR VPWR _20271_/Y sky130_fd_sc_hd__inv_2
X_22010_ _22014_/A _22010_/B VGND VGND VPWR VPWR _22010_/X sky130_fd_sc_hd__or2_4
XFILLER_89_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25077__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21864__B _21864_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25006__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15672__A3 _15643_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23961_ _24980_/CLK _23961_/D HRESETn VGND VGND VPWR VPWR _21012_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20402__B1 _20061_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22912_ _22774_/X _22907_/Y _22868_/X _22911_/X VGND VGND VPWR VPWR _22912_/X sky130_fd_sc_hd__a2bb2o_4
X_23892_ _23887_/CLK _18996_/X VGND VGND VPWR VPWR _23892_/Q sky130_fd_sc_hd__dfxtp_4
X_22843_ _14936_/A _22838_/X _22839_/X _22842_/X VGND VGND VPWR VPWR _22844_/C sky130_fd_sc_hd__a211o_4
XFILLER_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22774_ _22429_/X VGND VGND VPWR VPWR _22774_/X sky130_fd_sc_hd__buf_2
XFILLER_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20496__A _20496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_200_0_HCLK clkbuf_8_201_0_HCLK/A VGND VGND VPWR VPWR _24650_/CLK sky130_fd_sc_hd__clkbuf_1
X_21725_ _21725_/A VGND VGND VPWR VPWR _21725_/Y sky130_fd_sc_hd__inv_2
X_24513_ _24679_/CLK _24513_/D HRESETn VGND VGND VPWR VPWR _24513_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25493_ _25474_/CLK _25493_/D HRESETn VGND VGND VPWR VPWR _12019_/A sky130_fd_sc_hd__dfrtp_4
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24641__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11911__A _19606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_6_0_HCLK clkbuf_8_7_0_HCLK/A VGND VGND VPWR VPWR _23525_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_169_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21656_ _21656_/A _21654_/X _21656_/C VGND VGND VPWR VPWR _21656_/X sky130_fd_sc_hd__and3_4
X_24444_ _24477_/CLK _16797_/X HRESETn VGND VGND VPWR VPWR _16796_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12731__A2_N _24796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20607_ _20601_/A _20604_/Y _20605_/Y _14484_/X _20606_/X VGND VGND VPWR VPWR _20607_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_137_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24375_ _24725_/CLK _17157_/X HRESETn VGND VGND VPWR VPWR _24375_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_184_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21587_ _21587_/A _21587_/B VGND VGND VPWR VPWR _21601_/C sky130_fd_sc_hd__nor2_4
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23326_ _22686_/A _23326_/B VGND VGND VPWR VPWR _23326_/Y sky130_fd_sc_hd__nor2_4
XFILLER_181_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20538_ _20437_/C _20444_/B _20507_/X VGND VGND VPWR VPWR _24083_/D sky130_fd_sc_hd__a21o_4
XFILLER_181_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21120__A _21290_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23257_ _12204_/Y _22499_/X _23256_/X VGND VGND VPWR VPWR _23257_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_137_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20469_ _20469_/A _20453_/C _20466_/X VGND VGND VPWR VPWR _20469_/X sky130_fd_sc_hd__and3_4
XANTENNA__16214__A _22927_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13010_ _12285_/A _13009_/Y VGND VGND VPWR VPWR _13010_/X sky130_fd_sc_hd__or2_4
X_22208_ _22223_/A _22208_/B _22207_/X VGND VGND VPWR VPWR _22208_/X sky130_fd_sc_hd__and3_4
XFILLER_152_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15043__A2_N _16765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23188_ _22971_/X _23187_/X _22973_/X _12515_/A _22974_/X VGND VGND VPWR VPWR _23189_/B
+ sky130_fd_sc_hd__a32o_4
X_22139_ _22716_/A _22131_/X _22135_/X _22138_/X VGND VGND VPWR VPWR _22140_/B sky130_fd_sc_hd__a211o_4
XFILLER_0_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14961_ _25012_/Q VGND VGND VPWR VPWR _15244_/A sky130_fd_sc_hd__inv_2
XFILLER_181_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16700_ _16699_/Y _16697_/X _16518_/X _16697_/X VGND VGND VPWR VPWR _24486_/D sky130_fd_sc_hd__a2bb2o_4
X_13912_ _13931_/A _13931_/B _13930_/A _13932_/C VGND VGND VPWR VPWR _13912_/X sky130_fd_sc_hd__a211o_4
X_17680_ _17682_/A _17670_/X _17680_/C VGND VGND VPWR VPWR _17680_/X sky130_fd_sc_hd__and3_4
X_14892_ _14892_/A VGND VGND VPWR VPWR _15062_/D sky130_fd_sc_hd__inv_2
XFILLER_236_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16631_ _16631_/A _16632_/B VGND VGND VPWR VPWR _16631_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_10_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_21_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_13843_ _25254_/Q _13842_/B _13841_/X _13842_/Y VGND VGND VPWR VPWR _13843_/X sky130_fd_sc_hd__a211o_4
XANTENNA__24729__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19350_ _19350_/A VGND VGND VPWR VPWR _19350_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16562_ _24538_/Q VGND VGND VPWR VPWR _16562_/Y sky130_fd_sc_hd__inv_2
X_13774_ _25275_/Q VGND VGND VPWR VPWR _13774_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18301_ _18301_/A VGND VGND VPWR VPWR _18301_/X sky130_fd_sc_hd__buf_2
X_15513_ _15510_/Y _15506_/X HADDR[12] _15512_/X VGND VGND VPWR VPWR _15513_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12725_ _12721_/B _12725_/B _12722_/C VGND VGND VPWR VPWR _25402_/D sky130_fd_sc_hd__and3_4
X_19281_ _19281_/A VGND VGND VPWR VPWR _19281_/Y sky130_fd_sc_hd__inv_2
X_16493_ _16492_/Y _16488_/X _16402_/X _16488_/X VGND VGND VPWR VPWR _24564_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24382__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18232_ _17446_/X VGND VGND VPWR VPWR _20369_/A sky130_fd_sc_hd__buf_2
XANTENNA__14387__B1 _14262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15444_ _15432_/A VGND VGND VPWR VPWR _15444_/X sky130_fd_sc_hd__buf_2
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24311__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12656_ _12656_/A VGND VGND VPWR VPWR _12657_/B sky130_fd_sc_hd__inv_2
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14926__A2 _24443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18163_ _18099_/A _18163_/B _18163_/C VGND VGND VPWR VPWR _18164_/C sky130_fd_sc_hd__or3_4
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12587_ _12587_/A _12587_/B _12577_/X _12586_/X VGND VGND VPWR VPWR _12588_/B sky130_fd_sc_hd__or4_4
X_15375_ _15123_/Y _15375_/B VGND VGND VPWR VPWR _15376_/A sky130_fd_sc_hd__or2_4
XFILLER_8_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12241__A1_N _12240_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17114_ _17113_/X VGND VGND VPWR VPWR _17114_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14326_ _14326_/A VGND VGND VPWR VPWR _14329_/A sky130_fd_sc_hd__inv_2
X_18094_ _18094_/A _18094_/B _18093_/X VGND VGND VPWR VPWR _18099_/B sky130_fd_sc_hd__and3_4
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21030__A _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17045_ _17045_/A _17006_/Y _17026_/X _17045_/D VGND VGND VPWR VPWR _17045_/X sky130_fd_sc_hd__or4_4
XFILLER_99_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25517__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14257_ _14256_/Y _14252_/X _13788_/X _14252_/X VGND VGND VPWR VPWR _14257_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16124__A _16124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12652__A _12680_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14882__A2_N _24425_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13208_ _13392_/A _13208_/B VGND VGND VPWR VPWR _13209_/C sky130_fd_sc_hd__or2_4
X_14188_ _14187_/B _14185_/X _14189_/A VGND VGND VPWR VPWR _14188_/X sky130_fd_sc_hd__a21o_4
XFILLER_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13139_ _13249_/A VGND VGND VPWR VPWR _13421_/A sky130_fd_sc_hd__buf_2
XFILLER_97_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18996_ _18995_/Y _18993_/X _18951_/X _18993_/X VGND VGND VPWR VPWR _18996_/X sky130_fd_sc_hd__a2bb2o_4
X_17947_ _17947_/A _17947_/B _17947_/C VGND VGND VPWR VPWR _17947_/X sky130_fd_sc_hd__or3_4
XFILLER_227_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17878_ _17748_/Y _17852_/B _17793_/A _17876_/B VGND VGND VPWR VPWR _17878_/X sky130_fd_sc_hd__a211o_4
XANTENNA__22796__A _23328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16829_ _24427_/Q VGND VGND VPWR VPWR _16829_/Y sky130_fd_sc_hd__inv_2
X_19617_ _19617_/A VGND VGND VPWR VPWR _19617_/X sky130_fd_sc_hd__buf_2
XFILLER_93_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19548_ _19597_/A _19939_/B _19479_/X VGND VGND VPWR VPWR _19548_/X sky130_fd_sc_hd__or3_4
XFILLER_213_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19479_ _17711_/Y _18283_/X _18280_/C VGND VGND VPWR VPWR _19479_/X sky130_fd_sc_hd__or3_4
XFILLER_62_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12827__A _12967_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21510_ _21510_/A VGND VGND VPWR VPWR _21510_/X sky130_fd_sc_hd__buf_2
XFILLER_167_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14378__B1 _13829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22490_ _21127_/X VGND VGND VPWR VPWR _22490_/X sky130_fd_sc_hd__buf_2
XANTENNA__24052__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_30_0_HCLK clkbuf_8_31_0_HCLK/A VGND VGND VPWR VPWR _24305_/CLK sky130_fd_sc_hd__clkbuf_1
X_21441_ _21309_/A VGND VGND VPWR VPWR _21441_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_93_0_HCLK clkbuf_7_46_0_HCLK/X VGND VGND VPWR VPWR _25344_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24160_ _24325_/CLK _18593_/X HRESETn VGND VGND VPWR VPWR _18420_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_181_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17867__A1 _17849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21372_ _21372_/A _21372_/B _21369_/X _21372_/D VGND VGND VPWR VPWR _21372_/X sky130_fd_sc_hd__and4_4
XFILLER_147_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23111_ _23110_/X VGND VGND VPWR VPWR _23111_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15878__B1 _11721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20323_ _20322_/Y _20316_/X _11788_/X _20315_/Y VGND VGND VPWR VPWR _23419_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24091_ _25308_/CLK _24091_/D HRESETn VGND VGND VPWR VPWR _11977_/A sky130_fd_sc_hd__dfrtp_4
X_23042_ _22971_/X _23041_/X _22973_/X _24878_/Q _22974_/X VGND VGND VPWR VPWR _23043_/B
+ sky130_fd_sc_hd__a32o_4
X_20254_ _20254_/A VGND VGND VPWR VPWR _21633_/B sky130_fd_sc_hd__inv_2
XFILLER_115_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22612__B2 _22611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20185_ _20180_/A VGND VGND VPWR VPWR _20185_/X sky130_fd_sc_hd__buf_2
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24993_ _24597_/CLK _24993_/D HRESETn VGND VGND VPWR VPWR _15132_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_229_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11906__A _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23944_ _25140_/CLK _23944_/D HRESETn VGND VGND VPWR VPWR _23944_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24893__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23875_ _23875_/CLK _23875_/D VGND VGND VPWR VPWR _23875_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24822__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15802__B1 _11695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22826_ _21447_/X VGND VGND VPWR VPWR _22826_/X sky130_fd_sc_hd__buf_2
XANTENNA__22856__D _22856_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23340__A2 _25070_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25545_ _25538_/CLK _11686_/X HRESETn VGND VGND VPWR VPWR _11650_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_197_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22757_ _21592_/A _22755_/X _22111_/X _22756_/X VGND VGND VPWR VPWR _22758_/B sky130_fd_sc_hd__o22a_4
XFILLER_53_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16209__A _22996_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12737__A _12878_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12510_ _12664_/C _24871_/Q _12509_/A _24871_/Q VGND VGND VPWR VPWR _12519_/A sky130_fd_sc_hd__a2bb2o_4
X_13490_ _13490_/A VGND VGND VPWR VPWR _13490_/Y sky130_fd_sc_hd__inv_2
X_21708_ _21080_/X VGND VGND VPWR VPWR _21708_/X sky130_fd_sc_hd__buf_2
X_22688_ _22665_/X _22670_/Y _22687_/X VGND VGND VPWR VPWR HRDATA[13] sky130_fd_sc_hd__a21o_4
X_25476_ _24159_/CLK _12096_/X HRESETn VGND VGND VPWR VPWR _12094_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_212_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12456__B _12370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12441_ _12443_/B VGND VGND VPWR VPWR _12442_/B sky130_fd_sc_hd__inv_2
XFILLER_201_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21639_ _21635_/X _21638_/X _14744_/X VGND VGND VPWR VPWR _21639_/X sky130_fd_sc_hd__o21a_4
X_24427_ _24427_/CLK _16830_/X HRESETn VGND VGND VPWR VPWR _24427_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18646__A1_N _16584_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12372_ _12379_/A _12494_/A VGND VGND VPWR VPWR _12385_/B sky130_fd_sc_hd__or2_4
X_15160_ _15160_/A _15311_/B VGND VGND VPWR VPWR _15161_/D sky130_fd_sc_hd__or2_4
XFILLER_176_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24358_ _24357_/CLK _24358_/D HRESETn VGND VGND VPWR VPWR _17200_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22851__B2 _21051_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_1_0_HCLK clkbuf_5_1_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_3_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15869__B1 _11688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14111_ _23956_/Q VGND VGND VPWR VPWR _14111_/X sky130_fd_sc_hd__buf_2
X_15091_ _15091_/A VGND VGND VPWR VPWR _15091_/Y sky130_fd_sc_hd__inv_2
X_23309_ _23277_/A _23308_/X VGND VGND VPWR VPWR _23309_/X sky130_fd_sc_hd__and2_4
XFILLER_165_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24289_ _25444_/CLK _17772_/X HRESETn VGND VGND VPWR VPWR _23320_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14042_ _14001_/A _14038_/B _13999_/C VGND VGND VPWR VPWR _14042_/X sky130_fd_sc_hd__or3_4
XFILLER_69_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15884__A3 _16229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18850_ _16492_/A _18755_/B _16510_/Y _24136_/Q VGND VGND VPWR VPWR _18850_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17801_ _17790_/A _17801_/B _17801_/C VGND VGND VPWR VPWR _17801_/X sky130_fd_sc_hd__and3_4
X_18781_ _18780_/X VGND VGND VPWR VPWR _24138_/D sky130_fd_sc_hd__inv_2
X_15993_ _15993_/A VGND VGND VPWR VPWR _15993_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14399__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22186__A2_N _21849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17732_ _24219_/Q VGND VGND VPWR VPWR _17732_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14944_ _25022_/Q VGND VGND VPWR VPWR _14944_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16046__B1 _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17663_ _17663_/A VGND VGND VPWR VPWR _17663_/Y sky130_fd_sc_hd__inv_2
X_14875_ _14859_/C _14817_/X VGND VGND VPWR VPWR _14875_/Y sky130_fd_sc_hd__nand2_4
XFILLER_235_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24563__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19402_ _23749_/Q VGND VGND VPWR VPWR _19402_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16614_ _16613_/Y _16611_/X _16353_/X _16611_/X VGND VGND VPWR VPWR _24518_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_211_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13826_ _13826_/A VGND VGND VPWR VPWR _13826_/X sky130_fd_sc_hd__buf_2
X_17594_ _17587_/A _17586_/X _17589_/B _17593_/X VGND VGND VPWR VPWR _17595_/A sky130_fd_sc_hd__a211o_4
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19333_ _23773_/Q VGND VGND VPWR VPWR _19333_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21025__A _21024_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16545_ _16544_/Y _16542_/X _16373_/X _16542_/X VGND VGND VPWR VPWR _16545_/X sky130_fd_sc_hd__a2bb2o_4
X_13757_ _25276_/Q VGND VGND VPWR VPWR _13757_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17546__B1 _11710_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16939__A2_N _24284_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12708_ _12693_/A _12692_/X VGND VGND VPWR VPWR _12708_/Y sky130_fd_sc_hd__nand2_4
X_19264_ _21759_/B _19259_/X _16878_/X _19259_/X VGND VGND VPWR VPWR _23798_/D sky130_fd_sc_hd__a2bb2o_4
X_16476_ _16474_/Y _16470_/X _16386_/X _16475_/X VGND VGND VPWR VPWR _16476_/X sky130_fd_sc_hd__a2bb2o_4
X_13688_ _13687_/X VGND VGND VPWR VPWR _13688_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18215_ _18151_/A _23875_/Q VGND VGND VPWR VPWR _18215_/X sky130_fd_sc_hd__or2_4
XANTENNA__22124__A2_N _21849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15427_ _15426_/X VGND VGND VPWR VPWR _15427_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_17_0_HCLK clkbuf_6_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_35_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_12639_ _12608_/A _12638_/X VGND VGND VPWR VPWR _12639_/X sky130_fd_sc_hd__or2_4
X_19195_ _19193_/Y _19191_/X _19194_/X _19191_/X VGND VGND VPWR VPWR _19195_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23095__B2 _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18146_ _18146_/A _23901_/Q VGND VGND VPWR VPWR _18147_/C sky130_fd_sc_hd__or2_4
X_15358_ _15291_/A _15357_/X _15334_/X VGND VGND VPWR VPWR _15358_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_8_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14309_ _14295_/A _14308_/X _13475_/A _14300_/X VGND VGND VPWR VPWR _25173_/D sky130_fd_sc_hd__o22a_4
XFILLER_144_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25351__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18077_ _18054_/A VGND VGND VPWR VPWR _18146_/A sky130_fd_sc_hd__buf_2
X_15289_ _15075_/Y _15333_/A VGND VGND VPWR VPWR _15302_/C sky130_fd_sc_hd__or2_4
XFILLER_116_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23055__A1_N _17234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17028_ _24388_/Q VGND VGND VPWR VPWR _17030_/C sky130_fd_sc_hd__inv_2
XFILLER_236_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18979_ _18007_/B VGND VGND VPWR VPWR _18979_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11726__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21990_ _21841_/X _21867_/X _21882_/X _21990_/D VGND VGND VPWR VPWR HRDATA[4] sky130_fd_sc_hd__or4_4
X_20941_ _20941_/A _20941_/B VGND VGND VPWR VPWR _20941_/X sky130_fd_sc_hd__or2_4
XPHY_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20872_ _24045_/Q _13647_/B _20871_/Y VGND VGND VPWR VPWR _20872_/Y sky130_fd_sc_hd__a21oi_4
X_23660_ _24209_/CLK _19667_/X VGND VGND VPWR VPWR _19666_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__24233__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23322__A2 _21077_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22611_ _12830_/A _22572_/X _22610_/X VGND VGND VPWR VPWR _22611_/X sky130_fd_sc_hd__o21a_4
XFILLER_81_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20477__C _20477_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23591_ _23559_/CLK _19865_/X VGND VGND VPWR VPWR _19864_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_241_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17537__B1 _25541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16029__A _24733_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22542_ _21284_/X _22540_/X _21956_/X _22541_/X VGND VGND VPWR VPWR _22542_/X sky130_fd_sc_hd__o22a_4
X_25330_ _23456_/CLK _25330_/D HRESETn VGND VGND VPWR VPWR _25330_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_222_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22473_ _22443_/X _22449_/X _22457_/Y _22472_/X VGND VGND VPWR VPWR HRDATA[8] sky130_fd_sc_hd__a211o_4
X_25261_ _25089_/CLK _13827_/X HRESETn VGND VGND VPWR VPWR _13538_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21424_ _22451_/A VGND VGND VPWR VPWR _21424_/X sky130_fd_sc_hd__buf_2
X_24212_ _23678_/CLK _18312_/Y HRESETn VGND VGND VPWR VPWR _24212_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21097__B1 _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25192_ _25230_/CLK _14248_/X HRESETn VGND VGND VPWR VPWR _25192_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24143_ _24139_/CLK _24143_/D HRESETn VGND VGND VPWR VPWR _24143_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13388__A _13388_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25092__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21355_ _21354_/X VGND VGND VPWR VPWR _21355_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20306_ _18240_/A VGND VGND VPWR VPWR _20306_/X sky130_fd_sc_hd__buf_2
XANTENNA__25021__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24074_ _24074_/CLK _20530_/X HRESETn VGND VGND VPWR VPWR _24074_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21286_ _21131_/X _21224_/X _21286_/C _21285_/X VGND VGND VPWR VPWR _21287_/A sky130_fd_sc_hd__and4_4
XFILLER_135_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23025_ _22844_/A _23025_/B _23024_/X VGND VGND VPWR VPWR _23025_/X sky130_fd_sc_hd__and3_4
X_20237_ _20236_/Y _20234_/X _11788_/X _20234_/X VGND VGND VPWR VPWR _23452_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23309__B _23308_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20168_ _23478_/Q VGND VGND VPWR VPWR _20168_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23010__A1 _16564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19214__B1 _19122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12990_ _12990_/A _13059_/A _12989_/X VGND VGND VPWR VPWR _12993_/B sky130_fd_sc_hd__or3_4
X_20099_ _20099_/A VGND VGND VPWR VPWR _20099_/X sky130_fd_sc_hd__buf_2
X_24976_ _24976_/CLK _24976_/D HRESETn VGND VGND VPWR VPWR _15087_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_162_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16028__B1 _15951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11941_ _11945_/A _11940_/A _18901_/A _11929_/X VGND VGND VPWR VPWR _11942_/B sky130_fd_sc_hd__and4_4
X_23927_ _23927_/CLK _23927_/D HRESETn VGND VGND VPWR VPWR _23927_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_217_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19522__B _14181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17776__B1 _16952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14660_ _20199_/B VGND VGND VPWR VPWR _19141_/B sky130_fd_sc_hd__buf_2
X_11872_ _11797_/Y _11799_/A VGND VGND VPWR VPWR _11872_/X sky130_fd_sc_hd__and2_4
X_23858_ _23754_/CLK _23858_/D VGND VGND VPWR VPWR _23858_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__24122__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13611_ _25073_/Q VGND VGND VPWR VPWR _13612_/A sky130_fd_sc_hd__inv_2
X_22809_ _16578_/A _22807_/X _21737_/X _22808_/X VGND VGND VPWR VPWR _22810_/C sky130_fd_sc_hd__a211o_4
X_14591_ _13757_/Y VGND VGND VPWR VPWR _14591_/X sky130_fd_sc_hd__buf_2
XFILLER_232_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23789_ _23464_/CLK _19291_/X VGND VGND VPWR VPWR _23789_/Q sky130_fd_sc_hd__dfxtp_4
X_16330_ _16329_/Y _16325_/X _16236_/X _16325_/X VGND VGND VPWR VPWR _24624_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13542_ _13542_/A VGND VGND VPWR VPWR _22734_/A sky130_fd_sc_hd__inv_2
X_25528_ _24947_/CLK _25528_/D HRESETn VGND VGND VPWR VPWR _25528_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21875__A2 _21030_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23956__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16261_ _24649_/Q VGND VGND VPWR VPWR _16261_/Y sky130_fd_sc_hd__inv_2
X_13473_ _25320_/Q VGND VGND VPWR VPWR _13473_/Y sky130_fd_sc_hd__inv_2
X_25459_ _25453_/CLK _12401_/Y HRESETn VGND VGND VPWR VPWR _25459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14682__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18154__A _18014_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18000_ _18118_/A _19008_/A VGND VGND VPWR VPWR _18000_/X sky130_fd_sc_hd__or2_4
XFILLER_185_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15212_ _15207_/A _15207_/B _15194_/X _15209_/B VGND VGND VPWR VPWR _15212_/X sky130_fd_sc_hd__a211o_4
X_12424_ _12272_/Y _12422_/A VGND VGND VPWR VPWR _12424_/X sky130_fd_sc_hd__or2_4
XANTENNA__25109__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16192_ _16189_/Y _16185_/X _15996_/X _16191_/X VGND VGND VPWR VPWR _24676_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15143_ _15082_/Y _24606_/Q _24996_/Q _15142_/Y VGND VGND VPWR VPWR _15143_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13298__A _13199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17993__A _18054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12355_ _13005_/A _24846_/Q _25355_/Q _12354_/Y VGND VGND VPWR VPWR _12355_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_181_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12286_ _25341_/Q _12284_/Y _12285_/Y _24847_/Q VGND VGND VPWR VPWR _12289_/C sky130_fd_sc_hd__a2bb2o_4
X_15074_ _15153_/A _15072_/Y _15326_/A _15085_/A VGND VGND VPWR VPWR _15074_/X sky130_fd_sc_hd__a2bb2o_4
X_19951_ _21801_/B _19946_/X _19613_/X _19946_/X VGND VGND VPWR VPWR _23558_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22588__B1 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14025_ _23929_/Q _14020_/Y _14024_/Y VGND VGND VPWR VPWR _14532_/C sky130_fd_sc_hd__or3_4
X_18902_ _11945_/Y _18902_/B _18902_/C _18902_/D VGND VGND VPWR VPWR _18902_/X sky130_fd_sc_hd__or4_4
X_19882_ _22246_/B _19879_/X _19603_/X _19879_/X VGND VGND VPWR VPWR _23585_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16402__A HWDATA[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18833_ _16530_/Y _18683_/A _16530_/Y _18683_/A VGND VGND VPWR VPWR _18833_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24744__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18764_ _18752_/A _18764_/B _18763_/X VGND VGND VPWR VPWR _24143_/D sky130_fd_sc_hd__and3_4
XANTENNA__15018__A _15018_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15976_ _15472_/A VGND VGND VPWR VPWR _15976_/X sky130_fd_sc_hd__buf_2
XFILLER_48_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17715_ _21475_/A _17714_/X _21475_/A _17714_/X VGND VGND VPWR VPWR _18313_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_236_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14927_ _25017_/Q VGND VGND VPWR VPWR _15058_/A sky130_fd_sc_hd__inv_2
XFILLER_64_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18695_ _18745_/D _18695_/B VGND VGND VPWR VPWR _18695_/X sky130_fd_sc_hd__or2_4
XFILLER_63_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13761__A _13807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17646_ _17646_/A _17643_/B VGND VGND VPWR VPWR _17646_/Y sky130_fd_sc_hd__nand2_4
X_14858_ _14838_/A _14857_/Y _14808_/C _14838_/A VGND VGND VPWR VPWR _25045_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_17_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13809_ _13832_/A VGND VGND VPWR VPWR _13810_/A sky130_fd_sc_hd__buf_2
XFILLER_51_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17577_ _17575_/Y _17521_/Y _17577_/C _17499_/Y VGND VGND VPWR VPWR _17581_/B sky130_fd_sc_hd__or4_4
XFILLER_223_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14789_ _13579_/X _13588_/X _14788_/Y _25057_/Q _14611_/Y VGND VGND VPWR VPWR _25057_/D
+ sky130_fd_sc_hd__a32o_4
X_19316_ _19315_/Y _19313_/X _19203_/X _19313_/X VGND VGND VPWR VPWR _23780_/D sky130_fd_sc_hd__a2bb2o_4
X_16528_ _16453_/A VGND VGND VPWR VPWR _16528_/X sky130_fd_sc_hd__buf_2
XFILLER_176_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19247_ _19247_/A VGND VGND VPWR VPWR _21386_/B sky130_fd_sc_hd__inv_2
XFILLER_149_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25532__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16459_ HWDATA[29] VGND VGND VPWR VPWR _16459_/X sky130_fd_sc_hd__buf_2
X_19178_ _19176_/Y _19177_/X _19063_/X _19177_/X VGND VGND VPWR VPWR _23829_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_192_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18129_ _18097_/A _23822_/Q VGND VGND VPWR VPWR _18129_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_104_0_HCLK clkbuf_7_52_0_HCLK/X VGND VGND VPWR VPWR _24346_/CLK sky130_fd_sc_hd__clkbuf_1
X_21140_ _14481_/Y _21155_/B _14171_/Y _21365_/A VGND VGND VPWR VPWR _21141_/D sky130_fd_sc_hd__o22a_4
Xclkbuf_8_167_0_HCLK clkbuf_7_83_0_HCLK/X VGND VGND VPWR VPWR _23887_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_160_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21071_ _21040_/X _21069_/X _21047_/X _21070_/X VGND VGND VPWR VPWR _21072_/C sky130_fd_sc_hd__a211o_4
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16258__B1 _15466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20022_ _20022_/A VGND VGND VPWR VPWR _20022_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24485__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24830_ _24804_/CLK _24830_/D HRESETn VGND VGND VPWR VPWR _24830_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24414__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23145__A _22146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24761_ _24763_/CLK _15961_/X HRESETn VGND VGND VPWR VPWR _24761_/Q sky130_fd_sc_hd__dfrtp_4
X_21973_ _24230_/Q _21958_/B VGND VGND VPWR VPWR _21973_/X sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_2_0_0_HCLK_A clkbuf_1_0_1_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22751__B1 _16035_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23712_ _23437_/CLK _19509_/X VGND VGND VPWR VPWR _23712_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ _20919_/X _20922_/X _24500_/Q _20923_/X VGND VGND VPWR VPWR _24056_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24692_ _24744_/CLK _16137_/X HRESETn VGND VGND VPWR VPWR _22602_/A sky130_fd_sc_hd__dfrtp_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _20827_/A VGND VGND VPWR VPWR _20855_/X sky130_fd_sc_hd__buf_2
X_23643_ _23644_/CLK _19714_/X VGND VGND VPWR VPWR _13442_/B sky130_fd_sc_hd__dfxtp_4
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16981__A1 _24725_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20786_ _20754_/X _13122_/B VGND VGND VPWR VPWR _20786_/Y sky130_fd_sc_hd__nor2_4
X_23574_ _23575_/CLK _19910_/X VGND VGND VPWR VPWR _19909_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25313_ _25492_/CLK _25313_/D HRESETn VGND VGND VPWR VPWR _13490_/A sky130_fd_sc_hd__dfrtp_4
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22525_ _22525_/A _21748_/A VGND VGND VPWR VPWR _22525_/X sky130_fd_sc_hd__or2_4
XFILLER_194_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25244_ _25204_/CLK _13872_/X HRESETn VGND VGND VPWR VPWR _25244_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22456_ _22450_/X _22453_/X _22454_/X _22455_/X VGND VGND VPWR VPWR _22457_/B sky130_fd_sc_hd__o22a_4
XFILLER_148_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_7_63_0_HCLK clkbuf_7_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_63_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21407_ _21403_/X _21406_/X _21247_/X VGND VGND VPWR VPWR _21407_/X sky130_fd_sc_hd__o21a_4
X_22387_ _22387_/A _22387_/B VGND VGND VPWR VPWR _22387_/X sky130_fd_sc_hd__or2_4
X_25175_ _23884_/CLK _14305_/X HRESETn VGND VGND VPWR VPWR _25175_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19683__B1 _19587_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12140_ _12140_/A VGND VGND VPWR VPWR _12140_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16497__B1 _16320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21338_ _21338_/A VGND VGND VPWR VPWR _23178_/A sky130_fd_sc_hd__buf_2
X_24126_ _24133_/CLK _18824_/X HRESETn VGND VGND VPWR VPWR _18681_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__22224__A _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12071_ _25481_/Q VGND VGND VPWR VPWR _12071_/Y sky130_fd_sc_hd__inv_2
X_21269_ _21262_/A _21269_/B VGND VGND VPWR VPWR _21269_/X sky130_fd_sc_hd__or2_4
X_24057_ _24501_/CLK _24057_/D HRESETn VGND VGND VPWR VPWR _24057_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16956__A1_N _15980_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23008_ _16207_/A _22729_/B VGND VGND VPWR VPWR _23008_/X sky130_fd_sc_hd__or2_4
X_15830_ _11774_/A VGND VGND VPWR VPWR _15830_/X sky130_fd_sc_hd__buf_2
XANTENNA__24155__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15761_ _15699_/Y VGND VGND VPWR VPWR _15761_/X sky130_fd_sc_hd__buf_2
XFILLER_92_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15780__B _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12973_ _25363_/Q VGND VGND VPWR VPWR _13000_/A sky130_fd_sc_hd__inv_2
X_24959_ _24959_/CLK _24959_/D HRESETn VGND VGND VPWR VPWR _13876_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_73_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14677__A _22056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17500_ _24317_/Q VGND VGND VPWR VPWR _17585_/A sky130_fd_sc_hd__inv_2
XANTENNA__21545__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14712_ _13721_/Y _13747_/Y _25280_/Q _13746_/X VGND VGND VPWR VPWR _14712_/X sky130_fd_sc_hd__o22a_4
XFILLER_205_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17053__A _17381_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11924_ _19617_/A VGND VGND VPWR VPWR _11924_/X sky130_fd_sc_hd__buf_2
X_18480_ _18510_/D _18479_/X VGND VGND VPWR VPWR _18480_/X sky130_fd_sc_hd__or2_4
X_15692_ _15676_/Y _15686_/A _15691_/X VGND VGND VPWR VPWR _15692_/X sky130_fd_sc_hd__o21a_4
XANTENNA__16421__B1 _16420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17431_ _24327_/Q VGND VGND VPWR VPWR _17431_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14643_ _13592_/B _14630_/C _17942_/A _14642_/X VGND VGND VPWR VPWR _25076_/D sky130_fd_sc_hd__a22oi_4
X_11855_ _25514_/Q VGND VGND VPWR VPWR _11856_/A sky130_fd_sc_hd__inv_2
XANTENNA__13731__D _14764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12197__A _12197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17362_ _17346_/C _17346_/D VGND VGND VPWR VPWR _17366_/B sky130_fd_sc_hd__or2_4
XFILLER_220_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14574_ _14570_/B _14546_/X _14573_/X _13758_/X _14563_/A VGND VGND VPWR VPWR _25095_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21848__A2 _14212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11786_ _15472_/A VGND VGND VPWR VPWR _11786_/X sky130_fd_sc_hd__buf_2
XPHY_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19101_ _19101_/A VGND VGND VPWR VPWR _19101_/X sky130_fd_sc_hd__buf_2
XFILLER_201_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16313_ _24630_/Q VGND VGND VPWR VPWR _16313_/Y sky130_fd_sc_hd__inv_2
X_13525_ _15908_/A VGND VGND VPWR VPWR _13525_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21303__A _21303_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17293_ _17236_/A _17290_/X VGND VGND VPWR VPWR _17294_/C sky130_fd_sc_hd__or2_4
X_19032_ _18046_/B VGND VGND VPWR VPWR _19032_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16244_ _16244_/A VGND VGND VPWR VPWR _16244_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13456_ _13482_/B VGND VGND VPWR VPWR _13456_/X sky130_fd_sc_hd__buf_2
X_12407_ _12172_/Y _12405_/A VGND VGND VPWR VPWR _12408_/C sky130_fd_sc_hd__or2_4
X_16175_ _14758_/A _16174_/Y _14756_/A _16174_/Y VGND VGND VPWR VPWR _16175_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19708__A _11785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13387_ _13186_/X _13386_/X _25328_/Q _13245_/X VGND VGND VPWR VPWR _13387_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24996__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15126_ _15125_/Y _22701_/A _15125_/Y _22701_/A VGND VGND VPWR VPWR _15127_/D sky130_fd_sc_hd__a2bb2o_4
X_12338_ _12976_/D _24834_/Q _12976_/D _24834_/Q VGND VGND VPWR VPWR _12339_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24925__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15057_ _14970_/Y _15273_/A _15272_/A VGND VGND VPWR VPWR _15243_/A sky130_fd_sc_hd__or3_4
X_19934_ _19934_/A VGND VGND VPWR VPWR _21474_/B sky130_fd_sc_hd__inv_2
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21350__A1_N _14166_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12269_ _12269_/A _12211_/Y _12492_/A VGND VGND VPWR VPWR _12270_/D sky130_fd_sc_hd__or3_4
X_14008_ _14008_/A _14007_/D _14007_/A _13969_/Y VGND VGND VPWR VPWR _14008_/X sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_5_17_0_HCLK_A clkbuf_4_8_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19865_ _19864_/Y _19862_/X _19610_/X _19862_/X VGND VGND VPWR VPWR _19865_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22981__B1 _25541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18816_ _18819_/A _18815_/X VGND VGND VPWR VPWR _18820_/B sky130_fd_sc_hd__or2_4
XFILLER_96_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19796_ _19784_/A VGND VGND VPWR VPWR _19796_/X sky130_fd_sc_hd__buf_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15959_ _15955_/X _15958_/X _16226_/A _24763_/Q _15956_/X VGND VGND VPWR VPWR _24763_/D
+ sky130_fd_sc_hd__a32o_4
X_18747_ _18747_/A _18746_/X VGND VGND VPWR VPWR _18748_/B sky130_fd_sc_hd__or2_4
XFILLER_209_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13474__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_243_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18678_ _18733_/A _18730_/A VGND VGND VPWR VPWR _18696_/C sky130_fd_sc_hd__or2_4
XFILLER_36_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16412__B1 _16229_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17629_ _17570_/X _17637_/B VGND VGND VPWR VPWR _17629_/X sky130_fd_sc_hd__or2_4
X_20640_ _20640_/A _20639_/Y _20621_/C VGND VGND VPWR VPWR _20640_/X sky130_fd_sc_hd__and3_4
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21213__A _21178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20571_ _18877_/A _18876_/X VGND VGND VPWR VPWR _20571_/Y sky130_fd_sc_hd__nand2_4
XFILLER_177_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22310_ _24453_/Q _21309_/X _22891_/A VGND VGND VPWR VPWR _22310_/X sky130_fd_sc_hd__o21a_4
X_23290_ _23288_/X _23289_/X _22140_/A VGND VGND VPWR VPWR _23290_/X sky130_fd_sc_hd__or3_4
XFILLER_165_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22241_ _22007_/X _22238_/X _22241_/C VGND VGND VPWR VPWR _22241_/X sky130_fd_sc_hd__and3_4
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21867__B _21855_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19665__B1 _19540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22172_ _22171_/X VGND VGND VPWR VPWR _22174_/C sky130_fd_sc_hd__inv_2
XANTENNA__24666__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21318__A1_N _17203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21123_ _22840_/A VGND VGND VPWR VPWR _21124_/B sky130_fd_sc_hd__buf_2
XANTENNA__19417__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21054_ _11664_/B VGND VGND VPWR VPWR _22189_/A sky130_fd_sc_hd__inv_2
XFILLER_113_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11712__B1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20005_ _23540_/Q VGND VGND VPWR VPWR _21471_/B sky130_fd_sc_hd__inv_2
XFILLER_59_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_HCLK clkbuf_3_2_0_HCLK/X VGND VGND VPWR VPWR clkbuf_4_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__16651__B1 _16467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24813_ _25373_/CLK _24813_/D HRESETn VGND VGND VPWR VPWR _23219_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13465__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11914__A _19613_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24744_ _24744_/CLK _16002_/X HRESETn VGND VGND VPWR VPWR _24744_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21956_ _21956_/A VGND VGND VPWR VPWR _21956_/X sky130_fd_sc_hd__buf_2
XANTENNA__17304__C _17343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16403__B1 _16402_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _24052_/Q _24053_/Q _24051_/Q _20921_/C VGND VGND VPWR VPWR _20907_/X sky130_fd_sc_hd__or4_4
XFILLER_199_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25454__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24675_ _24675_/CLK _16194_/X HRESETn VGND VGND VPWR VPWR _23238_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21887_ _22056_/A VGND VGND VPWR VPWR _22083_/A sky130_fd_sc_hd__buf_2
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _23610_/CLK _23626_/D VGND VGND VPWR VPWR _19761_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _24038_/Q VGND VGND VPWR VPWR _20838_/Y sky130_fd_sc_hd__inv_2
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22219__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21123__A _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23557_ _25285_/CLK _23557_/D VGND VGND VPWR VPWR _23557_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_167_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20769_ _20767_/Y _20764_/X _20768_/X VGND VGND VPWR VPWR _20769_/X sky130_fd_sc_hd__o21a_4
XFILLER_50_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16217__A _22883_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _13433_/A VGND VGND VPWR VPWR _13310_/X sky130_fd_sc_hd__buf_2
XFILLER_156_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22508_ _21587_/A _22507_/X VGND VGND VPWR VPWR _22508_/Y sky130_fd_sc_hd__nor2_4
X_14290_ _14290_/A _14285_/X _14290_/C VGND VGND VPWR VPWR _25180_/D sky130_fd_sc_hd__and3_4
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23488_ _23490_/CLK _23488_/D VGND VGND VPWR VPWR _23488_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ _13150_/X _13236_/X _13241_/C VGND VGND VPWR VPWR _13241_/X sky130_fd_sc_hd__or3_4
X_25227_ _25238_/CLK _25227_/D HRESETn VGND VGND VPWR VPWR _14022_/B sky130_fd_sc_hd__dfrtp_4
X_22439_ _12192_/Y _22417_/B _22275_/X _12306_/Y _22129_/X VGND VGND VPWR VPWR _22439_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13172_ _13172_/A _13170_/X _13171_/X VGND VGND VPWR VPWR _13172_/X sky130_fd_sc_hd__and3_4
X_25158_ _25158_/CLK _25158_/D HRESETn VGND VGND VPWR VPWR _25158_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15775__B _15670_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12123_ _25473_/Q _20971_/A _12101_/Y _12122_/Y VGND VGND VPWR VPWR _12133_/A sky130_fd_sc_hd__o22a_4
X_24109_ _23932_/CLK MSI_S3 HRESETn VGND VGND VPWR VPWR _24109_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13576__A _14764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17980_ _17979_/X _17980_/B VGND VGND VPWR VPWR _17981_/C sky130_fd_sc_hd__or2_4
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25089_ _25089_/CLK _14589_/X HRESETn VGND VGND VPWR VPWR _13535_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_151_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23204__B2 _21315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_150_0_HCLK clkbuf_7_75_0_HCLK/X VGND VGND VPWR VPWR _25474_/CLK sky130_fd_sc_hd__clkbuf_1
X_12054_ _11667_/A VGND VGND VPWR VPWR _12083_/A sky130_fd_sc_hd__buf_2
X_16931_ _16106_/Y _17744_/A _16106_/Y _17744_/A VGND VGND VPWR VPWR _16934_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15791__A _15811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16862_ _24411_/Q VGND VGND VPWR VPWR _16863_/A sky130_fd_sc_hd__buf_2
X_19650_ _19650_/A VGND VGND VPWR VPWR _19650_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18631__A1 _24544_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15813_ _15813_/A VGND VGND VPWR VPWR _15813_/X sky130_fd_sc_hd__buf_2
X_18601_ _24157_/Q VGND VGND VPWR VPWR _18703_/A sky130_fd_sc_hd__buf_2
XFILLER_93_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19581_ _19576_/A VGND VGND VPWR VPWR _19581_/X sky130_fd_sc_hd__buf_2
XFILLER_92_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16793_ _16793_/A VGND VGND VPWR VPWR _16793_/X sky130_fd_sc_hd__buf_2
XFILLER_219_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18532_ _18531_/X VGND VGND VPWR VPWR _18532_/Y sky130_fd_sc_hd__inv_2
X_15744_ _15724_/X _15738_/X _15743_/X _24868_/Q _15736_/X VGND VGND VPWR VPWR _24868_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_80_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12956_ _12807_/X _12929_/X _12872_/A _12954_/B VGND VGND VPWR VPWR _12956_/X sky130_fd_sc_hd__a211o_4
XFILLER_18_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11907_ _11897_/X VGND VGND VPWR VPWR _11907_/X sky130_fd_sc_hd__buf_2
X_18463_ _24174_/Q VGND VGND VPWR VPWR _18466_/B sky130_fd_sc_hd__inv_2
XFILLER_34_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15675_ _15675_/A VGND VGND VPWR VPWR _15675_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12887_ _12887_/A _12884_/B _12886_/X VGND VGND VPWR VPWR _12888_/A sky130_fd_sc_hd__or3_4
XPHY_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17429_/A VGND VGND VPWR VPWR _17414_/X sky130_fd_sc_hd__buf_2
XPHY_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _18060_/A VGND VGND VPWR VPWR _17950_/A sky130_fd_sc_hd__buf_2
XFILLER_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25124__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11838_ _25290_/Q VGND VGND VPWR VPWR _13676_/A sky130_fd_sc_hd__inv_2
X_18394_ _16177_/Y _24189_/Q _16177_/Y _24189_/Q VGND VGND VPWR VPWR _18394_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22129__A _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17345_/A _17345_/B VGND VGND VPWR VPWR _17346_/D sky130_fd_sc_hd__or2_4
XPHY_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/A _14557_/B VGND VGND VPWR VPWR _14557_/X sky130_fd_sc_hd__or2_4
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11769_ HWDATA[5] VGND VGND VPWR VPWR _13829_/A sky130_fd_sc_hd__buf_2
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13508_ _25181_/Q _14289_/A _14278_/A _13508_/D VGND VGND VPWR VPWR _13509_/B sky130_fd_sc_hd__and4_4
X_17276_ _17284_/A VGND VGND VPWR VPWR _17276_/X sky130_fd_sc_hd__buf_2
X_14488_ _23393_/Q _20453_/C _14487_/A _25113_/Q _14487_/Y VGND VGND VPWR VPWR _14488_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19015_ _18118_/B VGND VGND VPWR VPWR _19015_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16227_ _16225_/Y _16223_/X _16226_/X _16223_/X VGND VGND VPWR VPWR _24662_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18859__A2_N _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13439_ _13234_/X _13439_/B VGND VGND VPWR VPWR _13439_/X sky130_fd_sc_hd__or2_4
XFILLER_162_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19647__B1 _19646_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16158_ _16157_/Y _16155_/X _15469_/X _16155_/X VGND VGND VPWR VPWR _16158_/X sky130_fd_sc_hd__a2bb2o_4
X_15109_ _24978_/Q VGND VGND VPWR VPWR _15296_/B sky130_fd_sc_hd__inv_2
X_16089_ _16088_/Y _16086_/X _15554_/X _16086_/X VGND VGND VPWR VPWR _16089_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24077__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19917_ _21260_/B _19912_/X _19852_/X _19900_/A VGND VGND VPWR VPWR _19917_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_244_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24006__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19848_ _19846_/Y _19847_/X _19824_/X _19847_/X VGND VGND VPWR VPWR _19848_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_229_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19779_ _19778_/Y _19776_/X _16885_/X _19776_/X VGND VGND VPWR VPWR _23620_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11734__A HWDATA[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21810_ _21677_/A _19976_/Y VGND VGND VPWR VPWR _21811_/C sky130_fd_sc_hd__or2_4
XFILLER_209_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17423__A2_N _17414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22790_ _22684_/B VGND VGND VPWR VPWR _22989_/B sky130_fd_sc_hd__buf_2
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22182__B2 _21351_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22965__C _22957_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21741_ _16530_/Y _21741_/B VGND VGND VPWR VPWR _21741_/X sky130_fd_sc_hd__and2_4
XFILLER_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17421__A _14407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24460_ _24460_/CLK _16761_/X HRESETn VGND VGND VPWR VPWR _24460_/Q sky130_fd_sc_hd__dfrtp_4
X_21672_ _21677_/A _21672_/B VGND VGND VPWR VPWR _21673_/C sky130_fd_sc_hd__or2_4
Xclkbuf_4_13_0_HCLK clkbuf_3_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_27_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23411_ _23411_/CLK _20344_/X VGND VGND VPWR VPWR _23411_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20623_ _20623_/A VGND VGND VPWR VPWR _23976_/D sky130_fd_sc_hd__inv_2
XFILLER_196_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24391_ _24315_/CLK _24391_/D HRESETn VGND VGND VPWR VPWR _24391_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16037__A _24730_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20554_ _14433_/Y _20543_/X _20600_/A _20553_/X VGND VGND VPWR VPWR _20555_/A sky130_fd_sc_hd__a211o_4
X_23342_ _13774_/Y _23342_/B VGND VGND VPWR VPWR _23342_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__24847__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19348__A _19343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20485_ _23966_/Q _20524_/B VGND VGND VPWR VPWR _20485_/X sky130_fd_sc_hd__and2_4
X_23273_ _23268_/Y _23272_/Y _22854_/X VGND VGND VPWR VPWR _23273_/X sky130_fd_sc_hd__o21a_4
X_25012_ _25015_/CLK _25012_/D HRESETn VGND VGND VPWR VPWR _25012_/Q sky130_fd_sc_hd__dfrtp_4
X_22224_ _22221_/A _22224_/B VGND VGND VPWR VPWR _22224_/X sky130_fd_sc_hd__or2_4
XANTENNA__24089__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22155_ _21055_/X _22154_/X VGND VGND VPWR VPWR _22155_/X sky130_fd_sc_hd__and2_4
XFILLER_133_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23198__B1 _12735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21106_ _21736_/A _21105_/Y _24644_/Q _21736_/A VGND VGND VPWR VPWR _21106_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_223_0_HCLK clkbuf_8_222_0_HCLK/A VGND VGND VPWR VPWR _25035_/CLK sky130_fd_sc_hd__clkbuf_1
X_22086_ _22378_/A _19839_/Y _21627_/A VGND VGND VPWR VPWR _22086_/X sky130_fd_sc_hd__o21a_4
XFILLER_154_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12489__A1 _12252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21037_ _24785_/Q _21064_/B VGND VGND VPWR VPWR _21037_/X sky130_fd_sc_hd__or2_4
XANTENNA__12331__A2_N _12329_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22960__A3 _22849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12810_ _24805_/Q VGND VGND VPWR VPWR _12810_/Y sky130_fd_sc_hd__inv_2
X_13790_ _25273_/Q VGND VGND VPWR VPWR _13790_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22988_ _16665_/Y _22921_/B VGND VGND VPWR VPWR _22988_/X sky130_fd_sc_hd__and2_4
XANTENNA__22173__B2 _22181_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12741_ _12838_/D VGND VGND VPWR VPWR _12741_/X sky130_fd_sc_hd__buf_2
X_24727_ _24266_/CLK _24727_/D HRESETn VGND VGND VPWR VPWR _24727_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23333__A _16363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_0_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_21939_ _21453_/X _21928_/X _21939_/C VGND VGND VPWR VPWR _21939_/X sky130_fd_sc_hd__or3_4
XFILLER_216_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15460_ _24957_/Q VGND VGND VPWR VPWR _15460_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14938__B1 _15261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12672_ _12677_/A _12672_/B _12671_/Y VGND VGND VPWR VPWR _25418_/D sky130_fd_sc_hd__and3_4
X_24658_ _24678_/CLK _16241_/X HRESETn VGND VGND VPWR VPWR _22590_/A sky130_fd_sc_hd__dfrtp_4
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14410_/Y _14408_/X _14380_/X _14408_/X VGND VGND VPWR VPWR _14411_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _23497_/CLK _19811_/X VGND VGND VPWR VPWR _23609_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _15068_/Y _15394_/B _15334_/X VGND VGND VPWR VPWR _15391_/Y sky130_fd_sc_hd__a21oi_4
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24589_ _24985_/CLK _16423_/X HRESETn VGND VGND VPWR VPWR _15107_/A sky130_fd_sc_hd__dfrtp_4
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _16971_/Y _17129_/X VGND VGND VPWR VPWR _17140_/B sky130_fd_sc_hd__or2_4
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _14342_/A VGND VGND VPWR VPWR _25162_/D sky130_fd_sc_hd__inv_2
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24588__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17061_ _17070_/A _17061_/B _17060_/X VGND VGND VPWR VPWR _24402_/D sky130_fd_sc_hd__and3_4
XFILLER_7_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15786__A _15811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14273_ _14273_/A VGND VGND VPWR VPWR _14273_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24517__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16012_ _15998_/A VGND VGND VPWR VPWR _16012_/X sky130_fd_sc_hd__buf_2
XFILLER_155_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13224_ _13219_/X _13224_/B _13223_/X VGND VGND VPWR VPWR _13224_/X sky130_fd_sc_hd__and3_4
XFILLER_124_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_33_0_HCLK clkbuf_6_33_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_67_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_3_0_HCLK_A clkbuf_3_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17501__A1_N _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13155_ _13172_/A _13152_/X _13155_/C VGND VGND VPWR VPWR _13155_/X sky130_fd_sc_hd__and3_4
XFILLER_151_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24170__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12106_ _25471_/Q VGND VGND VPWR VPWR _12106_/Y sky130_fd_sc_hd__inv_2
X_13086_ _12979_/D _13091_/A VGND VGND VPWR VPWR _13088_/B sky130_fd_sc_hd__nand2_4
X_17963_ _15673_/X _15680_/A _14608_/Y _15911_/X VGND VGND VPWR VPWR _17966_/A sky130_fd_sc_hd__a211o_4
XANTENNA__22412__A _24619_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19702_ _11774_/A VGND VGND VPWR VPWR _19702_/X sky130_fd_sc_hd__buf_2
X_12037_ _11660_/A VGND VGND VPWR VPWR _15636_/C sky130_fd_sc_hd__buf_2
X_16914_ _24710_/Q _16913_/A _16090_/Y _16913_/Y VGND VGND VPWR VPWR _16919_/B sky130_fd_sc_hd__o22a_4
XANTENNA__19801__B1 _19759_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17894_ _17892_/A VGND VGND VPWR VPWR _17894_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19633_ _18985_/A VGND VGND VPWR VPWR _19633_/X sky130_fd_sc_hd__buf_2
XANTENNA__21028__A _11701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25376__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16845_ _16793_/A VGND VGND VPWR VPWR _16845_/X sky130_fd_sc_hd__buf_2
XFILLER_226_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20962__A2 _14608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15026__A _15026_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16776_ _14986_/Y _16774_/X _16525_/X _16774_/X VGND VGND VPWR VPWR _24451_/D sky130_fd_sc_hd__a2bb2o_4
X_19564_ _23692_/Q VGND VGND VPWR VPWR _21495_/B sky130_fd_sc_hd__inv_2
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13988_ _13980_/A VGND VGND VPWR VPWR _13990_/C sky130_fd_sc_hd__buf_2
XFILLER_230_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22164__A1 _16520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15727_ _12574_/Y _15717_/X _11695_/X _15717_/X VGND VGND VPWR VPWR _15727_/X sky130_fd_sc_hd__a2bb2o_4
X_18515_ _18462_/B _18515_/B VGND VGND VPWR VPWR _18516_/C sky130_fd_sc_hd__nand2_4
X_12939_ _12939_/A VGND VGND VPWR VPWR _12939_/Y sky130_fd_sc_hd__inv_2
X_19495_ _19493_/Y _19494_/X _11924_/X _19494_/X VGND VGND VPWR VPWR _19495_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16918__A1 _21521_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16918__B2 _16917_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15658_ _21138_/A _17436_/C _11676_/B _15657_/X VGND VGND VPWR VPWR _15666_/A sky130_fd_sc_hd__or4_4
X_18446_ _18439_/X _18446_/B _18443_/X _18445_/X VGND VGND VPWR VPWR _18446_/X sky130_fd_sc_hd__or4_4
XFILLER_178_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14609_ _14608_/Y _15694_/A _13586_/A _13525_/Y VGND VGND VPWR VPWR _14610_/B sky130_fd_sc_hd__and4_4
X_18377_ _18376_/Y _18374_/X _24196_/Q _18374_/X VGND VGND VPWR VPWR _24197_/D sky130_fd_sc_hd__a2bb2o_4
X_15589_ _15576_/A VGND VGND VPWR VPWR _15589_/X sky130_fd_sc_hd__buf_2
XFILLER_194_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12385__A _12264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17328_ _24356_/Q _17327_/Y VGND VGND VPWR VPWR _17328_/X sky130_fd_sc_hd__or2_4
XFILLER_147_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_115_0_HCLK clkbuf_6_57_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_231_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__24940__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17259_ _17258_/X VGND VGND VPWR VPWR _17260_/B sky130_fd_sc_hd__inv_2
XFILLER_147_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24258__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20270_ _22259_/B _20267_/X _19967_/X _20267_/X VGND VGND VPWR VPWR _20270_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11729__A HWDATA[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21864__C _21864_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23960_ _23926_/CLK _23960_/D HRESETn VGND VGND VPWR VPWR _14369_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_57_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16320__A HWDATA[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22911_ _22908_/X _22909_/X _22495_/X _25539_/Q _22910_/X VGND VGND VPWR VPWR _22911_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_8_53_0_HCLK clkbuf_7_26_0_HCLK/X VGND VGND VPWR VPWR _25533_/CLK sky130_fd_sc_hd__clkbuf_1
X_23891_ _23889_/CLK _23891_/D VGND VGND VPWR VPWR _18218_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22842_ _15025_/A _23263_/B _23263_/C VGND VGND VPWR VPWR _22842_/X sky130_fd_sc_hd__and3_4
XANTENNA__25046__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24953__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22773_ _23043_/A _22773_/B VGND VGND VPWR VPWR _22781_/C sky130_fd_sc_hd__and2_4
XANTENNA__16909__A1 _22405_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24512_ _24679_/CLK _24512_/D HRESETn VGND VGND VPWR VPWR _13728_/A sky130_fd_sc_hd__dfrtp_4
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21724_ _21723_/Y _21159_/X _15468_/Y _21365_/X VGND VGND VPWR VPWR _21725_/A sky130_fd_sc_hd__o22a_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25492_ _25492_/CLK _25492_/D HRESETn VGND VGND VPWR VPWR _12022_/A sky130_fd_sc_hd__dfrtp_4
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22992__A _22992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24443_ _24443_/CLK _16800_/X HRESETn VGND VGND VPWR VPWR _24443_/Q sky130_fd_sc_hd__dfrtp_4
X_21655_ _21817_/A _21655_/B VGND VGND VPWR VPWR _21656_/C sky130_fd_sc_hd__or2_4
X_20606_ _20606_/A _20450_/X VGND VGND VPWR VPWR _20606_/X sky130_fd_sc_hd__or2_4
X_24374_ _24377_/CLK _24374_/D HRESETn VGND VGND VPWR VPWR _16990_/A sky130_fd_sc_hd__dfrtp_4
X_21586_ _16366_/B _21580_/X _16180_/X _21585_/X VGND VGND VPWR VPWR _21587_/B sky130_fd_sc_hd__o22a_4
XANTENNA__24681__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23325_ _22468_/A _23323_/Y _22469_/X _23324_/Y VGND VGND VPWR VPWR _23326_/B sky130_fd_sc_hd__o22a_4
X_20537_ _20436_/X _20505_/X _20453_/D _14484_/X _20444_/B VGND VGND VPWR VPWR _24084_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_181_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24610__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20468_ _20444_/X _20523_/B _20468_/C _20523_/A VGND VGND VPWR VPWR _20468_/X sky130_fd_sc_hd__or4_4
X_23256_ _12769_/Y _21879_/X _16913_/Y _22826_/X VGND VGND VPWR VPWR _23256_/X sky130_fd_sc_hd__o22a_4
XFILLER_165_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22207_ _22199_/A _19902_/Y VGND VGND VPWR VPWR _22207_/X sky130_fd_sc_hd__or2_4
XANTENNA__19806__A _19805_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20399_ _20398_/Y _20394_/X _15764_/X _20394_/X VGND VGND VPWR VPWR _20399_/X sky130_fd_sc_hd__a2bb2o_4
X_23187_ _23187_/A _23040_/X VGND VGND VPWR VPWR _23187_/X sky130_fd_sc_hd__or2_4
X_22138_ _21598_/X _22136_/X _22138_/C VGND VGND VPWR VPWR _22138_/X sky130_fd_sc_hd__and3_4
XANTENNA__23328__A _23328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22918__B1 _12766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14960_ _14995_/A _14966_/A _15026_/A _14895_/Y VGND VGND VPWR VPWR _14960_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22069_ _22069_/A VGND VGND VPWR VPWR _22383_/A sky130_fd_sc_hd__buf_2
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13911_ _13931_/A _13931_/B _13944_/A VGND VGND VPWR VPWR _13911_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_181_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14891_ _14882_/X _14891_/B _14891_/C _14891_/D VGND VGND VPWR VPWR _14935_/A sky130_fd_sc_hd__or4_4
X_16630_ _24513_/Q _16629_/Y _16624_/X VGND VGND VPWR VPWR _24513_/D sky130_fd_sc_hd__o21a_4
X_13842_ _25254_/Q _13842_/B VGND VGND VPWR VPWR _13842_/Y sky130_fd_sc_hd__nor2_4
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20687__A _20708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16561_ _16559_/Y _16555_/X _16386_/X _16560_/X VGND VGND VPWR VPWR _16561_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13773_ _13758_/X _13772_/X _13459_/X _13772_/X VGND VGND VPWR VPWR _13773_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13831__B1 _13785_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15512_ _15530_/A VGND VGND VPWR VPWR _15512_/X sky130_fd_sc_hd__buf_2
X_18300_ _18296_/A VGND VGND VPWR VPWR _18301_/A sky130_fd_sc_hd__buf_2
X_12724_ _12724_/A _12724_/B VGND VGND VPWR VPWR _12725_/B sky130_fd_sc_hd__or2_4
X_19280_ _19278_/Y _19276_/X _19279_/X _19276_/X VGND VGND VPWR VPWR _23793_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16492_ _16492_/A VGND VGND VPWR VPWR _16492_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24769__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18231_ _21958_/B VGND VGND VPWR VPWR _21962_/A sky130_fd_sc_hd__buf_2
XFILLER_230_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15443_ _14269_/X _24072_/Q _15436_/Y _13930_/A _15439_/X VGND VGND VPWR VPWR _24968_/D
+ sky130_fd_sc_hd__a32o_4
X_12655_ _12655_/A _12655_/B VGND VGND VPWR VPWR _12656_/A sky130_fd_sc_hd__or2_4
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17996__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18162_ _18098_/A _18160_/X _18161_/X VGND VGND VPWR VPWR _18163_/C sky130_fd_sc_hd__and3_4
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _15331_/A _15300_/C VGND VGND VPWR VPWR _15375_/B sky130_fd_sc_hd__or2_4
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _12586_/A _12581_/X _12582_/X _12586_/D VGND VGND VPWR VPWR _12586_/X sky130_fd_sc_hd__or4_4
XFILLER_196_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17113_ _17030_/D _17097_/B _17064_/X _17111_/B VGND VGND VPWR VPWR _17113_/X sky130_fd_sc_hd__a211o_4
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _25166_/Q _14339_/A _14332_/B VGND VGND VPWR VPWR _14325_/X sky130_fd_sc_hd__and3_4
XFILLER_209_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18093_ _18126_/A _23839_/Q VGND VGND VPWR VPWR _18093_/X sky130_fd_sc_hd__or2_4
XFILLER_128_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24351__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17044_ _17032_/X _17088_/B VGND VGND VPWR VPWR _17045_/D sky130_fd_sc_hd__or2_4
X_14256_ _14256_/A VGND VGND VPWR VPWR _14256_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13207_ _13249_/A VGND VGND VPWR VPWR _13392_/A sky130_fd_sc_hd__buf_2
XFILLER_125_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22082__B1 _14666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14187_ _20628_/A _14187_/B VGND VGND VPWR VPWR _14189_/A sky130_fd_sc_hd__nor2_4
XFILLER_125_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16836__B1 _15965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12238__A2_N _24763_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13138_ _13189_/A VGND VGND VPWR VPWR _13249_/A sky130_fd_sc_hd__inv_2
X_18995_ _23892_/Q VGND VGND VPWR VPWR _18995_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17236__A _17236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13069_ _13069_/A _13069_/B VGND VGND VPWR VPWR _13089_/A sky130_fd_sc_hd__or2_4
X_17946_ _17942_/X _17945_/X _18009_/A VGND VGND VPWR VPWR _17947_/C sky130_fd_sc_hd__o21a_4
XFILLER_112_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16140__A _22494_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13483__B _12086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17877_ _17866_/A _17873_/B _17877_/C VGND VGND VPWR VPWR _24263_/D sky130_fd_sc_hd__and3_4
XFILLER_227_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19616_ _19598_/Y VGND VGND VPWR VPWR _19616_/X sky130_fd_sc_hd__buf_2
X_16828_ _16826_/Y _16822_/X _15741_/X _16827_/X VGND VGND VPWR VPWR _16828_/X sky130_fd_sc_hd__a2bb2o_4
X_19547_ _19547_/A VGND VGND VPWR VPWR _22353_/B sky130_fd_sc_hd__inv_2
XFILLER_65_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16759_ _24460_/Q VGND VGND VPWR VPWR _16759_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19478_ _18285_/A VGND VGND VPWR VPWR _19939_/A sky130_fd_sc_hd__buf_2
XFILLER_61_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18429_ _24163_/Q VGND VGND VPWR VPWR _18563_/A sky130_fd_sc_hd__inv_2
XFILLER_22_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24439__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21440_ _21439_/X VGND VGND VPWR VPWR _23277_/A sky130_fd_sc_hd__buf_2
XANTENNA__22845__C1 _22844_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17316__A1 _17251_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18513__B1 _18489_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21371_ _14201_/Y _14182_/X _14261_/Y _21721_/B VGND VGND VPWR VPWR _21372_/D sky130_fd_sc_hd__o22a_4
XFILLER_135_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24092__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20322_ _23419_/Q VGND VGND VPWR VPWR _20322_/Y sky130_fd_sc_hd__inv_2
X_23110_ _23044_/X _23109_/X _23046_/X _16009_/A _22865_/X VGND VGND VPWR VPWR _23110_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24090_ _25308_/CLK _13633_/Y HRESETn VGND VGND VPWR VPWR _14290_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16034__A1_N _16031_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24021__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20253_ _21775_/B _20248_/X _19820_/A _20248_/X VGND VGND VPWR VPWR _23446_/D sky130_fd_sc_hd__a2bb2o_4
X_23041_ _24808_/Q _23040_/X VGND VGND VPWR VPWR _23041_/X sky130_fd_sc_hd__or2_4
XFILLER_115_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20184_ _20184_/A VGND VGND VPWR VPWR _22063_/B sky130_fd_sc_hd__inv_2
XFILLER_131_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23148__A _24811_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24992_ _24551_/CLK _24992_/D HRESETn VGND VGND VPWR VPWR _24992_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16050__A _16038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22987__A _22985_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23943_ _25140_/CLK _20575_/Y HRESETn VGND VGND VPWR VPWR _18877_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23874_ _23754_/CLK _23874_/D VGND VGND VPWR VPWR _19046_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23325__B1 _22469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22825_ _22721_/A VGND VGND VPWR VPWR _23268_/A sky130_fd_sc_hd__buf_2
XFILLER_56_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16602__A1_N _16600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22679__A2 _22992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25544_ _24310_/CLK _25544_/D HRESETn VGND VGND VPWR VPWR _11687_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_241_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22756_ _16679_/Y _22756_/B VGND VGND VPWR VPWR _22756_/X sky130_fd_sc_hd__and2_4
XANTENNA__24862__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21707_ _24615_/Q _22130_/B VGND VGND VPWR VPWR _21707_/X sky130_fd_sc_hd__or2_4
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25475_ _25474_/CLK _12098_/X HRESETn VGND VGND VPWR VPWR _12097_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_197_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22687_ _16272_/X _22676_/Y _22678_/Y _22682_/Y _22686_/Y VGND VGND VPWR VPWR _22687_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_200_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18705__A _18774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12440_ _12226_/X _12418_/X VGND VGND VPWR VPWR _12443_/B sky130_fd_sc_hd__or2_4
X_24426_ _24427_/CLK _16832_/X HRESETn VGND VGND VPWR VPWR _16831_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_212_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21638_ _21764_/A _21636_/X _21638_/C VGND VGND VPWR VPWR _21638_/X sky130_fd_sc_hd__and3_4
XFILLER_178_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24109__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22227__A _22212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13849__A _13839_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12371_ _12370_/X VGND VGND VPWR VPWR _12494_/A sky130_fd_sc_hd__buf_2
X_24357_ _24357_/CLK _17325_/Y HRESETn VGND VGND VPWR VPWR _24357_/Q sky130_fd_sc_hd__dfrtp_4
X_21569_ _21569_/A VGND VGND VPWR VPWR _21569_/X sky130_fd_sc_hd__buf_2
XANTENNA__22851__A2 _22523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14110_ _25145_/Q _14099_/X _14100_/X _14109_/Y VGND VGND VPWR VPWR _14110_/X sky130_fd_sc_hd__o22a_4
XFILLER_5_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23308_ _22129_/X _23307_/X _23145_/X _24851_/Q _22838_/X VGND VGND VPWR VPWR _23308_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_154_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15090_ _15090_/A VGND VGND VPWR VPWR _15291_/A sky130_fd_sc_hd__inv_2
X_24288_ _25444_/CLK _24288_/D HRESETn VGND VGND VPWR VPWR _24288_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14041_ _14004_/X _14041_/B VGND VGND VPWR VPWR _14049_/A sky130_fd_sc_hd__or2_4
X_23239_ _24575_/Q _23172_/X _23133_/X VGND VGND VPWR VPWR _23239_/X sky130_fd_sc_hd__o21a_4
XFILLER_192_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16818__B1 HWDATA[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22447__A1_N _17352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17800_ _17746_/A _17800_/B VGND VGND VPWR VPWR _17801_/C sky130_fd_sc_hd__or2_4
X_15992_ _15980_/Y _15990_/X _15991_/X _15990_/X VGND VGND VPWR VPWR _24747_/D sky130_fd_sc_hd__a2bb2o_4
X_18780_ _18694_/B _18774_/X _18735_/X _18777_/B VGND VGND VPWR VPWR _18780_/X sky130_fd_sc_hd__a211o_4
XFILLER_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22897__A _21087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14943_ _14942_/Y _16831_/A _14942_/Y _16831_/A VGND VGND VPWR VPWR _14943_/X sky130_fd_sc_hd__a2bb2o_4
X_17731_ _17730_/X VGND VGND VPWR VPWR _17731_/X sky130_fd_sc_hd__buf_2
XFILLER_236_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__20378__B1 _15762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14874_ _14874_/A VGND VGND VPWR VPWR _14874_/Y sky130_fd_sc_hd__inv_2
X_17662_ _17582_/B _17656_/X _17659_/B _17593_/X VGND VGND VPWR VPWR _17663_/A sky130_fd_sc_hd__a211o_4
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19401_ _19400_/Y _19396_/X _19377_/X _19396_/X VGND VGND VPWR VPWR _23750_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18991__B1 _18965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13825_ _13544_/Y _13822_/X _13824_/X _13822_/X VGND VGND VPWR VPWR _25262_/D sky130_fd_sc_hd__a2bb2o_4
X_16613_ _24518_/Q VGND VGND VPWR VPWR _16613_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21306__A _21303_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17593_ _17625_/A VGND VGND VPWR VPWR _17593_/X sky130_fd_sc_hd__buf_2
XFILLER_189_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16544_ _24545_/Q VGND VGND VPWR VPWR _16544_/Y sky130_fd_sc_hd__inv_2
X_19332_ _19331_/Y _19327_/X _19221_/X _19327_/X VGND VGND VPWR VPWR _19332_/X sky130_fd_sc_hd__a2bb2o_4
X_13756_ _13724_/X _14697_/A _13754_/X VGND VGND VPWR VPWR _13756_/X sky130_fd_sc_hd__o21a_4
XFILLER_204_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12707_ _12686_/A _12707_/B _12706_/Y VGND VGND VPWR VPWR _25408_/D sky130_fd_sc_hd__and3_4
XFILLER_149_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16475_ _16470_/A VGND VGND VPWR VPWR _16475_/X sky130_fd_sc_hd__buf_2
X_19263_ _23798_/Q VGND VGND VPWR VPWR _21759_/B sky130_fd_sc_hd__inv_2
X_13687_ _11820_/Y _13683_/A _13686_/X _13681_/X VGND VGND VPWR VPWR _13687_/X sky130_fd_sc_hd__o22a_4
XANTENNA__20550__B1 _20600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24532__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15426_ _15425_/X VGND VGND VPWR VPWR _15426_/X sky130_fd_sc_hd__buf_2
X_18214_ _18182_/A _19022_/A VGND VGND VPWR VPWR _18214_/X sky130_fd_sc_hd__or2_4
X_12638_ _12592_/Y _12606_/X _12638_/C _12599_/X VGND VGND VPWR VPWR _12638_/X sky130_fd_sc_hd__or4_4
X_19194_ _18942_/A VGND VGND VPWR VPWR _19194_/X sky130_fd_sc_hd__buf_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23095__A2 _21437_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22137__A _21427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21041__A _15660_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15357_ _15292_/A _15361_/A _15366_/A _15370_/B VGND VGND VPWR VPWR _15357_/X sky130_fd_sc_hd__or4_4
X_18145_ _18113_/A _19446_/A VGND VGND VPWR VPWR _18145_/X sky130_fd_sc_hd__or2_4
X_12569_ _12569_/A VGND VGND VPWR VPWR _12569_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16135__A _22602_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14308_ _25173_/Q _14288_/Y _25172_/Q _14296_/A VGND VGND VPWR VPWR _14308_/X sky130_fd_sc_hd__o22a_4
XFILLER_156_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12791__B1 _12912_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18076_ _18182_/A _19442_/A VGND VGND VPWR VPWR _18076_/X sky130_fd_sc_hd__or2_4
X_15288_ _15288_/A VGND VGND VPWR VPWR _15315_/A sky130_fd_sc_hd__inv_2
X_17027_ _17027_/A VGND VGND VPWR VPWR _17099_/C sky130_fd_sc_hd__inv_2
X_14239_ _14239_/A _14233_/B _15423_/A _14239_/D VGND VGND VPWR VPWR _14239_/X sky130_fd_sc_hd__or4_4
XANTENNA__12177__A2_N _24764_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16809__B1 HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25391__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25320__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18978_ _18974_/Y _18977_/X _17415_/X _18977_/X VGND VGND VPWR VPWR _23898_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_239_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17929_ _24251_/Q _17927_/Y _17917_/B _17928_/X VGND VGND VPWR VPWR _17929_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20940_ _20941_/B VGND VGND VPWR VPWR _20940_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18982__B1 _18981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20871_ _13648_/B VGND VGND VPWR VPWR _20871_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17413__B _14212_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12838__A _12838_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_127_0_HCLK clkbuf_7_63_0_HCLK/X VGND VGND VPWR VPWR _24032_/CLK sky130_fd_sc_hd__clkbuf_1
X_22610_ _17747_/Y _22435_/A _12266_/A _21448_/X VGND VGND VPWR VPWR _22610_/X sky130_fd_sc_hd__o22a_4
XFILLER_198_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11742__A HWDATA[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23590_ _23678_/CLK _19867_/X VGND VGND VPWR VPWR _19866_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_53_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22541_ _22541_/A _22735_/B VGND VGND VPWR VPWR _22541_/X sky130_fd_sc_hd__and2_4
XANTENNA__24273__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25260_ _25260_/CLK _25260_/D HRESETn VGND VGND VPWR VPWR _25260_/Q sky130_fd_sc_hd__dfrtp_4
X_22472_ _22472_/A _22472_/B _22472_/C _22472_/D VGND VGND VPWR VPWR _22472_/X sky130_fd_sc_hd__or4_4
XFILLER_10_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24202__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24211_ _24227_/CLK _24211_/D HRESETn VGND VGND VPWR VPWR _21822_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__21097__A1 _24820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21423_ _21423_/A VGND VGND VPWR VPWR _22298_/A sky130_fd_sc_hd__buf_2
X_25191_ _25230_/CLK _14250_/X HRESETn VGND VGND VPWR VPWR _25191_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16045__A _16038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12782__B1 _12781_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24142_ _24139_/CLK _24142_/D HRESETn VGND VGND VPWR VPWR _24142_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21886__A _22219_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21354_ _14386_/Y _14182_/X _14477_/Y _14245_/A VGND VGND VPWR VPWR _21354_/X sky130_fd_sc_hd__o22a_4
XANTENNA__23162__A1_N _17255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25479__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20305_ _21180_/B _20300_/X _20008_/X _20287_/Y VGND VGND VPWR VPWR _23426_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24073_ _24073_/CLK _24073_/D HRESETn VGND VGND VPWR VPWR _24073_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19356__A _19343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21285_ _21275_/X _21282_/X _21284_/X VGND VGND VPWR VPWR _21285_/X sky130_fd_sc_hd__a21o_4
XFILLER_116_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23024_ _14966_/A _22838_/X _22098_/X _23023_/X VGND VGND VPWR VPWR _23024_/X sky130_fd_sc_hd__a211o_4
XFILLER_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20236_ _13392_/B VGND VGND VPWR VPWR _20236_/Y sky130_fd_sc_hd__inv_2
X_20167_ _21906_/B _20164_/X _20099_/X _20164_/X VGND VGND VPWR VPWR _23479_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25061__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20098_ _23503_/Q VGND VGND VPWR VPWR _21898_/B sky130_fd_sc_hd__inv_2
X_24975_ _24973_/CLK _24975_/D HRESETn VGND VGND VPWR VPWR _24975_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22510__A _16272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11940_ _11940_/A VGND VGND VPWR VPWR _18902_/B sky130_fd_sc_hd__inv_2
X_23926_ _23926_/CLK _23926_/D HRESETn VGND VGND VPWR VPWR _23926_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17604__A _17625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_23_0_HCLK clkbuf_7_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_47_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18973__B1 _17440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_86_0_HCLK clkbuf_7_87_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_86_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11871_ _11851_/X VGND VGND VPWR VPWR _11896_/B sky130_fd_sc_hd__inv_2
X_23857_ _23873_/CLK _23857_/D VGND VGND VPWR VPWR _23857_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_233_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13610_ _13609_/X VGND VGND VPWR VPWR _13610_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11652__A _13807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22808_ _16494_/A _22431_/X _22535_/X VGND VGND VPWR VPWR _22808_/X sky130_fd_sc_hd__o21a_4
X_14590_ _14553_/A _14553_/B VGND VGND VPWR VPWR _14590_/Y sky130_fd_sc_hd__nand2_4
X_23788_ _23754_/CLK _19293_/X VGND VGND VPWR VPWR _23788_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12255__A1_N _12254_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13541_ _13541_/A _13541_/B _13537_/X _13540_/X VGND VGND VPWR VPWR _13575_/A sky130_fd_sc_hd__or4_4
X_25527_ _24947_/CLK _25527_/D HRESETn VGND VGND VPWR VPWR _25527_/Q sky130_fd_sc_hd__dfrtp_4
X_22739_ _22520_/A _22736_/X _22423_/X _22738_/X VGND VGND VPWR VPWR _22740_/A sky130_fd_sc_hd__o22a_4
XFILLER_186_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21875__A3 _22654_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16260_ _16259_/Y _16257_/X _15469_/X _16257_/X VGND VGND VPWR VPWR _24650_/D sky130_fd_sc_hd__a2bb2o_4
X_13472_ _13471_/Y _13469_/X _11775_/X _13469_/X VGND VGND VPWR VPWR _25321_/D sky130_fd_sc_hd__a2bb2o_4
X_25458_ _25382_/CLK _12408_/X HRESETn VGND VGND VPWR VPWR _12172_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_186_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15211_ _15203_/X _15211_/B _15211_/C VGND VGND VPWR VPWR _15211_/X sky130_fd_sc_hd__and3_4
X_12423_ _25454_/Q _12422_/Y VGND VGND VPWR VPWR _12425_/B sky130_fd_sc_hd__or2_4
X_24409_ _23808_/CLK _24409_/D HRESETn VGND VGND VPWR VPWR _20102_/A sky130_fd_sc_hd__dfrtp_4
X_16191_ _16190_/X VGND VGND VPWR VPWR _16191_/X sky130_fd_sc_hd__buf_2
X_25389_ _25387_/CLK _25389_/D HRESETn VGND VGND VPWR VPWR _12895_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19150__B1 _19125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23996__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15142_ _24600_/Q VGND VGND VPWR VPWR _15142_/Y sky130_fd_sc_hd__inv_2
X_12354_ _24840_/Q VGND VGND VPWR VPWR _12354_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21796__A _21484_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23925__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15073_ _25003_/Q VGND VGND VPWR VPWR _15326_/A sky130_fd_sc_hd__inv_2
X_19950_ _23558_/Q VGND VGND VPWR VPWR _21801_/B sky130_fd_sc_hd__inv_2
XANTENNA__19266__A _19253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12285_ _12285_/A VGND VGND VPWR VPWR _12285_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15711__B1 _24885_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14024_ _14023_/X VGND VGND VPWR VPWR _14024_/Y sky130_fd_sc_hd__inv_2
X_18901_ _18901_/A VGND VGND VPWR VPWR _18902_/C sky130_fd_sc_hd__inv_2
X_19881_ _19881_/A VGND VGND VPWR VPWR _22246_/B sky130_fd_sc_hd__inv_2
X_18832_ _16536_/Y _18616_/X _16536_/Y _18616_/X VGND VGND VPWR VPWR _18832_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18763_ _24143_/Q _18763_/B VGND VGND VPWR VPWR _18763_/X sky130_fd_sc_hd__or2_4
X_15975_ _15784_/X _15850_/A _15764_/X _24751_/Q _15925_/X VGND VGND VPWR VPWR _24751_/D
+ sky130_fd_sc_hd__a32o_4
X_17714_ _17711_/Y _18288_/A _17726_/B VGND VGND VPWR VPWR _17714_/X sky130_fd_sc_hd__a21o_4
XFILLER_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16509__A1_N _16507_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14926_ _25037_/Q _24443_/Q _15168_/A _14925_/Y VGND VGND VPWR VPWR _14934_/B sky130_fd_sc_hd__o22a_4
XFILLER_208_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18694_ _18778_/A _18694_/B _18694_/C _18747_/A VGND VGND VPWR VPWR _18695_/B sky130_fd_sc_hd__or4_4
XANTENNA__24784__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17645_ _17647_/A _17645_/B _17645_/C VGND VGND VPWR VPWR _17645_/X sky130_fd_sc_hd__and3_4
X_14857_ _14823_/X _14856_/X _15465_/A _14826_/A VGND VGND VPWR VPWR _14857_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__24713__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13808_ _13807_/X VGND VGND VPWR VPWR _13832_/A sky130_fd_sc_hd__buf_2
XFILLER_90_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14788_ _14788_/A VGND VGND VPWR VPWR _14788_/Y sky130_fd_sc_hd__inv_2
X_17576_ _24302_/Q VGND VGND VPWR VPWR _17577_/C sky130_fd_sc_hd__inv_2
XFILLER_223_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19315_ _18170_/B VGND VGND VPWR VPWR _19315_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13739_ _25279_/Q VGND VGND VPWR VPWR _13739_/Y sky130_fd_sc_hd__inv_2
X_16527_ _16527_/A VGND VGND VPWR VPWR _16527_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19246_ _21607_/B _19245_/X _16882_/X _19245_/X VGND VGND VPWR VPWR _23805_/D sky130_fd_sc_hd__a2bb2o_4
X_16458_ _24576_/Q VGND VGND VPWR VPWR _16458_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14202__B1 _13521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15409_ _15409_/A _15382_/X VGND VGND VPWR VPWR _15418_/A sky130_fd_sc_hd__or2_4
X_16389_ _24603_/Q VGND VGND VPWR VPWR _16389_/Y sky130_fd_sc_hd__inv_2
X_19177_ _19170_/A VGND VGND VPWR VPWR _19177_/X sky130_fd_sc_hd__buf_2
XANTENNA__15950__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18128_ _18128_/A _23830_/Q VGND VGND VPWR VPWR _18130_/B sky130_fd_sc_hd__or2_4
XFILLER_145_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14505__A1 _20601_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18059_ _18097_/A _19190_/A VGND VGND VPWR VPWR _18059_/X sky130_fd_sc_hd__or2_4
XANTENNA__25501__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18080__A _18227_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22579__A1 _16765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21070_ _21014_/B _21048_/Y VGND VGND VPWR VPWR _21070_/X sky130_fd_sc_hd__and2_4
X_20021_ _20020_/Y _20018_/X _19974_/X _20018_/X VGND VGND VPWR VPWR _20021_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18645__A1_N _16589_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24760_ _24763_/CLK _15962_/X HRESETn VGND VGND VPWR VPWR _24760_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21972_ _13763_/X _21972_/B VGND VGND VPWR VPWR _21972_/Y sky130_fd_sc_hd__nand2_4
XFILLER_132_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22751__A1 _21305_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23711_ _23437_/CLK _19511_/X VGND VGND VPWR VPWR _23711_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ _20923_/A VGND VGND VPWR VPWR _20923_/X sky130_fd_sc_hd__buf_2
XPHY_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24691_ _24744_/CLK _24691_/D HRESETn VGND VGND VPWR VPWR _22564_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24454__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ _25326_/CLK _19719_/X VGND VGND VPWR VPWR _23642_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20854_ _20853_/X VGND VGND VPWR VPWR _24041_/D sky130_fd_sc_hd__inv_2
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13244__A1 _11951_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23573_ _23526_/CLK _19913_/X VGND VGND VPWR VPWR _23573_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20785_ _20780_/X _20783_/X _24914_/Q _20784_/X VGND VGND VPWR VPWR _20785_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_168_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25312_ _25492_/CLK _25312_/D HRESETn VGND VGND VPWR VPWR _13492_/A sky130_fd_sc_hd__dfrtp_4
X_22524_ _22287_/X _22522_/X _21122_/X _22523_/X VGND VGND VPWR VPWR _22527_/A sky130_fd_sc_hd__o22a_4
XFILLER_179_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16194__B1 _16001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25243_ _25243_/CLK _13962_/X HRESETn VGND VGND VPWR VPWR scl_oen_o_S5 sky130_fd_sc_hd__dfstp_4
X_22455_ _16515_/Y _22282_/X _16724_/A _16600_/Y _16792_/A VGND VGND VPWR VPWR _22455_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21406_ _22196_/A _21404_/X _21405_/X VGND VGND VPWR VPWR _21406_/X sky130_fd_sc_hd__and3_4
X_25174_ _23884_/CLK _25174_/D HRESETn VGND VGND VPWR VPWR _25174_/Q sky130_fd_sc_hd__dfrtp_4
X_22386_ _22386_/A _22386_/B VGND VGND VPWR VPWR _22386_/X sky130_fd_sc_hd__or2_4
XFILLER_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24125_ _24146_/CLK _18869_/Y HRESETn VGND VGND VPWR VPWR pwm_S7 sky130_fd_sc_hd__dfrtp_4
X_21337_ _21309_/A VGND VGND VPWR VPWR _21337_/X sky130_fd_sc_hd__buf_2
XFILLER_191_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19086__A _19074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12070_ _12069_/Y _12065_/X _11781_/X _12065_/X VGND VGND VPWR VPWR _25482_/D sky130_fd_sc_hd__a2bb2o_4
X_24056_ _24501_/CLK _24056_/D HRESETn VGND VGND VPWR VPWR _24056_/Q sky130_fd_sc_hd__dfrtp_4
X_21268_ _14688_/A _21266_/X _21267_/X VGND VGND VPWR VPWR _21268_/X sky130_fd_sc_hd__and3_4
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23007_ _22983_/X _22987_/X _22991_/Y _23006_/X VGND VGND VPWR VPWR HRDATA[21] sky130_fd_sc_hd__a211o_4
X_20219_ _23458_/Q VGND VGND VPWR VPWR _20219_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19814__A _19805_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21199_ _24213_/Q _21199_/B _21199_/C VGND VGND VPWR VPWR _21199_/X sky130_fd_sc_hd__and3_4
XFILLER_237_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15760_ _12551_/Y _15759_/X _15623_/X _15759_/X VGND VGND VPWR VPWR _15760_/X sky130_fd_sc_hd__a2bb2o_4
X_12972_ _12971_/Y VGND VGND VPWR VPWR _13059_/A sky130_fd_sc_hd__buf_2
X_24958_ _24958_/CLK _15459_/X HRESETn VGND VGND VPWR VPWR _24958_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_64_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11923_ _19620_/A VGND VGND VPWR VPWR _11923_/Y sky130_fd_sc_hd__inv_2
X_14711_ _22228_/A VGND VGND VPWR VPWR _14711_/X sky130_fd_sc_hd__buf_2
X_15691_ _15691_/A VGND VGND VPWR VPWR _15691_/X sky130_fd_sc_hd__buf_2
X_23909_ _23853_/CLK _18949_/X VGND VGND VPWR VPWR _23909_/Q sky130_fd_sc_hd__dfxtp_4
X_24889_ _24889_/CLK _24889_/D HRESETn VGND VGND VPWR VPWR _15675_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24195__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14642_ _17944_/A _14632_/Y VGND VGND VPWR VPWR _14642_/X sky130_fd_sc_hd__or2_4
X_17430_ _21558_/A _17429_/X _16849_/X _17429_/X VGND VGND VPWR VPWR _17430_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11854_ _25519_/Q _11860_/A _11797_/A _11853_/X VGND VGND VPWR VPWR _11854_/X sky130_fd_sc_hd__and4_4
XFILLER_61_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14432__B1 _14407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_110_0_HCLK clkbuf_7_55_0_HCLK/X VGND VGND VPWR VPWR _24035_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ _14563_/A _14563_/B VGND VGND VPWR VPWR _14573_/X sky130_fd_sc_hd__or2_4
X_17361_ _17361_/A VGND VGND VPWR VPWR _24349_/D sky130_fd_sc_hd__inv_2
XANTENNA__15789__A _15783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ _11785_/A VGND VGND VPWR VPWR _15472_/A sky130_fd_sc_hd__buf_2
XPHY_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_173_0_HCLK clkbuf_7_86_0_HCLK/X VGND VGND VPWR VPWR _23844_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19100_ _19100_/A VGND VGND VPWR VPWR _19100_/Y sky130_fd_sc_hd__inv_2
X_13524_ _13630_/A _13520_/Y _13459_/X _13520_/Y VGND VGND VPWR VPWR _25303_/D sky130_fd_sc_hd__a2bb2o_4
X_16312_ _16310_/Y _16306_/X _15948_/X _16311_/X VGND VGND VPWR VPWR _24631_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17292_ _17292_/A _17292_/B VGND VGND VPWR VPWR _17292_/X sky130_fd_sc_hd__or2_4
XFILLER_201_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16243_ _16242_/Y _16239_/X _15965_/X _16239_/X VGND VGND VPWR VPWR _24657_/D sky130_fd_sc_hd__a2bb2o_4
X_19031_ _19030_/Y _19028_/X _18981_/X _19028_/X VGND VGND VPWR VPWR _19031_/X sky130_fd_sc_hd__a2bb2o_4
X_13455_ _21568_/B VGND VGND VPWR VPWR _13482_/B sky130_fd_sc_hd__buf_2
XANTENNA__19123__B1 _19122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12406_ _12172_/A _12405_/Y VGND VGND VPWR VPWR _12406_/X sky130_fd_sc_hd__or2_4
X_16174_ _16174_/A VGND VGND VPWR VPWR _16174_/Y sky130_fd_sc_hd__inv_2
X_13386_ _11951_/A _13370_/X _13385_/X _25329_/Q _13243_/X VGND VGND VPWR VPWR _13386_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_126_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15125_ _24990_/Q VGND VGND VPWR VPWR _15125_/Y sky130_fd_sc_hd__inv_2
X_12337_ _25349_/Q VGND VGND VPWR VPWR _12976_/D sky130_fd_sc_hd__inv_2
XFILLER_115_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15056_ _14880_/Y _15261_/A _15244_/A _15056_/D VGND VGND VPWR VPWR _15056_/X sky130_fd_sc_hd__or4_4
X_19933_ _21665_/B _19932_/X _19617_/X _19932_/X VGND VGND VPWR VPWR _23565_/D sky130_fd_sc_hd__a2bb2o_4
X_12268_ _12268_/A VGND VGND VPWR VPWR _12492_/A sky130_fd_sc_hd__inv_2
X_14007_ _14007_/A _14007_/B _14007_/C _14007_/D VGND VGND VPWR VPWR _14525_/A sky130_fd_sc_hd__or4_4
XFILLER_96_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19864_ _19864_/A VGND VGND VPWR VPWR _19864_/Y sky130_fd_sc_hd__inv_2
X_12199_ _12197_/A _22410_/A _12197_/Y _12198_/Y VGND VGND VPWR VPWR _12199_/X sky130_fd_sc_hd__o22a_4
XFILLER_233_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24965__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18815_ _18815_/A _18815_/B VGND VGND VPWR VPWR _18815_/X sky130_fd_sc_hd__or2_4
X_19795_ _13382_/B VGND VGND VPWR VPWR _19795_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15999__B1 _15996_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22150__A _22150_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13772__A _16721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18746_ _18689_/Y _18691_/B _18767_/B VGND VGND VPWR VPWR _18746_/X sky130_fd_sc_hd__or3_4
XFILLER_237_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15958_ _15958_/A VGND VGND VPWR VPWR _15958_/X sky130_fd_sc_hd__buf_2
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18937__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14909_ _25026_/Q _14908_/A _15219_/A _14908_/Y VGND VGND VPWR VPWR _14909_/X sky130_fd_sc_hd__o22a_4
X_18677_ _18677_/A VGND VGND VPWR VPWR _18730_/A sky130_fd_sc_hd__buf_2
X_15889_ _15889_/A VGND VGND VPWR VPWR _15889_/X sky130_fd_sc_hd__buf_2
XANTENNA__12388__A _12204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17628_ _17559_/Y _17628_/B VGND VGND VPWR VPWR _17637_/B sky130_fd_sc_hd__or2_4
XFILLER_24_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22497__B1 _22493_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17559_ _24714_/Q VGND VGND VPWR VPWR _17559_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14974__B2 _24418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20570_ _20570_/A VGND VGND VPWR VPWR _23942_/D sky130_fd_sc_hd__inv_2
XFILLER_20_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19229_ _19228_/Y _19224_/X _19138_/X _19224_/A VGND VGND VPWR VPWR _19229_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19114__B1 _18998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22240_ _22255_/A _22240_/B VGND VGND VPWR VPWR _22241_/C sky130_fd_sc_hd__or2_4
XFILLER_117_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21867__C _21859_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12273__D _12248_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22171_ _22170_/Y _21349_/A _14117_/Y _14209_/A VGND VGND VPWR VPWR _22171_/X sky130_fd_sc_hd__o22a_4
X_21122_ _22992_/A VGND VGND VPWR VPWR _21122_/X sky130_fd_sc_hd__buf_2
XFILLER_132_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21053_ _22632_/A _21027_/X _21053_/C VGND VGND VPWR VPWR _21288_/A sky130_fd_sc_hd__and3_4
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20004_ _21662_/B _20003_/X _19981_/X _20003_/X VGND VGND VPWR VPWR _20004_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16100__B1 _15567_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23156__A _22145_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22060__A _21627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24635__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24812_ _24804_/CLK _15866_/X HRESETn VGND VGND VPWR VPWR _23187_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18928__B1 _16787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24743_ _24744_/CLK _16005_/X HRESETn VGND VGND VPWR VPWR _24743_/Q sky130_fd_sc_hd__dfrtp_4
X_21955_ _21955_/A VGND VGND VPWR VPWR _21956_/A sky130_fd_sc_hd__buf_2
XFILLER_15_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _24053_/Q VGND VGND VPWR VPWR _20906_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25135__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24674_ _24678_/CLK _24674_/D HRESETn VGND VGND VPWR VPWR _23206_/A sky130_fd_sc_hd__dfrtp_4
X_21886_ _22219_/A _21883_/X _21885_/X VGND VGND VPWR VPWR _21886_/X sky130_fd_sc_hd__and3_4
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16954__A2 _16952_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25198__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23625_ _24413_/CLK _23625_/D VGND VGND VPWR VPWR _19766_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _20837_/A VGND VGND VPWR VPWR _24037_/D sky130_fd_sc_hd__inv_2
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14221__A1_N _14220_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23556_ _25285_/CLK _23556_/D VGND VGND VPWR VPWR _23556_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25494__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_246_0_HCLK clkbuf_8_247_0_HCLK/A VGND VGND VPWR VPWR _24073_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20768_ _13107_/A _20767_/A _13107_/C _20754_/X VGND VGND VPWR VPWR _20768_/X sky130_fd_sc_hd__or4_4
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22507_ _22450_/X _22504_/X _22454_/X _22506_/X VGND VGND VPWR VPWR _22507_/X sky130_fd_sc_hd__o22a_4
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23487_ _23487_/CLK _23487_/D VGND VGND VPWR VPWR _23487_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12561__A2_N _24878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20699_ _20698_/X VGND VGND VPWR VPWR _20699_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ _13169_/A _13240_/B _13239_/X VGND VGND VPWR VPWR _13241_/C sky130_fd_sc_hd__and3_4
X_25226_ _25226_/CLK _25226_/D HRESETn VGND VGND VPWR VPWR _13992_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_7_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22438_ _21448_/X VGND VGND VPWR VPWR _22721_/A sky130_fd_sc_hd__buf_2
XFILLER_108_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13171_ _13168_/A _23458_/Q VGND VGND VPWR VPWR _13171_/X sky130_fd_sc_hd__or2_4
X_25157_ _25158_/CLK _25157_/D HRESETn VGND VGND VPWR VPWR _25157_/Q sky130_fd_sc_hd__dfrtp_4
X_22369_ _22373_/A _22367_/X _22369_/C VGND VGND VPWR VPWR _22369_/X sky130_fd_sc_hd__and3_4
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12122_ _20971_/A VGND VGND VPWR VPWR _12122_/Y sky130_fd_sc_hd__inv_2
X_24108_ _24188_/CLK _12145_/C HRESETn VGND VGND VPWR VPWR _12140_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_123_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25088_ _25089_/CLK _14592_/X HRESETn VGND VGND VPWR VPWR _25088_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_184_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23204__A2 _21292_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17419__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12053_ _12043_/A VGND VGND VPWR VPWR _12081_/A sky130_fd_sc_hd__buf_2
X_16930_ _16131_/Y _17755_/A _16131_/Y _17755_/A VGND VGND VPWR VPWR _16930_/X sky130_fd_sc_hd__a2bb2o_4
X_24039_ _24486_/CLK _20845_/Y HRESETn VGND VGND VPWR VPWR _24039_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16861_ _16859_/Y _16856_/X _16860_/X _16856_/X VGND VGND VPWR VPWR _16861_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24376__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18600_ _16591_/Y _18791_/A _16591_/Y _18791_/A VGND VGND VPWR VPWR _18600_/X sky130_fd_sc_hd__a2bb2o_4
X_15812_ _15810_/X _15789_/X _15735_/X _24836_/Q _15811_/X VGND VGND VPWR VPWR _15812_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17064__A _17381_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24337__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19580_ _19580_/A VGND VGND VPWR VPWR _19580_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16792_ _16792_/A _16792_/B VGND VGND VPWR VPWR _16793_/A sky130_fd_sc_hd__nor2_4
XANTENNA__24305__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18919__B1 _17421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22715__A1 _24869_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18531_ _18442_/Y _18526_/B _18500_/X _18528_/B VGND VGND VPWR VPWR _18531_/X sky130_fd_sc_hd__a211o_4
X_12955_ _12952_/A _12948_/B _12954_/X VGND VGND VPWR VPWR _25373_/D sky130_fd_sc_hd__and3_4
X_15743_ HWDATA[13] VGND VGND VPWR VPWR _15743_/X sky130_fd_sc_hd__buf_2
XFILLER_218_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17999__A _17999_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11906_ _19603_/A VGND VGND VPWR VPWR _11906_/X sky130_fd_sc_hd__buf_2
XFILLER_45_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18462_ _18462_/A _18462_/B VGND VGND VPWR VPWR _18481_/C sky130_fd_sc_hd__or2_4
X_12886_ _12841_/D _12851_/B _12804_/Y VGND VGND VPWR VPWR _12886_/X sky130_fd_sc_hd__o21a_4
X_15674_ _13527_/B VGND VGND VPWR VPWR _15680_/A sky130_fd_sc_hd__buf_2
Xclkbuf_6_56_0_HCLK clkbuf_6_57_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_56_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17412_/X _14212_/B VGND VGND VPWR VPWR _17429_/A sky130_fd_sc_hd__nor2_4
XANTENNA__21314__A _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _13668_/B _24226_/Q _13668_/B _24226_/Q VGND VGND VPWR VPWR _11837_/X sky130_fd_sc_hd__a2bb2o_4
X_14625_ _18082_/A VGND VGND VPWR VPWR _18062_/A sky130_fd_sc_hd__buf_2
X_18393_ _16238_/Y _18473_/A _16238_/Y _18473_/A VGND VGND VPWR VPWR _18393_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__19344__B1 _19301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16408__A _24595_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _13563_/Y _14555_/X VGND VGND VPWR VPWR _14557_/B sky130_fd_sc_hd__or2_4
X_17344_ _17344_/A _17344_/B VGND VGND VPWR VPWR _17345_/B sky130_fd_sc_hd__or2_4
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16158__B1 _15469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _25525_/Q VGND VGND VPWR VPWR _11768_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23940__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ _12013_/B VGND VGND VPWR VPWR _13507_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14487_ _14487_/A VGND VGND VPWR VPWR _14487_/Y sky130_fd_sc_hd__inv_2
X_17275_ _17230_/X _17275_/B _17274_/X VGND VGND VPWR VPWR _17275_/X sky130_fd_sc_hd__and3_4
XFILLER_159_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11699_ _11699_/A VGND VGND VPWR VPWR _11699_/X sky130_fd_sc_hd__buf_2
XFILLER_174_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19014_ _19013_/Y _19011_/X _18942_/X _19011_/X VGND VGND VPWR VPWR _19014_/X sky130_fd_sc_hd__a2bb2o_4
X_13438_ _13438_/A _23787_/Q VGND VGND VPWR VPWR _13438_/X sky130_fd_sc_hd__or2_4
X_16226_ _16226_/A VGND VGND VPWR VPWR _16226_/X sky130_fd_sc_hd__buf_2
XFILLER_173_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22145__A _24617_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16157_ _21698_/A VGND VGND VPWR VPWR _16157_/Y sky130_fd_sc_hd__inv_2
X_13369_ _13369_/A _13365_/X _13369_/C VGND VGND VPWR VPWR _13370_/C sky130_fd_sc_hd__or3_4
XFILLER_155_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17239__A _17239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15108_ _15106_/A _15107_/A _15106_/Y _15107_/Y VGND VGND VPWR VPWR _15108_/X sky130_fd_sc_hd__o22a_4
X_16088_ _24711_/Q VGND VGND VPWR VPWR _16088_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16330__B1 _16236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15039_ _14944_/Y VGND VGND VPWR VPWR _15039_/X sky130_fd_sc_hd__buf_2
X_19916_ _19916_/A VGND VGND VPWR VPWR _21260_/B sky130_fd_sc_hd__inv_2
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14341__C1 _14340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19847_ _19835_/A VGND VGND VPWR VPWR _19847_/X sky130_fd_sc_hd__buf_2
XFILLER_229_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19778_ _23620_/Q VGND VGND VPWR VPWR _19778_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24046__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18729_ _18729_/A _18729_/B VGND VGND VPWR VPWR _18730_/B sky130_fd_sc_hd__or2_4
XFILLER_237_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21740_ _16847_/Y _15704_/A _21582_/A _21739_/X VGND VGND VPWR VPWR _21740_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22965__D _22965_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17594__C1 _17593_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21671_ _21670_/X _21671_/B VGND VGND VPWR VPWR _21671_/X sky130_fd_sc_hd__or2_4
XFILLER_240_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19335__B1 _19200_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23410_ _24302_/CLK _20346_/X VGND VGND VPWR VPWR _20345_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11750__A HWDATA[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20622_ _15468_/Y _20615_/X _20672_/A _20621_/X VGND VGND VPWR VPWR _20623_/A sky130_fd_sc_hd__a211o_4
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24390_ _24390_/CLK _17107_/X HRESETn VGND VGND VPWR VPWR _24390_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21142__B1 _17438_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23341_ _23341_/A VGND VGND VPWR VPWR _23341_/Y sky130_fd_sc_hd__inv_2
X_20553_ _20553_/A _20552_/Y _20553_/C VGND VGND VPWR VPWR _20553_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_13_0_HCLK clkbuf_7_6_0_HCLK/X VGND VGND VPWR VPWR _23415_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_164_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23272_ _23272_/A VGND VGND VPWR VPWR _23272_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_76_0_HCLK clkbuf_8_77_0_HCLK/A VGND VGND VPWR VPWR _24704_/CLK sky130_fd_sc_hd__clkbuf_1
X_20484_ _15451_/A _20515_/B _20479_/B VGND VGND VPWR VPWR _20529_/A sky130_fd_sc_hd__and3_4
X_25011_ _25015_/CLK _15275_/X HRESETn VGND VGND VPWR VPWR _25011_/Q sky130_fd_sc_hd__dfrtp_4
X_22223_ _22223_/A _22221_/X _22222_/X VGND VGND VPWR VPWR _22227_/B sky130_fd_sc_hd__and3_4
XANTENNA__24887__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22154_ _15704_/A _22153_/X _21427_/A _25525_/Q _23138_/A VGND VGND VPWR VPWR _22154_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__21894__A _22386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16321__B1 _16320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24816__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21105_ _21105_/A VGND VGND VPWR VPWR _21105_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22085_ _22365_/A _22085_/B VGND VGND VPWR VPWR _22085_/X sky130_fd_sc_hd__or2_4
XFILLER_120_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22945__A1 _24736_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21036_ _22132_/B VGND VGND VPWR VPWR _21051_/A sky130_fd_sc_hd__buf_2
XFILLER_247_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22987_ _22985_/X _22986_/X _22919_/X VGND VGND VPWR VPWR _22987_/X sky130_fd_sc_hd__or3_4
XFILLER_90_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ _12740_/A VGND VGND VPWR VPWR _12838_/D sky130_fd_sc_hd__inv_2
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17612__A _17625_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21938_ _21933_/X _21937_/X _18301_/A VGND VGND VPWR VPWR _21939_/C sky130_fd_sc_hd__o21a_4
X_24726_ _24266_/CLK _16048_/X HRESETn VGND VGND VPWR VPWR _24726_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16388__B1 _16386_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21134__A _21159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12671_ _12671_/A _12668_/B VGND VGND VPWR VPWR _12671_/Y sky130_fd_sc_hd__nand2_4
X_24657_ _24678_/CLK _24657_/D HRESETn VGND VGND VPWR VPWR _22548_/A sky130_fd_sc_hd__dfrtp_4
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21869_ _21047_/X VGND VGND VPWR VPWR _23075_/C sky130_fd_sc_hd__buf_2
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14938__B2 _14940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _25142_/Q VGND VGND VPWR VPWR _14410_/Y sky130_fd_sc_hd__inv_2
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12949__B1 _12854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23608_ _23610_/CLK _23608_/D VGND VGND VPWR VPWR _23608_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15390_/A _15390_/B VGND VGND VPWR VPWR _15394_/B sky130_fd_sc_hd__or2_4
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24588_ _24985_/CLK _16424_/X HRESETn VGND VGND VPWR VPWR _24588_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _14329_/C _14332_/B _14314_/X _14340_/X VGND VGND VPWR VPWR _14342_/A sky130_fd_sc_hd__a211o_4
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23539_ _24302_/CLK _23539_/D VGND VGND VPWR VPWR _20007_/A sky130_fd_sc_hd__dfxtp_4
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17060_ _16978_/Y _17057_/X VGND VGND VPWR VPWR _17060_/X sky130_fd_sc_hd__or2_4
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _13873_/X _20510_/B _13873_/X _14271_/X VGND VGND VPWR VPWR _14273_/A sky130_fd_sc_hd__o22a_4
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16011_ _24740_/Q VGND VGND VPWR VPWR _16011_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13223_ _13443_/A _13223_/B VGND VGND VPWR VPWR _13223_/X sky130_fd_sc_hd__or2_4
X_25209_ _25056_/CLK _14191_/X HRESETn VGND VGND VPWR VPWR _20503_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_143_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12177__B2 _24764_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_195_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13154_ _13175_/A _23642_/Q VGND VGND VPWR VPWR _13155_/C sky130_fd_sc_hd__or2_4
XANTENNA__16312__B1 _15948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24557__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12105_ _12104_/Y _12102_/X _11781_/X _12102_/X VGND VGND VPWR VPWR _12105_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13085_ _13085_/A _13073_/B _13084_/Y VGND VGND VPWR VPWR _13085_/X sky130_fd_sc_hd__and3_4
X_17962_ _18062_/A _17954_/X _17961_/X _15673_/X _15681_/X VGND VGND VPWR VPWR _17962_/X
+ sky130_fd_sc_hd__o32a_4
X_19701_ _13311_/B VGND VGND VPWR VPWR _19701_/Y sky130_fd_sc_hd__inv_2
X_12036_ _13454_/A VGND VGND VPWR VPWR _16364_/A sky130_fd_sc_hd__buf_2
X_16913_ _16913_/A VGND VGND VPWR VPWR _16913_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17893_ _17893_/A VGND VGND VPWR VPWR _17893_/Y sky130_fd_sc_hd__inv_2
X_19632_ _13270_/B VGND VGND VPWR VPWR _19632_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16844_ _24418_/Q VGND VGND VPWR VPWR _16844_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19563_ _21683_/B _19562_/X _11924_/X _19562_/X VGND VGND VPWR VPWR _19563_/X sky130_fd_sc_hd__a2bb2o_4
X_16775_ _15023_/Y _16774_/X _16522_/X _16774_/X VGND VGND VPWR VPWR _24452_/D sky130_fd_sc_hd__a2bb2o_4
X_13987_ _25236_/Q VGND VGND VPWR VPWR _13987_/X sky130_fd_sc_hd__buf_2
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22164__A2 _21309_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18514_ _18462_/A _18516_/B _18513_/Y VGND VGND VPWR VPWR _18514_/X sky130_fd_sc_hd__o21a_4
XFILLER_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15726_ _15724_/X _15709_/X _15725_/X _24878_/Q _15707_/X VGND VGND VPWR VPWR _15726_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12938_ _12834_/C _12937_/X _12872_/A _12934_/B VGND VGND VPWR VPWR _12939_/A sky130_fd_sc_hd__a211o_4
X_19494_ _19494_/A VGND VGND VPWR VPWR _19494_/X sky130_fd_sc_hd__buf_2
XANTENNA__16379__B1 _16004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16918__A2 _16917_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18445_ _16207_/A _18510_/C _16212_/Y _24178_/Q VGND VGND VPWR VPWR _18445_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15657_ _12083_/A _13800_/B VGND VGND VPWR VPWR _15657_/X sky130_fd_sc_hd__or2_4
XFILLER_22_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25345__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12869_ _12861_/A _12867_/X _12869_/C VGND VGND VPWR VPWR _12869_/X sky130_fd_sc_hd__and3_4
XFILLER_61_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16138__A _22564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14608_ _14608_/A VGND VGND VPWR VPWR _14608_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18376_ _18376_/A VGND VGND VPWR VPWR _18376_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15588_ _15588_/A VGND VGND VPWR VPWR _22878_/A sky130_fd_sc_hd__inv_2
XFILLER_159_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17327_ _17329_/B VGND VGND VPWR VPWR _17327_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14539_ _25099_/Q _14055_/X _14049_/X VGND VGND VPWR VPWR _25099_/D sky130_fd_sc_hd__a21bo_4
XANTENNA__21698__B _23002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17258_ _17191_/Y _17231_/X _17232_/Y _17271_/B VGND VGND VPWR VPWR _17258_/X sky130_fd_sc_hd__or4_4
XANTENNA__16551__B1 _16464_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16209_ _22996_/A VGND VGND VPWR VPWR _16209_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22624__B1 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17189_ _24360_/Q VGND VGND VPWR VPWR _17251_/C sky130_fd_sc_hd__inv_2
XFILLER_161_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24980__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24298__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16601__A HWDATA[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24227__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22910_ _23171_/A VGND VGND VPWR VPWR _22910_/X sky130_fd_sc_hd__buf_2
XANTENNA__19912__A _19900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23890_ _23890_/CLK _23890_/D VGND VGND VPWR VPWR _17932_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_245_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22841_ _21579_/B VGND VGND VPWR VPWR _23263_/C sky130_fd_sc_hd__buf_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22772_ _21424_/X _22771_/X _21427_/X _24871_/Q _21428_/X VGND VGND VPWR VPWR _22773_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16909__A2 _24265_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24511_ _24679_/CLK _24511_/D HRESETn VGND VGND VPWR VPWR _13728_/B sky130_fd_sc_hd__dfrtp_4
X_21723_ _21723_/A VGND VGND VPWR VPWR _21723_/Y sky130_fd_sc_hd__inv_2
X_25491_ _25466_/CLK _25491_/D HRESETn VGND VGND VPWR VPWR _12024_/A sky130_fd_sc_hd__dfrtp_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25086__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24442_ _24443_/CLK _24442_/D HRESETn VGND VGND VPWR VPWR _14962_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21654_ _21654_/A _19493_/Y VGND VGND VPWR VPWR _21654_/X sky130_fd_sc_hd__or2_4
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25015__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16790__B1 _16716_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_200_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20605_ _20605_/A VGND VGND VPWR VPWR _20605_/Y sky130_fd_sc_hd__inv_2
X_24373_ _24377_/CLK _24373_/D HRESETn VGND VGND VPWR VPWR _17040_/A sky130_fd_sc_hd__dfrtp_4
X_21585_ _16615_/Y _21581_/X _21582_/X _21584_/X VGND VGND VPWR VPWR _21585_/X sky130_fd_sc_hd__o22a_4
XFILLER_166_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23324_ _23324_/A _16792_/A VGND VGND VPWR VPWR _23324_/Y sky130_fd_sc_hd__nor2_4
XFILLER_165_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20536_ _20495_/C _20478_/Y _20492_/X _20535_/X VGND VGND VPWR VPWR _24073_/D sky130_fd_sc_hd__a211o_4
XFILLER_138_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23255_ _22141_/X _23252_/X _23254_/X VGND VGND VPWR VPWR _23274_/B sky130_fd_sc_hd__and3_4
XFILLER_192_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20467_ _20467_/A _20463_/B _20467_/C _20466_/X VGND VGND VPWR VPWR _20523_/A sky130_fd_sc_hd__and4_4
XFILLER_181_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22206_ _22209_/A _20140_/Y VGND VGND VPWR VPWR _22208_/B sky130_fd_sc_hd__or2_4
X_23186_ _23103_/A _23185_/X VGND VGND VPWR VPWR _23186_/X sky130_fd_sc_hd__and2_4
X_20398_ _13331_/B VGND VGND VPWR VPWR _20398_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24650__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22137_ _21427_/A VGND VGND VPWR VPWR _22138_/C sky130_fd_sc_hd__buf_2
X_22068_ _22373_/A _22066_/X _22068_/C VGND VGND VPWR VPWR _22068_/X sky130_fd_sc_hd__and3_4
XFILLER_247_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12331__B2 _24825_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13910_ _24975_/Q VGND VGND VPWR VPWR _13944_/A sky130_fd_sc_hd__inv_2
X_21019_ _15697_/B VGND VGND VPWR VPWR _21019_/X sky130_fd_sc_hd__buf_2
XFILLER_236_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14890_ _15192_/A _16806_/A _14888_/Y _16806_/A VGND VGND VPWR VPWR _14891_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15473__A1_N _14863_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13841_ _23995_/Q VGND VGND VPWR VPWR _13841_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_121_0_HCLK clkbuf_6_60_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_243_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13772_ _16721_/A _16721_/B _13772_/C _13772_/D VGND VGND VPWR VPWR _13772_/X sky130_fd_sc_hd__and4_4
X_16560_ _16548_/A VGND VGND VPWR VPWR _16560_/X sky130_fd_sc_hd__buf_2
X_15511_ _15511_/A VGND VGND VPWR VPWR _15530_/A sky130_fd_sc_hd__buf_2
X_12723_ _12716_/B VGND VGND VPWR VPWR _12724_/B sky130_fd_sc_hd__inv_2
X_24709_ _24704_/CLK _24709_/D HRESETn VGND VGND VPWR VPWR _23225_/A sky130_fd_sc_hd__dfrtp_4
X_16491_ _16490_/Y _16488_/X _16400_/X _16488_/X VGND VGND VPWR VPWR _24565_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_230_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18230_ _17966_/A _18229_/X _24242_/Q _18024_/A VGND VGND VPWR VPWR _24242_/D sky130_fd_sc_hd__o22a_4
XFILLER_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12654_ _12598_/X _12662_/B VGND VGND VPWR VPWR _12655_/B sky130_fd_sc_hd__or2_4
X_15442_ _13930_/A _15432_/X _15441_/X _13931_/B _15439_/X VGND VGND VPWR VPWR _15442_/X
+ sky130_fd_sc_hd__a32o_4
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18161_ _18097_/A _18161_/B VGND VGND VPWR VPWR _18161_/X sky130_fd_sc_hd__or2_4
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12693_/A _24861_/Q _12584_/X _24858_/Q VGND VGND VPWR VPWR _12586_/D sky130_fd_sc_hd__a2bb2o_4
X_15373_ _15281_/A VGND VGND VPWR VPWR _15379_/A sky130_fd_sc_hd__buf_2
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17112_ _17105_/A _17099_/D _17111_/X VGND VGND VPWR VPWR _17112_/X sky130_fd_sc_hd__and3_4
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14324_ _18372_/B _14324_/B VGND VGND VPWR VPWR _14332_/B sky130_fd_sc_hd__or2_4
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18092_ _18125_/A _19128_/A VGND VGND VPWR VPWR _18094_/B sky130_fd_sc_hd__or2_4
XANTENNA__16533__B1 _16435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24738__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14255_ _14254_/Y _14252_/X _13785_/X _14252_/X VGND VGND VPWR VPWR _14255_/X sky130_fd_sc_hd__a2bb2o_4
X_17043_ _17120_/A _17043_/B _17042_/X VGND VGND VPWR VPWR _17088_/B sky130_fd_sc_hd__or3_4
XFILLER_184_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13206_ _13363_/A _13206_/B VGND VGND VPWR VPWR _13209_/B sky130_fd_sc_hd__or2_4
XFILLER_125_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14186_ _20667_/A VGND VGND VPWR VPWR _20628_/A sky130_fd_sc_hd__inv_2
XANTENNA__24391__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22423__A _22423_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13137_ _13170_/A _23666_/Q VGND VGND VPWR VPWR _13137_/X sky130_fd_sc_hd__or2_4
XFILLER_151_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18994_ _18992_/Y _18993_/X _18948_/X _18993_/X VGND VGND VPWR VPWR _23893_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24320__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13068_ _13097_/A _12321_/Y _13068_/C _13068_/D VGND VGND VPWR VPWR _13069_/B sky130_fd_sc_hd__or4_4
X_17945_ _17950_/A _17945_/B _17945_/C VGND VGND VPWR VPWR _17945_/X sky130_fd_sc_hd__and3_4
XFILLER_112_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21039__A _21038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12019_ _12019_/A VGND VGND VPWR VPWR _12019_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17876_ _16925_/A _17876_/B VGND VGND VPWR VPWR _17877_/C sky130_fd_sc_hd__or2_4
XFILLER_241_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19615_ _23677_/Q VGND VGND VPWR VPWR _21684_/B sky130_fd_sc_hd__inv_2
X_16827_ _16841_/A VGND VGND VPWR VPWR _16827_/X sky130_fd_sc_hd__buf_2
XFILLER_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25526__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23334__A1 _24477_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19546_ _19545_/Y _19539_/X _19408_/X _19526_/A VGND VGND VPWR VPWR _23699_/D sky130_fd_sc_hd__a2bb2o_4
X_16758_ _16757_/Y _16755_/X _15739_/X _16755_/X VGND VGND VPWR VPWR _24461_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15709_ _15700_/X VGND VGND VPWR VPWR _15709_/X sky130_fd_sc_hd__buf_2
XFILLER_62_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19477_ _19477_/A VGND VGND VPWR VPWR _22336_/B sky130_fd_sc_hd__inv_2
X_16689_ _16689_/A VGND VGND VPWR VPWR _16689_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15024__B1 _25014_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_26_0_HCLK clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_26_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18428_ _18595_/A VGND VGND VPWR VPWR _18561_/C sky130_fd_sc_hd__inv_2
XFILLER_22_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18359_ _18350_/A _17480_/X _18358_/X VGND VGND VPWR VPWR _18359_/X sky130_fd_sc_hd__a21o_4
XFILLER_148_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22845__B1 _22835_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21370_ _21155_/B VGND VGND VPWR VPWR _21721_/B sky130_fd_sc_hd__buf_2
XFILLER_175_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24479__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20321_ _20320_/Y _20316_/X _20061_/X _20316_/X VGND VGND VPWR VPWR _20321_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24408__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23040_ _22638_/B VGND VGND VPWR VPWR _23040_/X sky130_fd_sc_hd__buf_2
X_20252_ _20252_/A VGND VGND VPWR VPWR _21775_/B sky130_fd_sc_hd__inv_2
XANTENNA__23270__B1 _17517_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12561__B2 _24878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20183_ _22225_/B _20180_/X _20092_/X _20180_/X VGND VGND VPWR VPWR _23473_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24061__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24991_ _25005_/CLK _24991_/D HRESETn VGND VGND VPWR VPWR _15369_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23942_ _25140_/CLK _23942_/D HRESETn VGND VGND VPWR VPWR _18876_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_97_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23873_ _23873_/CLK _23873_/D VGND VGND VPWR VPWR _23873_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23325__A1 _22468_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19529__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22824_ _21289_/X VGND VGND VPWR VPWR _22824_/X sky130_fd_sc_hd__buf_2
XFILLER_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22755_ _15595_/Y _15981_/A VGND VGND VPWR VPWR _22755_/X sky130_fd_sc_hd__and2_4
X_25543_ _25538_/CLK _11693_/X HRESETn VGND VGND VPWR VPWR _11690_/A sky130_fd_sc_hd__dfrtp_4
X_21706_ _21706_/A VGND VGND VPWR VPWR _21706_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25474_ _25474_/CLK _12100_/X HRESETn VGND VGND VPWR VPWR _25474_/Q sky130_fd_sc_hd__dfrtp_4
X_22686_ _22686_/A _22686_/B VGND VGND VPWR VPWR _22686_/Y sky130_fd_sc_hd__nor2_4
XFILLER_240_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22508__A _21587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24425_ _24419_/CLK _24425_/D HRESETn VGND VGND VPWR VPWR _24425_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21412__A _22202_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21637_ _21756_/A _21637_/B VGND VGND VPWR VPWR _21638_/C sky130_fd_sc_hd__or2_4
XFILLER_100_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12370_ _12370_/A _12370_/B VGND VGND VPWR VPWR _12370_/X sky130_fd_sc_hd__or2_4
X_24356_ _24341_/CLK _17330_/X HRESETn VGND VGND VPWR VPWR _24356_/Q sky130_fd_sc_hd__dfrtp_4
X_21568_ _21568_/A _21568_/B VGND VGND VPWR VPWR _21569_/A sky130_fd_sc_hd__or2_4
XFILLER_166_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24831__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22851__A3 _15855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23307_ _23307_/A _22658_/B VGND VGND VPWR VPWR _23307_/X sky130_fd_sc_hd__or2_4
X_20519_ _20519_/A _20518_/X VGND VGND VPWR VPWR _24077_/D sky130_fd_sc_hd__or2_4
X_24287_ _24275_/CLK _17782_/X HRESETn VGND VGND VPWR VPWR _16913_/A sky130_fd_sc_hd__dfrtp_4
X_21499_ _17731_/X _21490_/X _21498_/X VGND VGND VPWR VPWR _21499_/X sky130_fd_sc_hd__or3_4
XANTENNA__16771__A1_N _15003_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24149__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_46_0_HCLK clkbuf_7_47_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_46_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14040_ _14059_/A _14532_/C _14040_/C _14039_/X VGND VGND VPWR VPWR _14041_/B sky130_fd_sc_hd__or4_4
X_23238_ _23238_/A _23063_/X VGND VGND VPWR VPWR _23238_/X sky130_fd_sc_hd__or2_4
XFILLER_125_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23169_ _23169_/A _23169_/B VGND VGND VPWR VPWR _23169_/Y sky130_fd_sc_hd__nor2_4
XFILLER_106_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16156__A1_N _16154_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13584__B _14422_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15991_ HWDATA[31] VGND VGND VPWR VPWR _15991_/X sky130_fd_sc_hd__buf_2
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17730_ _18314_/A VGND VGND VPWR VPWR _17730_/X sky130_fd_sc_hd__buf_2
X_14942_ _25020_/Q VGND VGND VPWR VPWR _14942_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17661_ _17682_/A _17661_/B _17661_/C VGND VGND VPWR VPWR _24304_/D sky130_fd_sc_hd__and3_4
XFILLER_235_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14873_ _14871_/Y _14805_/X _14830_/X _14872_/Y VGND VGND VPWR VPWR _14874_/A sky130_fd_sc_hd__o22a_4
XFILLER_208_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19400_ _18110_/B VGND VGND VPWR VPWR _19400_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16612_ _16610_/Y _16606_/X _16349_/X _16611_/X VGND VGND VPWR VPWR _24519_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17072__A _17381_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13824_ _11760_/X VGND VGND VPWR VPWR _13824_/X sky130_fd_sc_hd__buf_2
XFILLER_91_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12068__B1 _11775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17592_ _17627_/A VGND VGND VPWR VPWR _17625_/A sky130_fd_sc_hd__inv_2
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12928__B _12588_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19331_ _18121_/B VGND VGND VPWR VPWR _19331_/Y sky130_fd_sc_hd__inv_2
X_16543_ _16538_/Y _16542_/X _15545_/X _16542_/X VGND VGND VPWR VPWR _24546_/D sky130_fd_sc_hd__a2bb2o_4
X_13755_ _13753_/X _13754_/X _13753_/X _13754_/X VGND VGND VPWR VPWR _13755_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ _12706_/A _12693_/X VGND VGND VPWR VPWR _12706_/Y sky130_fd_sc_hd__nand2_4
X_19262_ _19261_/Y _19259_/X _16873_/X _19259_/X VGND VGND VPWR VPWR _19262_/X sky130_fd_sc_hd__a2bb2o_4
X_16474_ _24571_/Q VGND VGND VPWR VPWR _16474_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13686_ _13686_/A _13686_/B VGND VGND VPWR VPWR _13686_/X sky130_fd_sc_hd__or2_4
XFILLER_189_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24919__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18213_ _13617_/X _18205_/X _18212_/X VGND VGND VPWR VPWR _18213_/X sky130_fd_sc_hd__and3_4
X_15425_ _23993_/Q _23967_/Q _14236_/D _15430_/A VGND VGND VPWR VPWR _15425_/X sky130_fd_sc_hd__o22a_4
X_12637_ _12636_/X VGND VGND VPWR VPWR _25427_/D sky130_fd_sc_hd__inv_2
X_19193_ _23823_/Q VGND VGND VPWR VPWR _19193_/Y sky130_fd_sc_hd__inv_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23095__A3 _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18144_ _14636_/A _18144_/B _18143_/X VGND VGND VPWR VPWR _18144_/X sky130_fd_sc_hd__and3_4
X_12568_ _12638_/C _24877_/Q _25411_/Q _12511_/Y VGND VGND VPWR VPWR _12568_/X sky130_fd_sc_hd__a2bb2o_4
X_15356_ _15356_/A _15355_/X VGND VGND VPWR VPWR _15370_/B sky130_fd_sc_hd__or2_4
XANTENNA__16506__B1 _16236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24572__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14307_ _14295_/A _14306_/X _25320_/Q _14300_/X VGND VGND VPWR VPWR _25174_/D sky130_fd_sc_hd__o22a_4
XFILLER_8_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12791__B2 _22714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18075_ _17984_/X _18073_/X _18075_/C VGND VGND VPWR VPWR _18075_/X sky130_fd_sc_hd__and3_4
XFILLER_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12499_ _12498_/Y _24866_/Q _12498_/Y _24866_/Q VGND VGND VPWR VPWR _12507_/A sky130_fd_sc_hd__a2bb2o_4
X_15287_ _15331_/A VGND VGND VPWR VPWR _15323_/A sky130_fd_sc_hd__buf_2
XFILLER_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24501__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17026_ _17026_/A _16973_/Y VGND VGND VPWR VPWR _17026_/X sky130_fd_sc_hd__or2_4
XANTENNA__18259__B1 _16849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14238_ _14238_/A _13939_/B _13948_/Y VGND VGND VPWR VPWR _14239_/D sky130_fd_sc_hd__or3_4
XANTENNA__23249__A _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22153__A _22153_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14169_ _14169_/A VGND VGND VPWR VPWR _14169_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_3_0_HCLK clkbuf_6_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_7_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_112_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18977_ _18986_/A VGND VGND VPWR VPWR _18977_/X sky130_fd_sc_hd__buf_2
XFILLER_239_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17928_ _17921_/Y _17926_/A _15905_/X VGND VGND VPWR VPWR _17928_/X sky130_fd_sc_hd__o21a_4
XFILLER_79_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17859_ _16915_/Y _17849_/X _17862_/B VGND VGND VPWR VPWR _17859_/X sky130_fd_sc_hd__or3_4
XANTENNA__25360__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20870_ _20919_/A VGND VGND VPWR VPWR _20870_/X sky130_fd_sc_hd__buf_2
XFILLER_199_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16993__B1 _16042_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12838__B _12838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19529_ _19528_/Y _19526_/X _19392_/X _19526_/X VGND VGND VPWR VPWR _23705_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22540_ _22540_/A _21642_/X VGND VGND VPWR VPWR _22540_/X sky130_fd_sc_hd__and2_4
XFILLER_201_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15548__A1 _15540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18860__A1_N _24568_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22471_ _22469_/X _22470_/X VGND VGND VPWR VPWR _22472_/D sky130_fd_sc_hd__nor2_4
X_24210_ _23912_/CLK _18332_/Y HRESETn VGND VGND VPWR VPWR _17452_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21422_ _21021_/A VGND VGND VPWR VPWR _21423_/A sky130_fd_sc_hd__buf_2
X_25190_ _25249_/CLK _14253_/X HRESETn VGND VGND VPWR VPWR _14251_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__12231__B1 _12418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21097__A2 _21082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24141_ _24340_/CLK _18771_/X HRESETn VGND VGND VPWR VPWR _18689_/A sky130_fd_sc_hd__dfrtp_4
X_21353_ _21353_/A VGND VGND VPWR VPWR _21356_/C sky130_fd_sc_hd__inv_2
XFILLER_107_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24242__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20304_ _20304_/A VGND VGND VPWR VPWR _21180_/B sky130_fd_sc_hd__inv_2
X_24072_ _24073_/CLK _24072_/D HRESETn VGND VGND VPWR VPWR _24072_/Q sky130_fd_sc_hd__dfrtp_4
X_21284_ _22515_/A VGND VGND VPWR VPWR _21284_/X sky130_fd_sc_hd__buf_2
XANTENNA__15720__A1 _15540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22063__A _22365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23023_ _16743_/A _23263_/B _23263_/C VGND VGND VPWR VPWR _23023_/X sky130_fd_sc_hd__and3_4
X_20235_ _20233_/Y _20234_/X _20061_/X _20234_/X VGND VGND VPWR VPWR _23453_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16061__A _24721_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20166_ _23479_/Q VGND VGND VPWR VPWR _21906_/B sky130_fd_sc_hd__inv_2
XANTENNA__25448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20097_ _22072_/B _20088_/X _20095_/X _20096_/X VGND VGND VPWR VPWR _20097_/X sky130_fd_sc_hd__a2bb2o_4
X_24974_ _24973_/CLK _15434_/X HRESETn VGND VGND VPWR VPWR _24974_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_217_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22510__B _22509_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23925_ _25113_/CLK _25113_/Q HRESETn VGND VGND VPWR VPWR _22317_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_242_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11870_ _11796_/B _11869_/Y _11864_/X VGND VGND VPWR VPWR _11870_/X sky130_fd_sc_hd__o21a_4
XANTENNA__25030__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23856_ _23873_/CLK _19102_/X VGND VGND VPWR VPWR _19100_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_217_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22807_ _22807_/A VGND VGND VPWR VPWR _22807_/X sky130_fd_sc_hd__buf_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20999_ _14817_/X _20998_/X _21006_/B VGND VGND VPWR VPWR _23994_/D sky130_fd_sc_hd__o21a_4
X_23787_ _23464_/CLK _19296_/X VGND VGND VPWR VPWR _23787_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13540_ _13538_/Y _13535_/A _25256_/Q _14549_/A VGND VGND VPWR VPWR _13540_/X sky130_fd_sc_hd__a2bb2o_4
X_25526_ _25524_/CLK _25526_/D HRESETn VGND VGND VPWR VPWR _25526_/Q sky130_fd_sc_hd__dfrtp_4
X_22738_ _17329_/A _22429_/X _22737_/Y VGND VGND VPWR VPWR _22738_/X sky130_fd_sc_hd__o21a_4
XFILLER_13_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16736__B1 _16382_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13471_ _25321_/Q VGND VGND VPWR VPWR _13471_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22669_ _22669_/A _22669_/B _22668_/X _22725_/A VGND VGND VPWR VPWR _22670_/A sky130_fd_sc_hd__and4_4
X_25457_ _25453_/CLK _12410_/Y HRESETn VGND VGND VPWR VPWR _25457_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_187_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16236__A _16236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12422_ _12422_/A VGND VGND VPWR VPWR _12422_/Y sky130_fd_sc_hd__inv_2
X_15210_ _15210_/A _15207_/X VGND VGND VPWR VPWR _15211_/C sky130_fd_sc_hd__or2_4
XFILLER_201_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24408_ _23378_/CLK _24408_/D HRESETn VGND VGND VPWR VPWR _16875_/A sky130_fd_sc_hd__dfrtp_4
X_16190_ _16183_/Y VGND VGND VPWR VPWR _16190_/X sky130_fd_sc_hd__buf_2
X_25388_ _25387_/CLK _12899_/Y HRESETn VGND VGND VPWR VPWR _25388_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12353_ _13069_/A _24824_/Q _25363_/Q _12352_/Y VGND VGND VPWR VPWR _12359_/B sky130_fd_sc_hd__a2bb2o_4
X_15141_ _15139_/Y _24584_/Q _15288_/A _15140_/Y VGND VGND VPWR VPWR _15141_/X sky130_fd_sc_hd__a2bb2o_4
X_24339_ _24340_/CLK _17403_/X HRESETn VGND VGND VPWR VPWR _24339_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_127_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15072_ _15072_/A VGND VGND VPWR VPWR _15072_/Y sky130_fd_sc_hd__inv_2
X_12284_ _24826_/Q VGND VGND VPWR VPWR _12284_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15711__A1 _15540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14023_ _14021_/Y _13975_/A _14034_/A _14014_/D VGND VGND VPWR VPWR _14023_/X sky130_fd_sc_hd__or4_4
X_18900_ _18900_/A _11948_/A VGND VGND VPWR VPWR _18900_/X sky130_fd_sc_hd__and2_4
XFILLER_141_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12525__B2 _12524_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19880_ _19876_/Y _19879_/X _19600_/X _19879_/X VGND VGND VPWR VPWR _19880_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18831_ _16472_/Y _18732_/A _16472_/Y _18732_/A VGND VGND VPWR VPWR _18835_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23965__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_133_0_HCLK clkbuf_7_66_0_HCLK/X VGND VGND VPWR VPWR _23912_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20063__A3 _14262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_196_0_HCLK clkbuf_7_98_0_HCLK/X VGND VGND VPWR VPWR _24037_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_121_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19282__A _18985_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18762_ _18758_/X VGND VGND VPWR VPWR _18763_/B sky130_fd_sc_hd__inv_2
X_15974_ _15784_/X _15850_/A _15830_/X _24752_/Q _15925_/X VGND VGND VPWR VPWR _24752_/D
+ sky130_fd_sc_hd__a32o_4
XANTENNA__25118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22420__B _22420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17713_ _24217_/Q _19455_/B VGND VGND VPWR VPWR _17726_/B sky130_fd_sc_hd__and2_4
X_14925_ _24443_/Q VGND VGND VPWR VPWR _14925_/Y sky130_fd_sc_hd__inv_2
X_18693_ _18760_/A _18755_/B _18693_/C _18692_/Y VGND VGND VPWR VPWR _18747_/A sky130_fd_sc_hd__or4_4
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17644_ _17523_/Y _17647_/B VGND VGND VPWR VPWR _17645_/C sky130_fd_sc_hd__nand2_4
X_14856_ _14808_/C _14808_/B _14808_/C _14808_/B VGND VGND VPWR VPWR _14856_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13807_ _13807_/A _13807_/B _13807_/C _13807_/D VGND VGND VPWR VPWR _13807_/X sky130_fd_sc_hd__and4_4
XANTENNA__13789__B1 _13788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17575_ _24294_/Q VGND VGND VPWR VPWR _17575_/Y sky130_fd_sc_hd__inv_2
X_14787_ _14787_/A _13609_/X _14783_/X _14787_/D VGND VGND VPWR VPWR _14788_/A sky130_fd_sc_hd__or4_4
X_11999_ _11976_/Y _11983_/B _11983_/Y _11998_/X VGND VGND VPWR VPWR _12012_/A sky130_fd_sc_hd__a211o_4
X_19314_ _19312_/Y _19313_/X _19200_/X _19313_/X VGND VGND VPWR VPWR _23781_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22512__A2 _22992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16526_ _16524_/Y _16521_/X _16525_/X _16521_/X VGND VGND VPWR VPWR _16526_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13738_ _25280_/Q VGND VGND VPWR VPWR _20157_/C sky130_fd_sc_hd__buf_2
XFILLER_220_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16727__B1 _15545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24753__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19245_ _19232_/Y VGND VGND VPWR VPWR _19245_/X sky130_fd_sc_hd__buf_2
X_16457_ _16456_/Y _16454_/X _16373_/X _16454_/X VGND VGND VPWR VPWR _24577_/D sky130_fd_sc_hd__a2bb2o_4
X_13669_ _13669_/A _13668_/X VGND VGND VPWR VPWR _13669_/X sky130_fd_sc_hd__or2_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15408_ _15407_/X VGND VGND VPWR VPWR _24980_/D sky130_fd_sc_hd__inv_2
X_19176_ _23829_/Q VGND VGND VPWR VPWR _19176_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16678__A1_N _16677_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12213__B1 _12211_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16388_ _15097_/Y _16381_/X _16386_/X _16387_/X VGND VGND VPWR VPWR _24604_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18127_ _18094_/A _18127_/B _18127_/C VGND VGND VPWR VPWR _18131_/B sky130_fd_sc_hd__and3_4
XANTENNA__15985__A _16366_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15339_ _15339_/A VGND VGND VPWR VPWR _15340_/B sky130_fd_sc_hd__inv_2
XFILLER_8_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19457__A _19456_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18058_ _18128_/A _19169_/A VGND VGND VPWR VPWR _18060_/B sky130_fd_sc_hd__or2_4
X_17009_ _16067_/Y _17036_/A _24717_/Q _17041_/C VGND VGND VPWR VPWR _17009_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_92_0_HCLK clkbuf_7_93_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_92_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_20020_ _20020_/A VGND VGND VPWR VPWR _20020_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25541__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17705__A _17704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21971_ _21649_/X _21958_/X _21962_/Y _13772_/D _21970_/X VGND VGND VPWR VPWR _21972_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__20211__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11753__A HWDATA[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20922_ _20920_/Y _20916_/X _20921_/X VGND VGND VPWR VPWR _20922_/X sky130_fd_sc_hd__o21a_4
X_23710_ _23437_/CLK _19513_/X VGND VGND VPWR VPWR _23710_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14767__C _14764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24690_ _24744_/CLK _16143_/X HRESETn VGND VGND VPWR VPWR _22494_/A sky130_fd_sc_hd__dfrtp_4
XPHY_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16966__B1 _24743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20853_ _16701_/Y _20846_/X _20834_/X _20852_/Y VGND VGND VPWR VPWR _20853_/X sky130_fd_sc_hd__o22a_4
X_23641_ _25326_/CLK _23641_/D VGND VGND VPWR VPWR _13235_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23572_ _23525_/CLK _19915_/X VGND VGND VPWR VPWR _19914_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20784_ _20784_/A VGND VGND VPWR VPWR _20784_/X sky130_fd_sc_hd__buf_2
XFILLER_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22058__A _22386_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19558__A1_N _21950_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21711__B1 _24261_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24494__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22523_ _15610_/Y _22523_/B VGND VGND VPWR VPWR _22523_/X sky130_fd_sc_hd__and2_4
X_25311_ _25466_/CLK _13495_/X HRESETn VGND VGND VPWR VPWR _25311_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24423__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22454_ _16180_/X VGND VGND VPWR VPWR _22454_/X sky130_fd_sc_hd__buf_2
X_25242_ _25238_/CLK _14050_/Y HRESETn VGND VGND VPWR VPWR _25242_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21405_ _21385_/X _21405_/B VGND VGND VPWR VPWR _21405_/X sky130_fd_sc_hd__or2_4
X_25173_ _25479_/CLK _25173_/D HRESETn VGND VGND VPWR VPWR _25173_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22385_ _22385_/A _20135_/Y VGND VGND VPWR VPWR _22385_/X sky130_fd_sc_hd__or2_4
XFILLER_157_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24124_ _23951_/CLK _18889_/X HRESETn VGND VGND VPWR VPWR _20984_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__22505__B _22505_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21336_ _21232_/X VGND VGND VPWR VPWR _21336_/X sky130_fd_sc_hd__buf_2
XFILLER_136_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24055_ _24501_/CLK _24055_/D HRESETn VGND VGND VPWR VPWR _24055_/Q sky130_fd_sc_hd__dfrtp_4
X_21267_ _21250_/A _20050_/Y VGND VGND VPWR VPWR _21267_/X sky130_fd_sc_hd__or2_4
XFILLER_135_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23006_ _23072_/A _22994_/Y _23006_/C _23006_/D VGND VGND VPWR VPWR _23006_/X sky130_fd_sc_hd__or4_4
XFILLER_150_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20218_ _20217_/Y _20213_/X _19759_/X _20200_/Y VGND VGND VPWR VPWR _20218_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21198_ _21189_/A _20283_/Y VGND VGND VPWR VPWR _21199_/C sky130_fd_sc_hd__or2_4
XFILLER_103_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_206_0_HCLK clkbuf_8_206_0_HCLK/A VGND VGND VPWR VPWR _24551_/CLK sky130_fd_sc_hd__clkbuf_1
X_20149_ _23485_/Q VGND VGND VPWR VPWR _21623_/B sky130_fd_sc_hd__inv_2
XFILLER_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25211__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12971_ _24781_/Q VGND VGND VPWR VPWR _12971_/Y sky130_fd_sc_hd__inv_2
X_24957_ _24958_/CLK _15461_/X HRESETn VGND VGND VPWR VPWR _24957_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_85_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12791__A2_N _22714_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20202__B1 _18250_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14710_ _14710_/A VGND VGND VPWR VPWR _22228_/A sky130_fd_sc_hd__buf_2
X_11922_ _19984_/A VGND VGND VPWR VPWR _19620_/A sky130_fd_sc_hd__buf_2
X_23908_ _23853_/CLK _18952_/X VGND VGND VPWR VPWR _23908_/Q sky130_fd_sc_hd__dfxtp_4
X_15690_ _15690_/A VGND VGND VPWR VPWR _15691_/A sky130_fd_sc_hd__buf_2
X_24888_ _23767_/CLK _15693_/X HRESETn VGND VGND VPWR VPWR _24888_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_205_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14641_ _17949_/A VGND VGND VPWR VPWR _17944_/A sky130_fd_sc_hd__buf_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11853_ _11852_/Y VGND VGND VPWR VPWR _11853_/X sky130_fd_sc_hd__buf_2
X_23839_ _23846_/CLK _19152_/X VGND VGND VPWR VPWR _23839_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _17352_/B _17352_/C _17284_/X _17357_/B VGND VGND VPWR VPWR _17361_/A sky130_fd_sc_hd__a211o_4
XFILLER_198_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ HWDATA[2] VGND VGND VPWR VPWR _11785_/A sky130_fd_sc_hd__buf_2
X_14572_ _14570_/X _14546_/X _14571_/X _13758_/X _14563_/C VGND VGND VPWR VPWR _25096_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21702__B1 _24858_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ _16284_/X VGND VGND VPWR VPWR _16311_/X sky130_fd_sc_hd__buf_2
XFILLER_201_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ _13523_/A VGND VGND VPWR VPWR _13630_/A sky130_fd_sc_hd__inv_2
X_25509_ _25510_/CLK _11903_/X HRESETn VGND VGND VPWR VPWR _19967_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_158_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17291_ _17290_/X VGND VGND VPWR VPWR _17292_/B sky130_fd_sc_hd__inv_2
XANTENNA__24164__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19030_ _18002_/B VGND VGND VPWR VPWR _19030_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16242_ _22548_/A VGND VGND VPWR VPWR _16242_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13454_ _13454_/A _14365_/B _11660_/A _12039_/D VGND VGND VPWR VPWR _21568_/B sky130_fd_sc_hd__or4_4
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12405_ _12405_/A VGND VGND VPWR VPWR _12405_/Y sky130_fd_sc_hd__inv_2
X_13385_ _13385_/A _13377_/X _13384_/X VGND VGND VPWR VPWR _13385_/X sky130_fd_sc_hd__and3_4
X_16173_ _16173_/A _16168_/X _16170_/X _16172_/X VGND VGND VPWR VPWR _16174_/A sky130_fd_sc_hd__or4_4
X_15124_ _15123_/Y _16415_/A _15123_/Y _16415_/A VGND VGND VPWR VPWR _15127_/C sky130_fd_sc_hd__a2bb2o_4
X_12336_ _12985_/B _24832_/Q _12985_/B _24832_/Q VGND VGND VPWR VPWR _12336_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23207__B1 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_16_0_HCLK clkbuf_5_8_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_33_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_12267_ _25443_/Q VGND VGND VPWR VPWR _12267_/Y sky130_fd_sc_hd__inv_2
X_15055_ _15192_/A _15189_/A VGND VGND VPWR VPWR _15055_/X sky130_fd_sc_hd__or2_4
X_19932_ _19932_/A VGND VGND VPWR VPWR _19932_/X sky130_fd_sc_hd__buf_2
XFILLER_141_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14006_ _14006_/A VGND VGND VPWR VPWR _14006_/Y sky130_fd_sc_hd__inv_2
X_19863_ _19861_/Y _19857_/X _19606_/X _19862_/X VGND VGND VPWR VPWR _23592_/D sky130_fd_sc_hd__a2bb2o_4
X_12198_ _22410_/A VGND VGND VPWR VPWR _12198_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22431__A _23172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18814_ _18813_/X VGND VGND VPWR VPWR _18814_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19794_ _19793_/Y _19789_/X _19728_/X _19789_/X VGND VGND VPWR VPWR _23614_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18745_ _18778_/A _18694_/B _18745_/C _18745_/D VGND VGND VPWR VPWR _18767_/B sky130_fd_sc_hd__or4_4
XANTENNA__21047__A _21579_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13772__B _16721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15957_ _15955_/X _15928_/X HWDATA[16] _24764_/Q _15956_/X VGND VGND VPWR VPWR _24764_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14908_ _14908_/A VGND VGND VPWR VPWR _14908_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19740__A _19740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18676_ _24151_/Q VGND VGND VPWR VPWR _18733_/A sky130_fd_sc_hd__inv_2
X_15888_ _15701_/X _15887_/X _16240_/A _24796_/Q _15857_/A VGND VGND VPWR VPWR _15888_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__24934__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17627_ _17627_/A VGND VGND VPWR VPWR _17647_/A sky130_fd_sc_hd__buf_2
X_14839_ _14820_/X _14837_/Y _25051_/Q _14838_/X VGND VGND VPWR VPWR _14839_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15620__B1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23143__C1 _23142_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17558_ _17627_/A VGND VGND VPWR VPWR _17620_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_5_26_0_HCLK_A clkbuf_5_27_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16509_ _16507_/Y _16508_/X _16240_/X _16508_/X VGND VGND VPWR VPWR _24558_/D sky130_fd_sc_hd__a2bb2o_4
X_17489_ _17488_/X VGND VGND VPWR VPWR _17489_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19228_ _23811_/Q VGND VGND VPWR VPWR _19228_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19159_ _19158_/Y _19156_/X _19067_/X _19156_/X VGND VGND VPWR VPWR _23836_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_191_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22170_ _23930_/Q VGND VGND VPWR VPWR _22170_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21121_ _21121_/A VGND VGND VPWR VPWR _22992_/A sky130_fd_sc_hd__buf_2
XANTENNA__11748__A _16240_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22957__C1 _22956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21052_ _24855_/Q _21031_/X _21034_/X _21051_/X VGND VGND VPWR VPWR _21053_/C sky130_fd_sc_hd__a211o_4
XANTENNA__22421__A1 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22421__B2 _22282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20003_ _19990_/Y VGND VGND VPWR VPWR _20003_/X sky130_fd_sc_hd__buf_2
XFILLER_101_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24811_ _24886_/CLK _15867_/X HRESETn VGND VGND VPWR VPWR _24811_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_36_0_HCLK clkbuf_8_37_0_HCLK/A VGND VGND VPWR VPWR _23528_/CLK sky130_fd_sc_hd__clkbuf_1
X_24742_ _24639_/CLK _16008_/X HRESETn VGND VGND VPWR VPWR _16006_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19050__B1 _19006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21954_ _21954_/A _21946_/X _21954_/C VGND VGND VPWR VPWR _21954_/X sky130_fd_sc_hd__or3_4
Xclkbuf_8_99_0_HCLK clkbuf_8_98_0_HCLK/A VGND VGND VPWR VPWR _24634_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24675__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23172__A _23172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20905_ _20892_/X _20904_/Y _24496_/Q _20896_/X VGND VGND VPWR VPWR _24052_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_242_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _21913_/A _19240_/Y VGND VGND VPWR VPWR _21885_/X sky130_fd_sc_hd__or2_4
X_24673_ _24678_/CLK _16199_/X HRESETn VGND VGND VPWR VPWR _23170_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24604__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15611__B1 _11753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _16711_/Y _20825_/X _20834_/X _20835_/X VGND VGND VPWR VPWR _20837_/A sky130_fd_sc_hd__o22a_4
X_23624_ _23610_/CLK _23624_/D VGND VGND VPWR VPWR _19768_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_230_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20499__B1 _20477_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20767_ _20767_/A VGND VGND VPWR VPWR _20767_/Y sky130_fd_sc_hd__inv_2
X_23555_ _23555_/CLK _19958_/X VGND VGND VPWR VPWR _19957_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17364__B1 _17268_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__A _13433_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22506_ _16596_/Y _22452_/X _21582_/X _22505_/X VGND VGND VPWR VPWR _22506_/X sky130_fd_sc_hd__o22a_4
XFILLER_183_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23486_ _23487_/CLK _20148_/X VGND VGND VPWR VPWR _23486_/Q sky130_fd_sc_hd__dfxtp_4
X_20698_ _21593_/A _20687_/X _20696_/X _20697_/X VGND VGND VPWR VPWR _20698_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22437_ _22437_/A _22437_/B VGND VGND VPWR VPWR _22443_/C sky130_fd_sc_hd__nor2_4
X_25225_ _23932_/CLK _14110_/X HRESETn VGND VGND VPWR VPWR _14094_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21420__A _22466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13170_ _13170_/A _19207_/A VGND VGND VPWR VPWR _13170_/X sky130_fd_sc_hd__or2_4
X_22368_ _22387_/A _20177_/Y VGND VGND VPWR VPWR _22369_/C sky130_fd_sc_hd__or2_4
X_25156_ _25158_/CLK _25156_/D HRESETn VGND VGND VPWR VPWR _25156_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12121_ _24101_/Q _24102_/Q _12120_/Y VGND VGND VPWR VPWR _20971_/A sky130_fd_sc_hd__o21a_4
XFILLER_184_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21319_ _21111_/A VGND VGND VPWR VPWR _21319_/X sky130_fd_sc_hd__buf_2
X_24107_ _24188_/CLK _24107_/D HRESETn VGND VGND VPWR VPWR _12139_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__11658__A _24067_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25087_ _25089_/CLK _25087_/D HRESETn VGND VGND VPWR VPWR _13569_/A sky130_fd_sc_hd__dfrtp_4
X_22299_ _21022_/A VGND VGND VPWR VPWR _22299_/X sky130_fd_sc_hd__buf_2
XFILLER_123_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12052_ _21568_/A VGND VGND VPWR VPWR _12058_/C sky130_fd_sc_hd__buf_2
X_24038_ _24594_/CLK _20841_/Y HRESETn VGND VGND VPWR VPWR _24038_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17419__B2 _17414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16860_ _16854_/X VGND VGND VPWR VPWR _16860_/X sky130_fd_sc_hd__buf_2
X_15811_ _15811_/A VGND VGND VPWR VPWR _15811_/X sky130_fd_sc_hd__buf_2
XFILLER_237_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16791_ _24445_/Q VGND VGND VPWR VPWR _16791_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18530_ _18523_/X _18530_/B _18530_/C VGND VGND VPWR VPWR _24179_/D sky130_fd_sc_hd__and3_4
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22715__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15742_ _15724_/X _15738_/X _15741_/X _24869_/Q _15736_/X VGND VGND VPWR VPWR _15742_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__19041__B1 _18948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12954_ _25373_/Q _12954_/B VGND VGND VPWR VPWR _12954_/X sky130_fd_sc_hd__or2_4
XFILLER_219_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11905_ _19606_/A VGND VGND VPWR VPWR _11905_/Y sky130_fd_sc_hd__inv_2
X_18461_ _18461_/A VGND VGND VPWR VPWR _18462_/A sky130_fd_sc_hd__inv_2
X_15673_ _15688_/A VGND VGND VPWR VPWR _15673_/X sky130_fd_sc_hd__buf_2
X_12885_ _12861_/A _12885_/B _12884_/X VGND VGND VPWR VPWR _25391_/D sky130_fd_sc_hd__and3_4
XFILLER_73_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24345__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_7_0_HCLK clkbuf_5_7_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_7_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15602__B1 _11739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17411_/X VGND VGND VPWR VPWR _17412_/X sky130_fd_sc_hd__buf_2
XFILLER_233_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14624_ _14623_/Y _14611_/Y _14606_/A _14610_/X VGND VGND VPWR VPWR _25079_/D sky130_fd_sc_hd__o22a_4
XFILLER_221_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11836_/A VGND VGND VPWR VPWR _13668_/B sky130_fd_sc_hd__inv_2
X_18392_ _21013_/B _17268_/X _18391_/Y VGND VGND VPWR VPWR _24190_/D sky130_fd_sc_hd__o21a_4
XFILLER_233_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17240_/D _17343_/B VGND VGND VPWR VPWR _17344_/B sky130_fd_sc_hd__or2_4
X_14555_ _14548_/Y _14554_/X VGND VGND VPWR VPWR _14555_/X sky130_fd_sc_hd__or2_4
XPHY_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11763_/Y _11756_/X _11765_/X _11766_/X VGND VGND VPWR VPWR _25526_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14209__A _14209_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _13506_/A VGND VGND VPWR VPWR _20964_/B sky130_fd_sc_hd__buf_2
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17274_ _17191_/Y _17272_/A VGND VGND VPWR VPWR _17274_/X sky130_fd_sc_hd__or2_4
XFILLER_159_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14486_ _14530_/A _14484_/X _14485_/X VGND VGND VPWR VPWR _14487_/A sky130_fd_sc_hd__o21a_4
XFILLER_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11698_ _11697_/Y VGND VGND VPWR VPWR _11699_/A sky130_fd_sc_hd__buf_2
XFILLER_158_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19013_ _18083_/B VGND VGND VPWR VPWR _19013_/Y sky130_fd_sc_hd__inv_2
X_16225_ _22741_/A VGND VGND VPWR VPWR _16225_/Y sky130_fd_sc_hd__inv_2
X_13437_ _13300_/A _13435_/X _13436_/X VGND VGND VPWR VPWR _13437_/X sky130_fd_sc_hd__and3_4
XFILLER_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18644__A1_N _24516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22100__B1 _22098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22145__B _22145_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23980__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16156_ _16154_/Y _16150_/X _15466_/X _16155_/X VGND VGND VPWR VPWR _24685_/D sky130_fd_sc_hd__a2bb2o_4
X_13368_ _13193_/A _13368_/B _13367_/X VGND VGND VPWR VPWR _13369_/C sky130_fd_sc_hd__and3_4
XANTENNA__13767__B _14208_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15107_ _15107_/A VGND VGND VPWR VPWR _15107_/Y sky130_fd_sc_hd__inv_2
X_12319_ _24829_/Q VGND VGND VPWR VPWR _12319_/Y sky130_fd_sc_hd__inv_2
X_16087_ _16081_/Y _16086_/X _15991_/X _16086_/X VGND VGND VPWR VPWR _24712_/D sky130_fd_sc_hd__a2bb2o_4
X_13299_ _13431_/A _13299_/B VGND VGND VPWR VPWR _13299_/X sky130_fd_sc_hd__or2_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15038_ _14913_/A _15037_/Y _14913_/A _15037_/Y VGND VGND VPWR VPWR _15038_/X sky130_fd_sc_hd__a2bb2o_4
X_19915_ _21402_/B _19912_/X _19827_/X _19912_/X VGND VGND VPWR VPWR _19915_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15684__A3 _15694_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25141__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14879__A pwm_S6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13783__A _16721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17255__A _17255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19846_ _23597_/Q VGND VGND VPWR VPWR _19846_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19280__B1 _19279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16989_ _24733_/Q _17103_/A _16061_/Y _16991_/A VGND VGND VPWR VPWR _16995_/A sky130_fd_sc_hd__a2bb2o_4
X_19777_ _21610_/B _19776_/X _16882_/X _19776_/X VGND VGND VPWR VPWR _23621_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_252_0_HCLK clkbuf_7_126_0_HCLK/X VGND VGND VPWR VPWR _24074_/CLK sky130_fd_sc_hd__clkbuf_1
X_18728_ _18728_/A _18695_/X _18745_/C VGND VGND VPWR VPWR _18729_/B sky130_fd_sc_hd__or3_4
XFILLER_243_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18659_ _16554_/Y _24152_/Q _16569_/A _18658_/Y VGND VGND VPWR VPWR _18662_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24086__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21670_ _21924_/A VGND VGND VPWR VPWR _21670_/X sky130_fd_sc_hd__buf_2
XFILLER_169_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24015__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20621_ _17385_/X _20619_/Y _20621_/C VGND VGND VPWR VPWR _20621_/X sky130_fd_sc_hd__and3_4
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21142__A1 _21343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23340_ _13790_/Y _25070_/Q _13794_/Y _25057_/Q VGND VGND VPWR VPWR _23341_/A sky130_fd_sc_hd__o22a_4
XFILLER_149_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16937__A2_N _24262_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20552_ _23939_/Q _18872_/X VGND VGND VPWR VPWR _20552_/Y sky130_fd_sc_hd__nand2_4
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23271_ _21446_/X _23269_/X _22691_/X _23270_/X VGND VGND VPWR VPWR _23272_/A sky130_fd_sc_hd__o22a_4
XANTENNA__19099__B1 _18981_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20483_ _20482_/X VGND VGND VPWR VPWR _20483_/X sky130_fd_sc_hd__buf_2
X_22222_ _22210_/A _22222_/B VGND VGND VPWR VPWR _22222_/X sky130_fd_sc_hd__or2_4
X_25010_ _24477_/CLK _25010_/D HRESETn VGND VGND VPWR VPWR _25010_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22153_ _22153_/A _22145_/B VGND VGND VPWR VPWR _22153_/X sky130_fd_sc_hd__or2_4
X_21104_ _24645_/Q _15651_/A _21103_/X _21042_/X VGND VGND VPWR VPWR _21105_/A sky130_fd_sc_hd__a211o_4
X_22084_ _22386_/A _22084_/B VGND VGND VPWR VPWR _22084_/X sky130_fd_sc_hd__or2_4
XANTENNA__22071__A _22199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_62_0_HCLK clkbuf_6_63_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_62_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_21035_ _11678_/X VGND VGND VPWR VPWR _22132_/B sky130_fd_sc_hd__buf_2
XFILLER_120_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24856__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15832__B1 _24823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19023__B1 _18998_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22986_ _17249_/C _22916_/X _12895_/A _22917_/X VGND VGND VPWR VPWR _22986_/X sky130_fd_sc_hd__a2bb2o_4
X_24725_ _24725_/CLK _24725_/D HRESETn VGND VGND VPWR VPWR _24725_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21937_ _21937_/A _21937_/B _21937_/C VGND VGND VPWR VPWR _21937_/X sky130_fd_sc_hd__and3_4
XFILLER_28_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12670_ _12677_/A _12670_/B _12670_/C VGND VGND VPWR VPWR _25419_/D sky130_fd_sc_hd__and3_4
X_24656_ _24654_/CLK _24656_/D HRESETn VGND VGND VPWR VPWR _16244_/A sky130_fd_sc_hd__dfrtp_4
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21868_ _21537_/X VGND VGND VPWR VPWR _21868_/X sky130_fd_sc_hd__buf_2
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ _23487_/CLK _23607_/D VGND VGND VPWR VPWR _19816_/A sky130_fd_sc_hd__dfxtp_4
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20819_ _20817_/Y _20818_/Y _13125_/X VGND VGND VPWR VPWR _20819_/X sky130_fd_sc_hd__o21a_4
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21799_ _21662_/A _21799_/B VGND VGND VPWR VPWR _21799_/X sky130_fd_sc_hd__or2_4
X_24587_ _24591_/CLK _16425_/X HRESETn VGND VGND VPWR VPWR _24587_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22330__B1 _20673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ _14338_/B VGND VGND VPWR VPWR _14340_/X sky130_fd_sc_hd__buf_2
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23538_ _23415_/CLK _23538_/D VGND VGND VPWR VPWR _23538_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22881__B2 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14271_ _23966_/Q VGND VGND VPWR VPWR _14271_/X sky130_fd_sc_hd__buf_2
X_23469_ _23378_/CLK _20193_/X VGND VGND VPWR VPWR _20191_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12772__A _12772_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16010_ _16009_/Y _16007_/X _11685_/X _16007_/X VGND VGND VPWR VPWR _16010_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13222_ _13199_/A VGND VGND VPWR VPWR _13443_/A sky130_fd_sc_hd__buf_2
X_25208_ _24146_/CLK _14193_/X HRESETn VGND VGND VPWR VPWR _20516_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_183_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13153_ _13168_/A VGND VGND VPWR VPWR _13175_/A sky130_fd_sc_hd__buf_2
X_25139_ _25140_/CLK _25139_/D HRESETn VGND VGND VPWR VPWR _14417_/A sky130_fd_sc_hd__dfstp_4
XFILLER_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12104_ _25472_/Q VGND VGND VPWR VPWR _12104_/Y sky130_fd_sc_hd__inv_2
X_13084_ _13072_/A _13072_/B VGND VGND VPWR VPWR _13084_/Y sky130_fd_sc_hd__nand2_4
X_17961_ _17957_/X _17960_/X _18009_/A VGND VGND VPWR VPWR _17961_/X sky130_fd_sc_hd__o21a_4
XFILLER_97_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14699__A _13731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12035_ _15636_/A VGND VGND VPWR VPWR _13454_/A sky130_fd_sc_hd__inv_2
X_16912_ _22909_/A _24277_/Q _16115_/Y _16911_/Y VGND VGND VPWR VPWR _16919_/A sky130_fd_sc_hd__o22a_4
X_19700_ _19698_/Y _19694_/X _19633_/X _19699_/X VGND VGND VPWR VPWR _23648_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17892_ _17892_/A VGND VGND VPWR VPWR _17906_/B sky130_fd_sc_hd__buf_2
XFILLER_238_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24597__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16843_ _14940_/Y _16841_/X _16525_/X _16841_/X VGND VGND VPWR VPWR _24419_/D sky130_fd_sc_hd__a2bb2o_4
X_19631_ _19629_/Y _19627_/X _19630_/X _19627_/X VGND VGND VPWR VPWR _19631_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24526__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19562_ _19549_/Y VGND VGND VPWR VPWR _19562_/X sky130_fd_sc_hd__buf_2
XANTENNA__19014__B1 _18942_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16774_ _16766_/A VGND VGND VPWR VPWR _16774_/X sky130_fd_sc_hd__buf_2
X_13986_ _25237_/Q VGND VGND VPWR VPWR _13986_/X sky130_fd_sc_hd__buf_2
X_18513_ _18462_/A _18516_/B _18489_/X VGND VGND VPWR VPWR _18513_/Y sky130_fd_sc_hd__a21oi_4
X_15725_ HWDATA[23] VGND VGND VPWR VPWR _15725_/X sky130_fd_sc_hd__buf_2
X_12937_ _12834_/A _12756_/X _12931_/X VGND VGND VPWR VPWR _12937_/X sky130_fd_sc_hd__or3_4
X_19493_ _23717_/Q VGND VGND VPWR VPWR _19493_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12947__A _12781_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_82_0_HCLK clkbuf_8_83_0_HCLK/A VGND VGND VPWR VPWR _24765_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_160_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11851__A _11934_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18444_ _24180_/Q VGND VGND VPWR VPWR _18510_/C sky130_fd_sc_hd__inv_2
XFILLER_222_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15656_ _15639_/Y _15651_/X _15643_/X _20822_/A _15655_/X VGND VGND VPWR VPWR _15656_/X
+ sky130_fd_sc_hd__a32o_4
X_12868_ _12735_/Y _12868_/B VGND VGND VPWR VPWR _12869_/C sky130_fd_sc_hd__or2_4
XFILLER_233_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14604_/Y _14610_/A _14606_/Y VGND VGND VPWR VPWR _14607_/Y sky130_fd_sc_hd__o21ai_4
X_11819_ _25296_/Q _22735_/A _11804_/A _22584_/A VGND VGND VPWR VPWR _11822_/C sky130_fd_sc_hd__a2bb2o_4
X_18375_ _18371_/Y _18374_/X _18376_/A _18374_/X VGND VGND VPWR VPWR _24198_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15587_ _22922_/A _15584_/X _11715_/X _15584_/X VGND VGND VPWR VPWR _24912_/D sky130_fd_sc_hd__a2bb2o_4
X_12799_ _12838_/B _24802_/Q _12895_/A _12746_/Y VGND VGND VPWR VPWR _12799_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22321__B1 _12197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17326_ _17248_/Y _17304_/X VGND VGND VPWR VPWR _17329_/B sky130_fd_sc_hd__or2_4
X_14538_ _14531_/X _14537_/Y sda_oen_o_S4 _14531_/X VGND VGND VPWR VPWR _25100_/D
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25385__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_HCLK clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_5_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_186_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21060__A _22807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17257_ _17333_/A _17265_/A VGND VGND VPWR VPWR _17271_/B sky130_fd_sc_hd__or2_4
X_14469_ _14467_/Y _14463_/X _14407_/X _14468_/X VGND VGND VPWR VPWR _14469_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16208_ _16207_/Y _16203_/X _15942_/X _16203_/X VGND VGND VPWR VPWR _16208_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18828__B1 _24552_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17188_ _17180_/X _17188_/B _17184_/X _17188_/D VGND VGND VPWR VPWR _17188_/X sky130_fd_sc_hd__or4_4
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16139_ _16138_/Y _16136_/X _15965_/X _16136_/X VGND VGND VPWR VPWR _24691_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14402__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19829_ _19829_/A VGND VGND VPWR VPWR _21238_/B sky130_fd_sc_hd__inv_2
XFILLER_110_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24267__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15814__B1 _24835_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22840_ _22840_/A VGND VGND VPWR VPWR _23263_/B sky130_fd_sc_hd__buf_2
XANTENNA__12628__B1 _12627_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22771_ _24801_/Q _22901_/B VGND VGND VPWR VPWR _22771_/X sky130_fd_sc_hd__or2_4
XFILLER_240_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22560__B1 _24830_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24510_ _24910_/CLK _16638_/X HRESETn VGND VGND VPWR VPWR _23323_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15233__A _15059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11761__A _11760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21722_ _21722_/A _21722_/B VGND VGND VPWR VPWR _21722_/Y sky130_fd_sc_hd__nor2_4
X_25490_ _25466_/CLK _12028_/X HRESETn VGND VGND VPWR VPWR _25490_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21653_ _21641_/Y _21652_/Y _13772_/C VGND VGND VPWR VPWR _21697_/C sky130_fd_sc_hd__o21a_4
X_24441_ _24443_/CLK _24441_/D HRESETn VGND VGND VPWR VPWR _24441_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_220_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21115__A1 _17239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_200_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20604_ _20603_/A VGND VGND VPWR VPWR _20604_/Y sky130_fd_sc_hd__inv_2
X_21584_ _16532_/Y _21741_/B VGND VGND VPWR VPWR _21584_/X sky130_fd_sc_hd__and2_4
X_24372_ _24641_/CLK _24372_/D HRESETn VGND VGND VPWR VPWR _17261_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_177_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20535_ _24073_/Q _20535_/B VGND VGND VPWR VPWR _20535_/X sky130_fd_sc_hd__and2_4
X_23323_ _23323_/A _16792_/A VGND VGND VPWR VPWR _23323_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__25055__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16064__A _24720_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20466_ _20437_/A _20466_/B VGND VGND VPWR VPWR _20466_/X sky130_fd_sc_hd__and2_4
X_23254_ _24745_/Q _21031_/X _21034_/X _23253_/X VGND VGND VPWR VPWR _23254_/X sky130_fd_sc_hd__a211o_4
XFILLER_153_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__20626__B1 _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22205_ _22205_/A _22205_/B _22204_/X VGND VGND VPWR VPWR _22213_/B sky130_fd_sc_hd__or3_4
XFILLER_180_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23185_ _23035_/X _23184_/X _23145_/X _24847_/Q _23037_/X VGND VGND VPWR VPWR _23185_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_180_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20397_ _20396_/Y _20394_/X _15762_/X _20394_/X VGND VGND VPWR VPWR _23389_/D sky130_fd_sc_hd__a2bb2o_4
X_22136_ _24898_/Q _22136_/B VGND VGND VPWR VPWR _22136_/X sky130_fd_sc_hd__or2_4
XFILLER_106_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22067_ _22365_/A _22067_/B VGND VGND VPWR VPWR _22068_/C sky130_fd_sc_hd__or2_4
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24690__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21018_ _25299_/Q _21018_/B VGND VGND VPWR VPWR _23371_/A sky130_fd_sc_hd__and2_4
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15805__B1 _11711_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18719__A _18774_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13840_ _20476_/A _20476_/B _13840_/C VGND VGND VPWR VPWR _13842_/B sky130_fd_sc_hd__or3_4
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23343__A2 _21970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13771_ _13771_/A VGND VGND VPWR VPWR _13772_/D sky130_fd_sc_hd__buf_2
X_22969_ _22474_/X _22968_/X _22858_/X _12296_/A _22478_/X VGND VGND VPWR VPWR _22969_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_43_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21354__B2 _14245_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15510_ _24937_/Q VGND VGND VPWR VPWR _15510_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_69_0_HCLK clkbuf_7_69_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_69_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_12722_ _12722_/A _12721_/Y _12722_/C VGND VGND VPWR VPWR _25403_/D sky130_fd_sc_hd__and3_4
X_24708_ _24704_/CLK _24708_/D HRESETn VGND VGND VPWR VPWR _23193_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_231_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16490_ _24565_/Q VGND VGND VPWR VPWR _16490_/Y sky130_fd_sc_hd__inv_2
X_15441_ _15426_/X VGND VGND VPWR VPWR _15441_/X sky130_fd_sc_hd__buf_2
XANTENNA__23360__A _23344_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12653_ _12592_/Y _12606_/X VGND VGND VPWR VPWR _12662_/B sky130_fd_sc_hd__or2_4
X_24639_ _24639_/CLK _24639_/D HRESETn VGND VGND VPWR VPWR _23190_/A sky130_fd_sc_hd__dfrtp_4
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22303__B1 _22140_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21106__B2 _21736_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18454__A _18745_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18160_ _18128_/A _23829_/Q VGND VGND VPWR VPWR _18160_/X sky130_fd_sc_hd__or2_4
XFILLER_157_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ _15371_/X VGND VGND VPWR VPWR _24990_/D sky130_fd_sc_hd__inv_2
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12578_/Y VGND VGND VPWR VPWR _12584_/X sky130_fd_sc_hd__buf_2
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17111_ _24388_/Q _17111_/B VGND VGND VPWR VPWR _17111_/X sky130_fd_sc_hd__or2_4
XFILLER_156_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _18372_/B _14324_/B _14314_/X VGND VGND VPWR VPWR _25167_/D sky130_fd_sc_hd__a21o_4
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18091_ _18057_/A VGND VGND VPWR VPWR _18125_/A sky130_fd_sc_hd__buf_2
XFILLER_156_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17042_ _17042_/A _17038_/X _17042_/C VGND VGND VPWR VPWR _17042_/X sky130_fd_sc_hd__or3_4
X_14254_ _25189_/Q VGND VGND VPWR VPWR _14254_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13205_ _13289_/A VGND VGND VPWR VPWR _13363_/A sky130_fd_sc_hd__buf_2
XANTENNA__20617__B1 _20672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14185_ _13873_/X _23998_/Q VGND VGND VPWR VPWR _14185_/X sky130_fd_sc_hd__or2_4
XFILLER_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24778__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13136_ _13167_/A VGND VGND VPWR VPWR _13170_/A sky130_fd_sc_hd__buf_2
XFILLER_124_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18993_ _18986_/A VGND VGND VPWR VPWR _18993_/X sky130_fd_sc_hd__buf_2
XFILLER_3_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24707__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13067_ _12983_/D _12971_/Y VGND VGND VPWR VPWR _13068_/D sky130_fd_sc_hd__or2_4
X_17944_ _17944_/A _23826_/Q VGND VGND VPWR VPWR _17945_/C sky130_fd_sc_hd__or2_4
XFILLER_78_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12018_ _12017_/Y _12015_/X _12019_/A _12015_/X VGND VGND VPWR VPWR _25494_/D sky130_fd_sc_hd__a2bb2o_4
X_17875_ _17853_/D VGND VGND VPWR VPWR _17876_/B sky130_fd_sc_hd__inv_2
XFILLER_120_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24360__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19614_ _21817_/B _19607_/X _19613_/X _19607_/X VGND VGND VPWR VPWR _23678_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_241_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16826_ _24428_/Q VGND VGND VPWR VPWR _16826_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23334__A2 _22661_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16757_ _24461_/Q VGND VGND VPWR VPWR _16757_/Y sky130_fd_sc_hd__inv_2
X_19545_ _23699_/Q VGND VGND VPWR VPWR _19545_/Y sky130_fd_sc_hd__inv_2
X_13969_ _14007_/B VGND VGND VPWR VPWR _13969_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22542__B1 _21956_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16149__A _22191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15708_ _15540_/X _15701_/X _15702_/X _24886_/Q _15707_/X VGND VGND VPWR VPWR _15708_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__14679__A2_N _14678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16688_ _16687_/Y _16685_/X _15746_/X _16685_/X VGND VGND VPWR VPWR _16688_/X sky130_fd_sc_hd__a2bb2o_4
X_19476_ _21188_/B _19470_/X _19475_/X _19457_/Y VGND VGND VPWR VPWR _23723_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15639_ _15671_/A VGND VGND VPWR VPWR _15639_/Y sky130_fd_sc_hd__inv_2
X_18427_ _22814_/A _18467_/B _16254_/Y _24163_/Q VGND VGND VPWR VPWR _18433_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18358_ _18365_/A _18365_/B _18357_/Y VGND VGND VPWR VPWR _18358_/X sky130_fd_sc_hd__a21o_4
XANTENNA__14783__B1 _18020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17309_ _17174_/A _17309_/B VGND VGND VPWR VPWR _17311_/B sky130_fd_sc_hd__or2_4
X_18289_ _18288_/X VGND VGND VPWR VPWR _18289_/X sky130_fd_sc_hd__buf_2
X_20320_ _23420_/Q VGND VGND VPWR VPWR _20320_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22614__A _22581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20251_ _20250_/Y _20248_/X _16867_/X _20248_/X VGND VGND VPWR VPWR _23447_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23270__B2 _22821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16288__B1 _16001_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20084__B2 _20067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20182_ _23473_/Q VGND VGND VPWR VPWR _22225_/B sky130_fd_sc_hd__inv_2
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24448__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17544__A2_N _25546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24990_ _25005_/CLK _24990_/D HRESETn VGND VGND VPWR VPWR _24990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12313__A2 _24827_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23941_ _23938_/CLK _23941_/D HRESETn VGND VGND VPWR VPWR _18875_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_130_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18539__A _18467_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23872_ _23853_/CLK _23872_/D VGND VGND VPWR VPWR _23872_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_244_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24030__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22823_ _22946_/A _22820_/X _22822_/X VGND VGND VPWR VPWR _22856_/B sky130_fd_sc_hd__and3_4
XANTENNA__16059__A _14403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25542_ _24310_/CLK _25542_/D HRESETn VGND VGND VPWR VPWR _25542_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22754_ _22149_/X _22753_/X _22146_/X _25535_/Q _22554_/X VGND VGND VPWR VPWR _22754_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_197_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21705_ _21581_/X _21704_/X _21436_/X _24823_/Q _21336_/X VGND VGND VPWR VPWR _21706_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_212_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25473_ _24325_/CLK _12103_/X HRESETn VGND VGND VPWR VPWR _25473_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22685_ _21122_/X _22683_/X _21227_/X _22684_/X VGND VGND VPWR VPWR _22686_/B sky130_fd_sc_hd__o22a_4
XFILLER_198_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_201_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24424_ _24463_/CLK _24424_/D HRESETn VGND VGND VPWR VPWR _24424_/Q sky130_fd_sc_hd__dfrtp_4
X_21636_ _21609_/X _21636_/B VGND VGND VPWR VPWR _21636_/X sky130_fd_sc_hd__or2_4
XFILLER_166_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24355_ _24341_/CLK _17332_/Y HRESETn VGND VGND VPWR VPWR _22709_/A sky130_fd_sc_hd__dfrtp_4
X_21567_ _21730_/A _21567_/B VGND VGND VPWR VPWR _21567_/X sky130_fd_sc_hd__and2_4
XANTENNA__13211__A _13289_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23306_ _23287_/X _23290_/X _23294_/Y _23305_/X VGND VGND VPWR VPWR HRDATA[30] sky130_fd_sc_hd__a211o_4
XFILLER_176_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20518_ _20516_/X _20517_/X _15451_/X VGND VGND VPWR VPWR _20518_/X sky130_fd_sc_hd__o21a_4
X_21498_ _21493_/X _21497_/X _18301_/X VGND VGND VPWR VPWR _21498_/X sky130_fd_sc_hd__o21a_4
X_24286_ _24275_/CLK _24286_/D HRESETn VGND VGND VPWR VPWR _24286_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20449_ _23928_/Q VGND VGND VPWR VPWR _20449_/X sky130_fd_sc_hd__buf_2
X_23237_ _23169_/A _23236_/X VGND VGND VPWR VPWR _23237_/Y sky130_fd_sc_hd__nor2_4
XFILLER_134_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16522__A _14403_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24871__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21272__B1 _14672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23168_ _20800_/Y _22992_/X _20939_/Y _22794_/X VGND VGND VPWR VPWR _23169_/B sky130_fd_sc_hd__o22a_4
XANTENNA__24189__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24800__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22119_ _25249_/Q _22119_/B VGND VGND VPWR VPWR _22119_/X sky130_fd_sc_hd__and2_4
XANTENNA__19217__B1 _19125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15990_ _15990_/A VGND VGND VPWR VPWR _15990_/X sky130_fd_sc_hd__buf_2
X_23099_ _23094_/Y _23098_/Y _22854_/X VGND VGND VPWR VPWR _23099_/X sky130_fd_sc_hd__o21a_4
XANTENNA__24118__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14941_ _25009_/Q _14939_/Y _25013_/Q _14940_/Y VGND VGND VPWR VPWR _14946_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_248_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17660_ _17660_/A _17660_/B VGND VGND VPWR VPWR _17661_/C sky130_fd_sc_hd__or2_4
XFILLER_235_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14872_ _14859_/B _14866_/X _14867_/Y VGND VGND VPWR VPWR _14872_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_48_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16611_ _16547_/A VGND VGND VPWR VPWR _16611_/X sky130_fd_sc_hd__buf_2
X_13823_ _13562_/Y _13817_/X _11757_/X _13822_/X VGND VGND VPWR VPWR _13823_/X sky130_fd_sc_hd__a2bb2o_4
X_17591_ _17620_/A _17589_/X _17590_/X VGND VGND VPWR VPWR _24322_/D sky130_fd_sc_hd__and3_4
XFILLER_235_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21306__C _21306_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22524__B1 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16542_ _16541_/X VGND VGND VPWR VPWR _16542_/X sky130_fd_sc_hd__buf_2
X_19330_ _19329_/Y _19327_/X _19194_/X _19327_/X VGND VGND VPWR VPWR _23775_/D sky130_fd_sc_hd__a2bb2o_4
X_13754_ _13737_/X VGND VGND VPWR VPWR _13754_/X sky130_fd_sc_hd__buf_2
XFILLER_189_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15006__B2 _15005_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12705_ _12686_/A _12696_/B _12705_/C VGND VGND VPWR VPWR _25409_/D sky130_fd_sc_hd__and3_4
X_19261_ _19261_/A VGND VGND VPWR VPWR _19261_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21603__A _22056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16473_ _16472_/Y _16470_/X _16295_/X _16470_/X VGND VGND VPWR VPWR _16473_/X sky130_fd_sc_hd__a2bb2o_4
X_13685_ _11806_/Y _13679_/A VGND VGND VPWR VPWR _13686_/B sky130_fd_sc_hd__or2_4
XFILLER_71_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18212_ _18052_/A _18208_/X _18211_/X VGND VGND VPWR VPWR _18212_/X sky130_fd_sc_hd__or3_4
X_15424_ _13939_/X _15424_/B _15424_/C _14234_/B VGND VGND VPWR VPWR _15430_/A sky130_fd_sc_hd__or4_4
X_12636_ _12627_/X _12632_/B _12636_/C VGND VGND VPWR VPWR _12636_/X sky130_fd_sc_hd__or3_4
X_19192_ _19190_/Y _19186_/X _19125_/X _19191_/X VGND VGND VPWR VPWR _19192_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22827__A1 _12838_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_156_0_HCLK clkbuf_7_78_0_HCLK/X VGND VGND VPWR VPWR _25471_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ _17972_/A _18143_/B VGND VGND VPWR VPWR _18143_/X sky130_fd_sc_hd__or2_4
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _15125_/Y _15347_/B VGND VGND VPWR VPWR _15355_/X sky130_fd_sc_hd__or2_4
X_12567_ _12567_/A VGND VGND VPWR VPWR _12638_/C sky130_fd_sc_hd__inv_2
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14217__A _20664_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24959__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ _25174_/Q _14288_/Y _25173_/Q _14296_/A VGND VGND VPWR VPWR _14306_/X sky130_fd_sc_hd__o22a_4
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18074_ _17987_/X _23743_/Q VGND VGND VPWR VPWR _18075_/C sky130_fd_sc_hd__or2_4
X_15286_ _15285_/Y VGND VGND VPWR VPWR _15331_/A sky130_fd_sc_hd__buf_2
XANTENNA__17007__A1_N _24738_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12498_ _25412_/Q VGND VGND VPWR VPWR _12498_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17025_ _24398_/Q VGND VGND VPWR VPWR _17026_/A sky130_fd_sc_hd__inv_2
X_14237_ _23967_/Q _13953_/A VGND VGND VPWR VPWR _15423_/A sky130_fd_sc_hd__or2_4
XFILLER_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23249__B _23075_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22153__B _22145_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24071__D _20471_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14168_ _14166_/Y _14099_/X _14125_/X _14167_/Y VGND VGND VPWR VPWR _14169_/A sky130_fd_sc_hd__o22a_4
XANTENNA__11751__B1 _25530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24541__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13119_ _20738_/A _13119_/B VGND VGND VPWR VPWR _13120_/B sky130_fd_sc_hd__or2_4
XFILLER_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19743__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14099_ _14099_/A VGND VGND VPWR VPWR _14099_/X sky130_fd_sc_hd__buf_2
X_18976_ _18975_/X VGND VGND VPWR VPWR _18986_/A sky130_fd_sc_hd__inv_2
XANTENNA__16690__B1 _15748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17927_ _17926_/X VGND VGND VPWR VPWR _17927_/Y sky130_fd_sc_hd__inv_2
XFILLER_239_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17858_ _17866_/A _17858_/B _17858_/C VGND VGND VPWR VPWR _24269_/D sky130_fd_sc_hd__and3_4
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16809_ _14914_/Y _16804_/X HWDATA[24] _16808_/X VGND VGND VPWR VPWR _16809_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_82_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17789_ _16898_/Y _17787_/A VGND VGND VPWR VPWR _17790_/C sky130_fd_sc_hd__or2_4
XANTENNA__21318__B2 _21317_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12838__C _12766_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19528_ _19528_/A VGND VGND VPWR VPWR _19528_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_52_0_HCLK clkbuf_7_53_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_52_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19459_ _22350_/B _19458_/X _11902_/X _19458_/X VGND VGND VPWR VPWR _23730_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_167_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22818__A1 _16576_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22470_ _20723_/A _21596_/X _15612_/Y _22452_/X VGND VGND VPWR VPWR _22470_/X sky130_fd_sc_hd__o22a_4
XFILLER_194_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21421_ _21421_/A VGND VGND VPWR VPWR _23328_/A sky130_fd_sc_hd__buf_2
XANTENNA__12231__B2 _24761_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21352_ _14417_/Y _21351_/X _14457_/Y _17411_/X VGND VGND VPWR VPWR _21353_/A sky130_fd_sc_hd__o22a_4
X_24140_ _24340_/CLK _24140_/D HRESETn VGND VGND VPWR VPWR _24140_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20303_ _21482_/B _20300_/X _19984_/X _20300_/X VGND VGND VPWR VPWR _20303_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24629__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21283_ _21283_/A VGND VGND VPWR VPWR _22515_/A sky130_fd_sc_hd__buf_2
X_24071_ _23427_/CLK _20471_/X HRESETn VGND VGND VPWR VPWR _13807_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__17438__A _14212_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23243__A1 _24474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20234_ _20227_/A VGND VGND VPWR VPWR _20234_/X sky130_fd_sc_hd__buf_2
X_23022_ _24602_/Q _23022_/B VGND VGND VPWR VPWR _23025_/B sky130_fd_sc_hd__or2_4
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24282__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20165_ _22085_/B _20159_/X _20095_/X _20164_/X VGND VGND VPWR VPWR _23480_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16681__B1 _15739_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20096_ _20088_/A VGND VGND VPWR VPWR _20096_/X sky130_fd_sc_hd__buf_2
X_24973_ _24973_/CLK _15435_/X HRESETn VGND VGND VPWR VPWR _24973_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_218_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13495__B1 _11775_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22754__B1 _25535_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23924_ _23926_/CLK _20977_/X HRESETn VGND VGND VPWR VPWR _23924_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25488__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16433__B1 _16353_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23855_ _23735_/CLK _23855_/D VGND VGND VPWR VPWR _23855_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22506__B1 _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22806_ _22806_/A _22890_/B VGND VGND VPWR VPWR _22806_/X sky130_fd_sc_hd__or2_4
XFILLER_26_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23786_ _25073_/CLK _19302_/X VGND VGND VPWR VPWR _17951_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_60_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20998_ scl_oen_o_S5 _20998_/B VGND VGND VPWR VPWR _20998_/X sky130_fd_sc_hd__and2_4
XFILLER_198_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25525_ _25524_/CLK _11771_/X HRESETn VGND VGND VPWR VPWR _25525_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22737_ _13650_/C _21303_/X _13121_/C _21317_/X VGND VGND VPWR VPWR _22737_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_201_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13470_ _13468_/Y _13464_/X _11770_/X _13469_/X VGND VGND VPWR VPWR _25322_/D sky130_fd_sc_hd__a2bb2o_4
X_25456_ _25382_/CLK _25456_/D HRESETn VGND VGND VPWR VPWR _25456_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22668_ _12418_/A _21532_/X _17755_/Y _22437_/A VGND VGND VPWR VPWR _22668_/X sky130_fd_sc_hd__o22a_4
XFILLER_185_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20039__A _20034_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_229_0_HCLK clkbuf_8_229_0_HCLK/A VGND VGND VPWR VPWR _24520_/CLK sky130_fd_sc_hd__clkbuf_1
X_12421_ _12248_/Y _12420_/X VGND VGND VPWR VPWR _12422_/A sky130_fd_sc_hd__or2_4
X_24407_ _23378_/CLK _24407_/D HRESETn VGND VGND VPWR VPWR _16880_/A sky130_fd_sc_hd__dfrtp_4
X_21619_ _21764_/A _21617_/X _21618_/X VGND VGND VPWR VPWR _21619_/X sky130_fd_sc_hd__and3_4
X_25387_ _25387_/CLK _12902_/X HRESETn VGND VGND VPWR VPWR _12766_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__19686__B1 _19540_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22599_ _24623_/Q _21337_/X VGND VGND VPWR VPWR _22599_/X sky130_fd_sc_hd__or2_4
XFILLER_139_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15140_ _23242_/A VGND VGND VPWR VPWR _15140_/Y sky130_fd_sc_hd__inv_2
X_12352_ _24848_/Q VGND VGND VPWR VPWR _12352_/Y sky130_fd_sc_hd__inv_2
X_24338_ _24340_/CLK _24338_/D HRESETn VGND VGND VPWR VPWR _21002_/B sky130_fd_sc_hd__dfstp_4
XFILLER_5_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15071_ _15070_/Y _16363_/A _15070_/Y _16363_/A VGND VGND VPWR VPWR _15077_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19438__B1 _19392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12283_ _12993_/A _24851_/Q _12993_/A _24851_/Q VGND VGND VPWR VPWR _12283_/X sky130_fd_sc_hd__a2bb2o_4
X_24269_ _24725_/CLK _24269_/D HRESETn VGND VGND VPWR VPWR _17747_/A sky130_fd_sc_hd__dfrtp_4
X_14022_ _25242_/Q _14022_/B VGND VGND VPWR VPWR _14034_/A sky130_fd_sc_hd__or2_4
XFILLER_106_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18830_ _18826_/X _18830_/B _18828_/X _18830_/D VGND VGND VPWR VPWR _18830_/X sky130_fd_sc_hd__or4_4
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18661__B2 _24146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15973_ _12220_/Y _15972_/X _15623_/X _15972_/X VGND VGND VPWR VPWR _15973_/X sky130_fd_sc_hd__a2bb2o_4
X_18761_ _18752_/A _18755_/X _18761_/C VGND VGND VPWR VPWR _18761_/X sky130_fd_sc_hd__and3_4
XANTENNA__13486__B1 _11753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21548__A1 _21289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14924_ _25037_/Q VGND VGND VPWR VPWR _15168_/A sky130_fd_sc_hd__inv_2
X_17712_ _19455_/B VGND VGND VPWR VPWR _18288_/A sky130_fd_sc_hd__inv_2
XFILLER_208_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18692_ _24142_/Q VGND VGND VPWR VPWR _18692_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16424__B1 _16145_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14855_ _14840_/X _14854_/Y _24956_/Q _14806_/X VGND VGND VPWR VPWR _14855_/X sky130_fd_sc_hd__a2bb2o_4
X_17643_ _17646_/A _17643_/B VGND VGND VPWR VPWR _17647_/B sky130_fd_sc_hd__or2_4
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13806_ _21642_/A VGND VGND VPWR VPWR _13807_/D sky130_fd_sc_hd__buf_2
XANTENNA__17811__A _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17574_ _17519_/Y _17670_/A _17513_/Y _17574_/D VGND VGND VPWR VPWR _17581_/A sky130_fd_sc_hd__or4_4
X_14786_ _19320_/A _14785_/X _19320_/A _14785_/X VGND VGND VPWR VPWR _14787_/D sky130_fd_sc_hd__a2bb2o_4
X_11998_ _11998_/A _11998_/B _11993_/X _11997_/X VGND VGND VPWR VPWR _11998_/X sky130_fd_sc_hd__or4_4
X_16525_ _14407_/A VGND VGND VPWR VPWR _16525_/X sky130_fd_sc_hd__buf_2
X_19313_ _19299_/Y VGND VGND VPWR VPWR _19313_/X sky130_fd_sc_hd__buf_2
XFILLER_204_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13737_ _13736_/Y _13732_/X VGND VGND VPWR VPWR _13737_/X sky130_fd_sc_hd__or2_4
XFILLER_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_39_0_HCLK clkbuf_5_19_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_79_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__23251__C _23250_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15331__A _15331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16456_ _16456_/A VGND VGND VPWR VPWR _16456_/Y sky130_fd_sc_hd__inv_2
X_19244_ _23805_/Q VGND VGND VPWR VPWR _21607_/B sky130_fd_sc_hd__inv_2
XFILLER_189_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13668_ _11829_/Y _13668_/B VGND VGND VPWR VPWR _13668_/X sky130_fd_sc_hd__or2_4
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15407_ _15139_/Y _15383_/X _15405_/B _15334_/X VGND VGND VPWR VPWR _15407_/X sky130_fd_sc_hd__a211o_4
X_12619_ _12613_/B _12650_/A _12618_/X VGND VGND VPWR VPWR _12620_/A sky130_fd_sc_hd__or3_4
X_19175_ _19174_/Y _19170_/X _19106_/X _19170_/X VGND VGND VPWR VPWR _19175_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16387_ _16387_/A VGND VGND VPWR VPWR _16387_/X sky130_fd_sc_hd__buf_2
X_13599_ _18016_/A VGND VGND VPWR VPWR _17943_/A sky130_fd_sc_hd__buf_2
XFILLER_247_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24793__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18126_ _18126_/A _18126_/B VGND VGND VPWR VPWR _18127_/C sky130_fd_sc_hd__or2_4
X_15338_ _15338_/A _15338_/B _15337_/Y VGND VGND VPWR VPWR _15338_/X sky130_fd_sc_hd__and3_4
XFILLER_247_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24722__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18057_ _18057_/A VGND VGND VPWR VPWR _18128_/A sky130_fd_sc_hd__buf_2
X_15269_ _15269_/A _15269_/B _15268_/X VGND VGND VPWR VPWR _15269_/X sky130_fd_sc_hd__and3_4
XANTENNA__19429__B1 _19360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17008_ _17008_/A _17008_/B _17005_/X _17008_/D VGND VGND VPWR VPWR _17008_/X sky130_fd_sc_hd__or4_4
XANTENNA__21236__B1 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11724__B1 _11721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18959_ _18040_/B VGND VGND VPWR VPWR _18959_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13477__B1 _11786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15506__A _15489_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21970_ _21966_/Y _21967_/X _21968_/X _21969_/X VGND VGND VPWR VPWR _21970_/X sky130_fd_sc_hd__a211o_4
XFILLER_66_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20921_ _24056_/Q _24055_/Q _20921_/C _13637_/D VGND VGND VPWR VPWR _20921_/X sky130_fd_sc_hd__or4_4
XANTENNA__22751__A3 _21312_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25510__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16770__A1_N _15008_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23640_ _23644_/CLK _23640_/D VGND VGND VPWR VPWR _13275_/B sky130_fd_sc_hd__dfxtp_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20852_ _24041_/Q _13644_/X _20862_/B VGND VGND VPWR VPWR _20852_/Y sky130_fd_sc_hd__a21oi_4
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23161__B1 _24284_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23571_ _23525_/CLK _19917_/X VGND VGND VPWR VPWR _19916_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20783_ _20781_/Y _20777_/X _20782_/X VGND VGND VPWR VPWR _20783_/X sky130_fd_sc_hd__o21a_4
XANTENNA__17915__B1 _14608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12865__A _12617_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25310_ _25308_/CLK _25310_/D HRESETn VGND VGND VPWR VPWR _25310_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21711__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22522_ _16694_/Y _22522_/B VGND VGND VPWR VPWR _22522_/X sky130_fd_sc_hd__and2_4
XFILLER_167_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16785__A1_N _15005_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25241_ _25238_/CLK _14056_/X HRESETn VGND VGND VPWR VPWR _13980_/A sky130_fd_sc_hd__dfrtp_4
X_22453_ _15003_/Y _21082_/X _16724_/A _14911_/Y _22452_/X VGND VGND VPWR VPWR _22453_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15941__A2 _15928_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21404_ _14668_/X _19849_/Y VGND VGND VPWR VPWR _21404_/X sky130_fd_sc_hd__or2_4
XFILLER_108_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25172_ _25171_/CLK _14311_/X HRESETn VGND VGND VPWR VPWR _25172_/Q sky130_fd_sc_hd__dfrtp_4
X_22384_ _22380_/X _22383_/X _14666_/X VGND VGND VPWR VPWR _22384_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_163_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24463__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24123_ _23951_/CLK _18890_/X HRESETn VGND VGND VPWR VPWR _24123_/Q sky130_fd_sc_hd__dfstp_4
Xclkbuf_8_59_0_HCLK clkbuf_8_59_0_HCLK/A VGND VGND VPWR VPWR _25260_/CLK sky130_fd_sc_hd__clkbuf_1
X_21335_ _21335_/A _22701_/B VGND VGND VPWR VPWR _21335_/X sky130_fd_sc_hd__or2_4
XFILLER_190_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24054_ _24501_/CLK _24054_/D HRESETn VGND VGND VPWR VPWR _13636_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21266_ _21262_/A _21266_/B VGND VGND VPWR VPWR _21266_/X sky130_fd_sc_hd__or2_4
X_23005_ _23005_/A _23000_/X _23005_/C VGND VGND VPWR VPWR _23006_/D sky130_fd_sc_hd__and3_4
X_20217_ _18203_/B VGND VGND VPWR VPWR _20217_/Y sky130_fd_sc_hd__inv_2
X_21197_ _24212_/Q _21197_/B VGND VGND VPWR VPWR _21199_/B sky130_fd_sc_hd__or2_4
XFILLER_106_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20148_ _20147_/Y _20143_/X _20102_/X _20143_/X VGND VGND VPWR VPWR _20148_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21418__A _21418_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22188__D1 _22187_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12970_ _13087_/A VGND VGND VPWR VPWR _12970_/X sky130_fd_sc_hd__buf_2
X_20079_ _20067_/A VGND VGND VPWR VPWR _20079_/X sky130_fd_sc_hd__buf_2
X_24956_ _24958_/CLK _15464_/X HRESETn VGND VGND VPWR VPWR _24956_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11921_ _11918_/Y _11919_/X _11920_/X _11919_/X VGND VGND VPWR VPWR _11921_/X sky130_fd_sc_hd__a2bb2o_4
X_23907_ _23853_/CLK _23907_/D VGND VGND VPWR VPWR _18953_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_73_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24887_ _23767_/CLK _24887_/D HRESETn VGND VGND VPWR VPWR _24887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_246_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14640_ _18017_/A VGND VGND VPWR VPWR _17949_/A sky130_fd_sc_hd__buf_2
XFILLER_205_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11852_ _11934_/C VGND VGND VPWR VPWR _11852_/Y sky130_fd_sc_hd__inv_2
X_23838_ _23846_/CLK _19154_/X VGND VGND VPWR VPWR _18126_/B sky130_fd_sc_hd__dfxtp_4
XPHY_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14563_/C _14569_/A VGND VGND VPWR VPWR _14571_/X sky130_fd_sc_hd__or2_4
XPHY_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _25522_/Q VGND VGND VPWR VPWR _11783_/Y sky130_fd_sc_hd__inv_2
X_23769_ _24088_/CLK _19346_/X VGND VGND VPWR VPWR _23769_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15994__A1_N _15993_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16310_ _24631_/Q VGND VGND VPWR VPWR _16310_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21702__B2 _22522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13522_ SSn_S2 _13520_/Y _13521_/X _13520_/Y VGND VGND VPWR VPWR _25304_/D sky130_fd_sc_hd__a2bb2o_4
X_25508_ _23406_/CLK _11908_/X HRESETn VGND VGND VPWR VPWR _19970_/A sky130_fd_sc_hd__dfrtp_4
X_17290_ _17183_/Y _17299_/B VGND VGND VPWR VPWR _17290_/X sky130_fd_sc_hd__or2_4
XFILLER_198_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16241_ _16238_/Y _16239_/X _16240_/X _16239_/X VGND VGND VPWR VPWR _16241_/X sky130_fd_sc_hd__a2bb2o_4
X_13453_ _13453_/A VGND VGND VPWR VPWR _14365_/B sky130_fd_sc_hd__buf_2
X_25439_ _25450_/CLK _12480_/X HRESETn VGND VGND VPWR VPWR _25439_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12404_ _12194_/Y _12413_/B VGND VGND VPWR VPWR _12405_/A sky130_fd_sc_hd__or2_4
XFILLER_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16172_ _13577_/B _16171_/X VGND VGND VPWR VPWR _16172_/X sky130_fd_sc_hd__and2_4
X_13384_ _13310_/X _13380_/X _13384_/C VGND VGND VPWR VPWR _13384_/X sky130_fd_sc_hd__or3_4
XFILLER_126_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15123_ _24988_/Q VGND VGND VPWR VPWR _15123_/Y sky130_fd_sc_hd__inv_2
X_12335_ _12335_/A VGND VGND VPWR VPWR _12985_/B sky130_fd_sc_hd__inv_2
XFILLER_147_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24133__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15054_ _15241_/A VGND VGND VPWR VPWR _15165_/A sky130_fd_sc_hd__buf_2
X_19931_ _19931_/A VGND VGND VPWR VPWR _21665_/B sky130_fd_sc_hd__inv_2
X_12266_ _12266_/A _12217_/Y _12266_/C _12184_/Y VGND VGND VPWR VPWR _12271_/C sky130_fd_sc_hd__or4_4
XANTENNA__22712__A _22712_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14005_ _14005_/A _14005_/B VGND VGND VPWR VPWR _14005_/Y sky130_fd_sc_hd__nand2_4
X_19862_ _19856_/Y VGND VGND VPWR VPWR _19862_/X sky130_fd_sc_hd__buf_2
X_12197_ _12197_/A VGND VGND VPWR VPWR _12197_/Y sky130_fd_sc_hd__inv_2
X_18813_ _18787_/A _18786_/X _18724_/X _18811_/B VGND VGND VPWR VPWR _18813_/X sky130_fd_sc_hd__a211o_4
XFILLER_110_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19793_ _13350_/B VGND VGND VPWR VPWR _19793_/Y sky130_fd_sc_hd__inv_2
XANTENNA__25339__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18744_ _18744_/A VGND VGND VPWR VPWR _18752_/A sky130_fd_sc_hd__buf_2
X_15956_ _15924_/X VGND VGND VPWR VPWR _15956_/X sky130_fd_sc_hd__buf_2
XANTENNA__13772__C _13772_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14907_ _15062_/A VGND VGND VPWR VPWR _15219_/A sky130_fd_sc_hd__buf_2
X_15887_ _15958_/A VGND VGND VPWR VPWR _15887_/X sky130_fd_sc_hd__buf_2
X_18675_ _18739_/A VGND VGND VPWR VPWR _18729_/A sky130_fd_sc_hd__inv_2
XFILLER_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17626_ _17625_/X VGND VGND VPWR VPWR _17626_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14838_ _14838_/A VGND VGND VPWR VPWR _14838_/X sky130_fd_sc_hd__buf_2
XFILLER_17_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23143__B1 _23127_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21063__A _22136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14769_ _25059_/Q _14769_/B _14769_/C VGND VGND VPWR VPWR _14769_/X sky130_fd_sc_hd__and3_4
X_17557_ _17602_/B VGND VGND VPWR VPWR _17627_/A sky130_fd_sc_hd__buf_2
XFILLER_189_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24974__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25101__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16508_ _16521_/A VGND VGND VPWR VPWR _16508_/X sky130_fd_sc_hd__buf_2
XFILLER_232_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17488_ _17478_/Y _18356_/B _17480_/X _17487_/X VGND VGND VPWR VPWR _17488_/X sky130_fd_sc_hd__o22a_4
XFILLER_177_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24903__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19227_ _19226_/Y _19224_/X _19203_/X _19224_/X VGND VGND VPWR VPWR _23812_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_177_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15996__A HWDATA[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16439_ _16438_/Y _16370_/A _16361_/X _16370_/A VGND VGND VPWR VPWR _24580_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_8_212_0_HCLK clkbuf_7_106_0_HCLK/X VGND VGND VPWR VPWR _24501_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_192_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19158_ _19158_/A VGND VGND VPWR VPWR _19158_/Y sky130_fd_sc_hd__inv_2
X_18109_ _18220_/A _18109_/B _18108_/X VGND VGND VPWR VPWR _18109_/X sky130_fd_sc_hd__or3_4
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19089_ _19088_/Y _19086_/X _16885_/X _19086_/X VGND VGND VPWR VPWR _23860_/D sky130_fd_sc_hd__a2bb2o_4
X_21120_ _21290_/A VGND VGND VPWR VPWR _21121_/A sky130_fd_sc_hd__buf_2
X_21051_ _21051_/A _21037_/X _21051_/C VGND VGND VPWR VPWR _21051_/X sky130_fd_sc_hd__and3_4
XFILLER_87_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18827__A1_N _16498_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20002_ _23541_/Q VGND VGND VPWR VPWR _21662_/B sky130_fd_sc_hd__inv_2
XFILLER_101_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24810_ _24834_/CLK _15868_/X HRESETn VGND VGND VPWR VPWR _24810_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11764__A HWDATA[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25009__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24741_ _24639_/CLK _16010_/X HRESETn VGND VGND VPWR VPWR _16009_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_28_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21953_ _21949_/X _21952_/X _18301_/A VGND VGND VPWR VPWR _21954_/C sky130_fd_sc_hd__o21a_4
XFILLER_227_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20904_ _24052_/Q _20899_/X _20903_/X VGND VGND VPWR VPWR _20904_/Y sky130_fd_sc_hd__a21oi_4
X_24672_ _24678_/CLK _16201_/X HRESETn VGND VGND VPWR VPWR _23132_/A sky130_fd_sc_hd__dfrtp_4
X_21884_ _21884_/A VGND VGND VPWR VPWR _21913_/A sky130_fd_sc_hd__buf_2
XFILLER_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22069__A _22069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23134__B1 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _23808_/CLK _23623_/D VGND VGND VPWR VPWR _19771_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ _13640_/A _13640_/B _13641_/Y VGND VGND VPWR VPWR _20835_/X sky130_fd_sc_hd__o21a_4
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16067__A _24719_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23554_ _23441_/CLK _19965_/X VGND VGND VPWR VPWR _23554_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_168_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_22_0_HCLK clkbuf_6_23_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_45_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20766_ _20753_/X _20765_/Y _24910_/Q _20757_/X VGND VGND VPWR VPWR _20766_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21160__A2 _14181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24644__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22505_ _16512_/Y _22505_/B VGND VGND VPWR VPWR _22505_/X sky130_fd_sc_hd__and2_4
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23485_ _25510_/CLK _20151_/X VGND VGND VPWR VPWR _23485_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20697_ _13111_/A _13111_/B _13113_/B VGND VGND VPWR VPWR _20697_/X sky130_fd_sc_hd__o21a_4
XFILLER_210_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25224_ _25224_/CLK _25224_/D HRESETn VGND VGND VPWR VPWR _14086_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_195_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22436_ _16144_/Y _21833_/X _22432_/X _11755_/Y _22274_/X VGND VGND VPWR VPWR _22437_/B
+ sky130_fd_sc_hd__o32a_4
XFILLER_108_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25155_ _25158_/CLK _14360_/X HRESETn VGND VGND VPWR VPWR _25155_/Q sky130_fd_sc_hd__dfrtp_4
X_22367_ _22367_/A _19761_/Y VGND VGND VPWR VPWR _22367_/X sky130_fd_sc_hd__or2_4
XANTENNA__18864__B2 _24146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12120_ _12120_/A VGND VGND VPWR VPWR _12120_/Y sky130_fd_sc_hd__inv_2
X_24106_ _24159_/CLK _24106_/D HRESETn VGND VGND VPWR VPWR _12135_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__20671__A1 _14207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21318_ _17203_/X _22543_/A _13110_/A _21317_/X VGND VGND VPWR VPWR _21318_/X sky130_fd_sc_hd__a2bb2o_4
X_25086_ _25098_/CLK _25086_/D HRESETn VGND VGND VPWR VPWR _13560_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22298_ _22298_/A _22298_/B VGND VGND VPWR VPWR _22298_/X sky130_fd_sc_hd__and2_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16662__A1_N _16659_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12051_ _13800_/B VGND VGND VPWR VPWR _21568_/A sky130_fd_sc_hd__buf_2
X_24037_ _24037_/CLK _24037_/D HRESETn VGND VGND VPWR VPWR _13638_/A sky130_fd_sc_hd__dfrtp_4
X_21249_ _21622_/A _21249_/B VGND VGND VPWR VPWR _21249_/X sky130_fd_sc_hd__or2_4
XFILLER_78_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15810_ _11706_/X VGND VGND VPWR VPWR _15810_/X sky130_fd_sc_hd__buf_2
X_16790_ _16789_/Y _16726_/A _16716_/X _16726_/A VGND VGND VPWR VPWR _24446_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15741_ HWDATA[14] VGND VGND VPWR VPWR _15741_/X sky130_fd_sc_hd__buf_2
XANTENNA__23363__A _23363_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12953_ _12947_/B VGND VGND VPWR VPWR _12954_/B sky130_fd_sc_hd__inv_2
X_24939_ _25510_/CLK _15507_/X HRESETn VGND VGND VPWR VPWR _24939_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_246_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_7_104_0_HCLK clkbuf_6_52_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_104_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_11904_ _19970_/A VGND VGND VPWR VPWR _19606_/A sky130_fd_sc_hd__buf_2
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15672_ _15639_/Y _15665_/X _15643_/X _13658_/A _15671_/X VGND VGND VPWR VPWR _15672_/X
+ sky130_fd_sc_hd__a32o_4
X_18460_ _24181_/Q VGND VGND VPWR VPWR _18481_/A sky130_fd_sc_hd__inv_2
XFILLER_206_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12884_ _12796_/A _12884_/B VGND VGND VPWR VPWR _12884_/X sky130_fd_sc_hd__or2_4
XPHY_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14606_/A VGND VGND VPWR VPWR _14623_/Y sky130_fd_sc_hd__inv_2
X_17411_ _21368_/A VGND VGND VPWR VPWR _17411_/X sky130_fd_sc_hd__buf_2
XFILLER_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11825_/X _11835_/B _11831_/X _11834_/X VGND VGND VPWR VPWR _11835_/X sky130_fd_sc_hd__or4_4
X_18391_ _24644_/Q VGND VGND VPWR VPWR _18391_/Y sky130_fd_sc_hd__inv_2
XPHY_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17243_/B VGND VGND VPWR VPWR _17352_/B sky130_fd_sc_hd__buf_2
XPHY_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14554_/A _14554_/B VGND VGND VPWR VPWR _14554_/X sky130_fd_sc_hd__or2_4
XPHY_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11766_/A VGND VGND VPWR VPWR _11766_/X sky130_fd_sc_hd__buf_2
XPHY_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24385__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _12013_/B VGND VGND VPWR VPWR _13506_/A sky130_fd_sc_hd__buf_2
X_17273_ _17273_/A _17273_/B VGND VGND VPWR VPWR _17275_/B sky130_fd_sc_hd__or2_4
XFILLER_186_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _23929_/Q _23928_/Q VGND VGND VPWR VPWR _14485_/X sky130_fd_sc_hd__or2_4
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11697_ _16077_/A VGND VGND VPWR VPWR _11697_/Y sky130_fd_sc_hd__inv_2
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24314__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16224_ _16221_/Y _16223_/X _11726_/X _16223_/X VGND VGND VPWR VPWR _16224_/X sky130_fd_sc_hd__a2bb2o_4
X_19012_ _19010_/Y _19004_/X _18985_/X _19011_/X VGND VGND VPWR VPWR _23888_/D sky130_fd_sc_hd__a2bb2o_4
X_13436_ _13260_/A _13436_/B VGND VGND VPWR VPWR _13436_/X sky130_fd_sc_hd__or2_4
XANTENNA__22100__A1 _24520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_HCLK_A clkbuf_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16155_ _16084_/X VGND VGND VPWR VPWR _16155_/X sky130_fd_sc_hd__buf_2
X_13367_ _13431_/A _13367_/B VGND VGND VPWR VPWR _13367_/X sky130_fd_sc_hd__or2_4
XANTENNA__18855__B2 _24138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15106_ _15106_/A VGND VGND VPWR VPWR _15106_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20662__A1 _14220_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12318_ _25344_/Q VGND VGND VPWR VPWR _13074_/A sky130_fd_sc_hd__inv_2
XFILLER_6_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_42_0_HCLK clkbuf_8_43_0_HCLK/A VGND VGND VPWR VPWR _23665_/CLK sky130_fd_sc_hd__clkbuf_1
X_16086_ _16086_/A VGND VGND VPWR VPWR _16086_/X sky130_fd_sc_hd__buf_2
X_13298_ _13199_/A VGND VGND VPWR VPWR _13431_/A sky130_fd_sc_hd__buf_2
X_15037_ _15037_/A VGND VGND VPWR VPWR _15037_/Y sky130_fd_sc_hd__inv_2
X_19914_ _19914_/A VGND VGND VPWR VPWR _21402_/B sky130_fd_sc_hd__inv_2
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12249_ _12240_/A _12247_/Y _12248_/Y _24768_/Q VGND VGND VPWR VPWR _12249_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16618__B1 _16358_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21058__A _21111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19845_ _21770_/B _19840_/X _19820_/X _19840_/X VGND VGND VPWR VPWR _23598_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13783__B _16721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22445__A1_N _17849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24507__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19776_ _19764_/A VGND VGND VPWR VPWR _19776_/X sky130_fd_sc_hd__buf_2
XANTENNA__25102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16988_ _24390_/Q VGND VGND VPWR VPWR _17103_/A sky130_fd_sc_hd__inv_2
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14644__A2 _14630_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_237_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18727_ _18726_/X VGND VGND VPWR VPWR _24152_/D sky130_fd_sc_hd__inv_2
X_15939_ HWDATA[24] VGND VGND VPWR VPWR _15939_/X sky130_fd_sc_hd__buf_2
XFILLER_92_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__17271__A _17231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18658_ _24146_/Q VGND VGND VPWR VPWR _18658_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__23116__B1 _24283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17609_ _17494_/Y _17597_/B VGND VGND VPWR VPWR _17610_/C sky130_fd_sc_hd__or2_4
XFILLER_52_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18589_ _18589_/A _18593_/A VGND VGND VPWR VPWR _18591_/A sky130_fd_sc_hd__nand2_4
X_20620_ _17399_/X VGND VGND VPWR VPWR _20621_/C sky130_fd_sc_hd__buf_2
XANTENNA__15824__A1_N _12306_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17205__A2_N _17203_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21521__A _21521_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20551_ _20550_/X VGND VGND VPWR VPWR _20551_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24055__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23270_ _16090_/Y _22559_/X _22849_/X _17517_/Y _22821_/B VGND VGND VPWR VPWR _23270_/X
+ sky130_fd_sc_hd__o32a_4
X_20482_ _25207_/Q _20489_/B VGND VGND VPWR VPWR _20482_/X sky130_fd_sc_hd__or2_4
X_22221_ _22221_/A _19809_/Y VGND VGND VPWR VPWR _22221_/X sky130_fd_sc_hd__or2_4
XANTENNA__11759__A _25527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16857__B1 RsRx_S0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22152_ _21439_/X _22151_/X VGND VGND VPWR VPWR _22152_/X sky130_fd_sc_hd__and2_4
X_21103_ _21013_/A _21089_/B VGND VGND VPWR VPWR _21103_/X sky130_fd_sc_hd__and2_4
XANTENNA__17446__A _14364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22083_ _22083_/A _20142_/Y VGND VGND VPWR VPWR _22083_/X sky130_fd_sc_hd__or2_4
XFILLER_121_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16609__B1 _16525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21034_ _22525_/A VGND VGND VPWR VPWR _21034_/X sky130_fd_sc_hd__buf_2
XFILLER_160_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__19271__B2 _19253_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15832__B2 _15786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_216_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22985_ _12272_/Y _22984_/X _24279_/Q _22914_/X VGND VGND VPWR VPWR _22985_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20600__A _20600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24896__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24724_ _24725_/CLK _24724_/D HRESETn VGND VGND VPWR VPWR _16052_/A sky130_fd_sc_hd__dfrtp_4
X_21936_ _21936_/A _19927_/Y VGND VGND VPWR VPWR _21937_/C sky130_fd_sc_hd__or2_4
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24825__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24655_ _24650_/CLK _24655_/D HRESETn VGND VGND VPWR VPWR _24655_/Q sky130_fd_sc_hd__dfrtp_4
X_21867_ _21845_/X _21855_/Y _21859_/X _21867_/D VGND VGND VPWR VPWR _21867_/X sky130_fd_sc_hd__or4_4
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23808_/CLK _23606_/D VGND VGND VPWR VPWR _19819_/A sky130_fd_sc_hd__dfxtp_4
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20818_ _20814_/X VGND VGND VPWR VPWR _20818_/Y sky130_fd_sc_hd__inv_2
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24586_ _24591_/CLK _24586_/D HRESETn VGND VGND VPWR VPWR _15072_/A sky130_fd_sc_hd__dfrtp_4
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21798_ _21661_/A _21798_/B VGND VGND VPWR VPWR _21800_/B sky130_fd_sc_hd__or2_4
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15040__A2_N _24460_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22330__B2 _22181_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23537_ _23415_/CLK _23537_/D VGND VGND VPWR VPWR _23537_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20749_ _20749_/A VGND VGND VPWR VPWR _20749_/Y sky130_fd_sc_hd__inv_2
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16525__A _14407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22881__A2 _21122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _20525_/B VGND VGND VPWR VPWR _20510_/B sky130_fd_sc_hd__buf_2
XFILLER_184_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23468_ _23476_/CLK _23468_/D VGND VGND VPWR VPWR _23468_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ _13220_/X _13221_/B VGND VGND VPWR VPWR _13224_/B sky130_fd_sc_hd__or2_4
X_25207_ _24146_/CLK _14195_/X HRESETn VGND VGND VPWR VPWR _25207_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_195_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22419_ _21748_/A _22419_/B VGND VGND VPWR VPWR _22419_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__22094__B1 _21730_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18837__A1 _24576_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23399_ _25272_/CLK _23399_/D VGND VGND VPWR VPWR _20374_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16848__B1 _16783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12582__B1 _12569_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13152_ _13170_/A _13152_/B VGND VGND VPWR VPWR _13152_/X sky130_fd_sc_hd__or2_4
X_25138_ _25140_/CLK _14420_/X HRESETn VGND VGND VPWR VPWR _25138_/Q sky130_fd_sc_hd__dfstp_4
Xclkbuf_8_1_0_HCLK clkbuf_7_0_0_HCLK/X VGND VGND VPWR VPWR _23476_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_29_0_HCLK clkbuf_7_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_59_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22262__A _22262_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12103_ _12101_/Y _12102_/X _11775_/X _12102_/X VGND VGND VPWR VPWR _12103_/X sky130_fd_sc_hd__a2bb2o_4
X_13083_ _13085_/A _13074_/B _13082_/Y VGND VGND VPWR VPWR _13083_/X sky130_fd_sc_hd__and3_4
X_17960_ _17950_/A _17958_/X _17959_/X VGND VGND VPWR VPWR _17960_/X sky130_fd_sc_hd__and3_4
X_25069_ _25070_/CLK _25069_/D HRESETn VGND VGND VPWR VPWR _13726_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_124_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15520__B1 HADDR[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12034_ _16181_/A VGND VGND VPWR VPWR _13462_/C sky130_fd_sc_hd__buf_2
X_16911_ _24277_/Q VGND VGND VPWR VPWR _16911_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17891_ _17703_/X _17706_/A VGND VGND VPWR VPWR _17892_/A sky130_fd_sc_hd__and2_4
XFILLER_239_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19630_ _18981_/A VGND VGND VPWR VPWR _19630_/X sky130_fd_sc_hd__buf_2
X_16842_ _14885_/Y _16841_/X _16522_/X _16841_/X VGND VGND VPWR VPWR _16842_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19561_ _19561_/A VGND VGND VPWR VPWR _21683_/B sky130_fd_sc_hd__inv_2
XANTENNA__21606__A _22225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13985_ _13979_/C VGND VGND VPWR VPWR _13995_/B sky130_fd_sc_hd__inv_2
X_16773_ _16772_/Y _16769_/X _16518_/X _16769_/X VGND VGND VPWR VPWR _16773_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__20510__A _20510_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13834__B1 _13791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18187__A _18056_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18512_ _18462_/B _18515_/B VGND VGND VPWR VPWR _18516_/B sky130_fd_sc_hd__or2_4
XFILLER_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12936_ _12952_/A _12936_/B _12936_/C VGND VGND VPWR VPWR _25379_/D sky130_fd_sc_hd__and3_4
X_15724_ _15724_/A VGND VGND VPWR VPWR _15724_/X sky130_fd_sc_hd__buf_2
XFILLER_234_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19492_ _21791_/B _19487_/X _11920_/X _19487_/X VGND VGND VPWR VPWR _23718_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_234_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24566__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18443_ _16197_/Y _18459_/A _22939_/A _18442_/Y VGND VGND VPWR VPWR _18443_/X sky130_fd_sc_hd__a2bb2o_4
X_12867_ _12735_/A _12872_/B VGND VGND VPWR VPWR _12867_/X sky130_fd_sc_hd__or2_4
X_15655_ _15671_/A _15773_/B VGND VGND VPWR VPWR _15655_/X sky130_fd_sc_hd__or2_4
XANTENNA__15587__B1 _11715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15051__A2 _15185_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _24237_/Q VGND VGND VPWR VPWR _22584_/A sky130_fd_sc_hd__inv_2
X_14606_ _14606_/A _14605_/X VGND VGND VPWR VPWR _14606_/Y sky130_fd_sc_hd__nand2_4
X_15586_ _24912_/Q VGND VGND VPWR VPWR _22922_/A sky130_fd_sc_hd__inv_2
X_18374_ _18373_/Y VGND VGND VPWR VPWR _18374_/X sky130_fd_sc_hd__buf_2
XANTENNA__20816__A1_N _20690_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12798_ _25385_/Q VGND VGND VPWR VPWR _12838_/B sky130_fd_sc_hd__inv_2
XANTENNA__12253__A1_N _12252_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14536_/X VGND VGND VPWR VPWR _14537_/Y sky130_fd_sc_hd__inv_2
X_17325_ _17325_/A VGND VGND VPWR VPWR _17325_/Y sky130_fd_sc_hd__inv_2
X_11749_ _11746_/Y _11744_/X _11748_/X _11744_/X VGND VGND VPWR VPWR _25531_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_239_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__20332__B1 _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16435__A _19063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ _14468_/A VGND VGND VPWR VPWR _14468_/X sky130_fd_sc_hd__buf_2
X_17256_ _17175_/Y _17256_/B VGND VGND VPWR VPWR _17265_/A sky130_fd_sc_hd__or2_4
X_13419_ _13186_/A _13418_/X _25327_/Q _13184_/A VGND VGND VPWR VPWR _25327_/D sky130_fd_sc_hd__o22a_4
X_16207_ _16207_/A VGND VGND VPWR VPWR _16207_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17187_ _24619_/Q _24348_/Q _16341_/Y _17346_/A VGND VGND VPWR VPWR _17188_/D sky130_fd_sc_hd__o22a_4
XANTENNA__19746__A HWDATA[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14399_ HWDATA[7] VGND VGND VPWR VPWR _14400_/A sky130_fd_sc_hd__buf_2
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16839__B1 _16601_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16138_ _22564_/A VGND VGND VPWR VPWR _16138_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25354__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16069_ _24718_/Q VGND VGND VPWR VPWR _16069_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16170__A _14764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20399__B1 _15764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19828_ _21384_/B _19823_/X _19827_/X _19823_/X VGND VGND VPWR VPWR _23604_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19481__A _19480_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19759_ _19646_/A VGND VGND VPWR VPWR _19759_/X sky130_fd_sc_hd__buf_2
XFILLER_204_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13825__B1 _13824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22770_ _21022_/A VGND VGND VPWR VPWR _23043_/A sky130_fd_sc_hd__buf_2
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22560__B2 _22559_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21721_ _14256_/Y _21721_/B VGND VGND VPWR VPWR _21721_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15233__B _15311_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18825__A pwm_S7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24236__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24440_ _24460_/CLK _16805_/X HRESETn VGND VGND VPWR VPWR _24440_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21652_ _21652_/A VGND VGND VPWR VPWR _21652_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_5_10_0_HCLK_A clkbuf_4_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14250__B1 _13826_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22347__A _21936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21115__A2 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20603_ _20603_/A _20603_/B _20602_/Y VGND VGND VPWR VPWR _20603_/X sky130_fd_sc_hd__and3_4
XANTENNA__21251__A _21627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24371_ _24641_/CLK _24371_/D HRESETn VGND VGND VPWR VPWR _24371_/Q sky130_fd_sc_hd__dfrtp_4
X_21583_ _21583_/A VGND VGND VPWR VPWR _21741_/B sky130_fd_sc_hd__buf_2
XANTENNA__20323__B1 _11788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23322_ _12167_/A _21077_/X _23320_/X _23321_/X _22876_/C VGND VGND VPWR VPWR _23322_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_166_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20534_ _24072_/Q _20528_/X _20501_/B _20533_/X VGND VGND VPWR VPWR _24072_/D sky130_fd_sc_hd__a211o_4
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23253_ _23253_/A _22817_/B _22817_/C VGND VGND VPWR VPWR _23253_/X sky130_fd_sc_hd__and3_4
X_20465_ _14054_/A _20465_/B VGND VGND VPWR VPWR _20468_/C sky130_fd_sc_hd__and2_4
XFILLER_193_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18560__A _18560_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22204_ _22223_/A _22204_/B _22204_/C VGND VGND VPWR VPWR _22204_/X sky130_fd_sc_hd__and3_4
XANTENNA__20626__A1 _15465_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23184_ _23184_/A _22658_/B VGND VGND VPWR VPWR _23184_/X sky130_fd_sc_hd__or2_4
XFILLER_161_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20396_ _13294_/B VGND VGND VPWR VPWR _20396_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22135_ _21303_/A _22135_/B _22135_/C VGND VGND VPWR VPWR _22135_/X sky130_fd_sc_hd__and3_4
XANTENNA__15502__B1 HADDR[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25024__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22066_ _22385_/A _22066_/B VGND VGND VPWR VPWR _22066_/X sky130_fd_sc_hd__or2_4
XFILLER_87_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21017_ _25334_/Q _21017_/B VGND VGND VPWR VPWR _21017_/X sky130_fd_sc_hd__and2_4
XFILLER_248_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13816__B1 _11748_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13770_ _13769_/Y VGND VGND VPWR VPWR _13771_/A sky130_fd_sc_hd__buf_2
X_22968_ _22968_/A _22897_/X VGND VGND VPWR VPWR _22968_/X sky130_fd_sc_hd__or2_4
XANTENNA__21354__A2 _14182_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12721_ _12717_/A _12721_/B VGND VGND VPWR VPWR _12721_/Y sky130_fd_sc_hd__nand2_4
XFILLER_231_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21919_ _17720_/A _21919_/B VGND VGND VPWR VPWR _21919_/X sky130_fd_sc_hd__or2_4
X_24707_ _24639_/CLK _16100_/X HRESETn VGND VGND VPWR VPWR _23157_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_204_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22899_ _22474_/X _22898_/X _22858_/X _24839_/Q _22478_/X VGND VGND VPWR VPWR _22899_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15440_ _13931_/B _15432_/X _15427_/X _13931_/A _15439_/X VGND VGND VPWR VPWR _15440_/X
+ sky130_fd_sc_hd__a32o_4
X_12652_ _12680_/A VGND VGND VPWR VPWR _12677_/A sky130_fd_sc_hd__buf_2
X_24638_ _24639_/CLK _24638_/D HRESETn VGND VGND VPWR VPWR _16291_/A sky130_fd_sc_hd__dfrtp_4
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21546__A1_N _17242_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _15125_/Y _15347_/B _15313_/A _15369_/B VGND VGND VPWR VPWR _15371_/X sky130_fd_sc_hd__a211o_4
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _25407_/Q VGND VGND VPWR VPWR _12693_/A sky130_fd_sc_hd__inv_2
X_24569_ _24573_/CLK _24569_/D HRESETn VGND VGND VPWR VPWR _24569_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19180__B1 _19067_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14322_ _12149_/X _18372_/D VGND VGND VPWR VPWR _14324_/B sky130_fd_sc_hd__or2_4
X_17110_ _17098_/B VGND VGND VPWR VPWR _17111_/B sky130_fd_sc_hd__inv_2
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18090_ _18090_/A VGND VGND VPWR VPWR _18094_/A sky130_fd_sc_hd__buf_2
XFILLER_184_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__23959__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17041_ _16991_/Y _17039_/Y _17041_/C _17040_/Y VGND VGND VPWR VPWR _17042_/C sky130_fd_sc_hd__or4_4
XFILLER_156_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ _14251_/Y _14247_/X _13829_/X _14252_/X VGND VGND VPWR VPWR _14253_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_109_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13204_ _13288_/A VGND VGND VPWR VPWR _13365_/A sky130_fd_sc_hd__buf_2
XANTENNA__20617__A1 _14863_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23088__A _24604_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14184_ _14184_/A _14183_/X VGND VGND VPWR VPWR _14187_/B sky130_fd_sc_hd__or2_4
XFILLER_125_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13135_ _13225_/A VGND VGND VPWR VPWR _13167_/A sky130_fd_sc_hd__buf_2
XFILLER_152_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18992_ _18154_/B VGND VGND VPWR VPWR _18992_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13066_ _13065_/X VGND VGND VPWR VPWR _25347_/D sky130_fd_sc_hd__inv_2
X_17943_ _17943_/A _19162_/A VGND VGND VPWR VPWR _17945_/B sky130_fd_sc_hd__or2_4
XANTENNA__23031__A2 _23029_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_116_0_HCLK clkbuf_7_58_0_HCLK/X VGND VGND VPWR VPWR _24874_/CLK sky130_fd_sc_hd__clkbuf_1
X_12017_ _25494_/Q VGND VGND VPWR VPWR _12017_/Y sky130_fd_sc_hd__inv_2
X_17874_ _17866_/A _17874_/B _17873_/Y VGND VGND VPWR VPWR _17874_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_179_0_HCLK clkbuf_7_89_0_HCLK/X VGND VGND VPWR VPWR _25134_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__18994__B1 _18948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19613_ _19613_/A VGND VGND VPWR VPWR _19613_/X sky130_fd_sc_hd__buf_2
XANTENNA__24747__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16825_ _16824_/Y _16822_/X _15739_/X _16822_/X VGND VGND VPWR VPWR _16825_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_226_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21336__A _21232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19544_ _19542_/Y _19539_/X _19543_/X _19539_/X VGND VGND VPWR VPWR _19544_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_235_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15334__A _15282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16756_ _14998_/Y _16755_/X _15735_/X _16755_/X VGND VGND VPWR VPWR _24462_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13968_ _13991_/D VGND VGND VPWR VPWR _14007_/B sky130_fd_sc_hd__buf_2
XFILLER_80_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14480__B1 _14479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22542__A1 _21284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15707_ _15706_/X VGND VGND VPWR VPWR _15707_/X sky130_fd_sc_hd__buf_2
X_12919_ _12617_/B _12835_/X VGND VGND VPWR VPWR _12919_/X sky130_fd_sc_hd__or2_4
X_19475_ _19874_/A VGND VGND VPWR VPWR _19475_/X sky130_fd_sc_hd__buf_2
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13899_ _13917_/B VGND VGND VPWR VPWR _13907_/C sky130_fd_sc_hd__inv_2
X_16687_ _24491_/Q VGND VGND VPWR VPWR _16687_/Y sky130_fd_sc_hd__inv_2
X_18426_ _24175_/Q VGND VGND VPWR VPWR _18467_/B sky130_fd_sc_hd__inv_2
XFILLER_62_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15638_ _14366_/A _22829_/A VGND VGND VPWR VPWR _15671_/A sky130_fd_sc_hd__or2_4
X_18357_ _18356_/X VGND VGND VPWR VPWR _18357_/Y sky130_fd_sc_hd__inv_2
X_15569_ _24918_/Q VGND VGND VPWR VPWR _15569_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22845__A2 _22828_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19171__B1 _19125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17308_ _17310_/B VGND VGND VPWR VPWR _17309_/B sky130_fd_sc_hd__inv_2
XFILLER_147_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18288_ _18288_/A _17704_/X VGND VGND VPWR VPWR _18288_/X sky130_fd_sc_hd__or2_4
XANTENNA__25535__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17721__B2 _21473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17239_ _17239_/A VGND VGND VPWR VPWR _17240_/D sky130_fd_sc_hd__inv_2
XANTENNA__15732__B1 _11715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13504__A1_N _13503_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20250_ _23447_/Q VGND VGND VPWR VPWR _20250_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23270__A2 _22559_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20415__A _20409_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20181_ _20177_/Y _20180_/X _20089_/X _20180_/X VGND VGND VPWR VPWR _23474_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__23007__C1 _23006_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_12_0_HCLK clkbuf_6_6_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_12_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_7_75_0_HCLK clkbuf_7_75_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_75_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__22630__A _24797_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23940_ _23938_/CLK _23940_/D HRESETn VGND VGND VPWR VPWR _20558_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_215_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24488__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21246__A _21627_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23871_ _23735_/CLK _23871_/D VGND VGND VPWR VPWR _23871_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_217_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20150__A _20137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24417__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22822_ _24733_/Q _21061_/X _21062_/X _22821_/X VGND VGND VPWR VPWR _22822_/X sky130_fd_sc_hd__a211o_4
XFILLER_84_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14471__B1 _14380_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_HCLK_A clkbuf_2_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25541_ _24626_/CLK _25541_/D HRESETn VGND VGND VPWR VPWR _25541_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_241_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22753_ _22753_/A _22638_/B VGND VGND VPWR VPWR _22753_/X sky130_fd_sc_hd__or2_4
XFILLER_25_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21704_ _24751_/Q _23172_/A VGND VGND VPWR VPWR _21704_/X sky130_fd_sc_hd__or2_4
X_25472_ _25471_/CLK _12105_/X HRESETn VGND VGND VPWR VPWR _25472_/Q sky130_fd_sc_hd__dfrtp_4
X_22684_ _22684_/A _22684_/B VGND VGND VPWR VPWR _22684_/X sky130_fd_sc_hd__and2_4
XANTENNA__14223__B1 _13788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24423_ _24419_/CLK _16838_/X HRESETn VGND VGND VPWR VPWR _24423_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21635_ _22380_/A _21633_/X _21635_/C VGND VGND VPWR VPWR _21635_/X sky130_fd_sc_hd__and3_4
XFILLER_212_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15971__B1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24354_ _24346_/CLK _17338_/X HRESETn VGND VGND VPWR VPWR _17336_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_100_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21566_ _16261_/Y _16180_/A _15110_/A _16719_/A VGND VGND VPWR VPWR _21567_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20311__A3 _11760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23305_ _23182_/A _23296_/Y _23305_/C _23305_/D VGND VGND VPWR VPWR _23305_/X sky130_fd_sc_hd__or4_4
XFILLER_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20517_ _20517_/A _20517_/B _20496_/A _20503_/C VGND VGND VPWR VPWR _20517_/X sky130_fd_sc_hd__and4_4
XANTENNA__19386__A _17955_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24285_ _24278_/CLK _17790_/X HRESETn VGND VGND VPWR VPWR _24285_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15723__B1 _11688_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21497_ _21803_/A _21495_/X _21496_/X VGND VGND VPWR VPWR _21497_/X sky130_fd_sc_hd__and3_4
XANTENNA__25205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16803__A _24440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23236_ _20810_/A _22992_/X _20948_/Y _22794_/X VGND VGND VPWR VPWR _23236_/X sky130_fd_sc_hd__o22a_4
X_20448_ _14053_/A _20435_/X _20439_/Y _20447_/X VGND VGND VPWR VPWR _20448_/X sky130_fd_sc_hd__a211o_4
XFILLER_181_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23167_ _23235_/A _23167_/B VGND VGND VPWR VPWR _23167_/Y sky130_fd_sc_hd__nor2_4
X_20379_ _20372_/X _20368_/X _18257_/X _23397_/Q _20370_/X VGND VGND VPWR VPWR _20379_/X
+ sky130_fd_sc_hd__a32o_4
X_22118_ _21111_/A _22114_/X _22117_/X VGND VGND VPWR VPWR _22118_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23098_ _23097_/X VGND VGND VPWR VPWR _23098_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14940_ _14940_/A VGND VGND VPWR VPWR _14940_/Y sky130_fd_sc_hd__inv_2
X_22049_ _22046_/Y _22047_/X _21969_/X _22048_/X VGND VGND VPWR VPWR _23342_/B sky130_fd_sc_hd__a211o_4
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24840__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14871_ _24952_/Q VGND VGND VPWR VPWR _14871_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24158__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16610_ _16610_/A VGND VGND VPWR VPWR _16610_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13822_ _13832_/A VGND VGND VPWR VPWR _13822_/X sky130_fd_sc_hd__buf_2
X_17590_ _17590_/A _17587_/X VGND VGND VPWR VPWR _17590_/X sky130_fd_sc_hd__or2_4
XFILLER_232_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23371__A _23371_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13753_ _14683_/A VGND VGND VPWR VPWR _13753_/X sky130_fd_sc_hd__buf_2
X_16541_ _16547_/A VGND VGND VPWR VPWR _16541_/X sky130_fd_sc_hd__buf_2
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12704_ _12704_/A _12707_/B VGND VGND VPWR VPWR _12705_/C sky130_fd_sc_hd__nand2_4
XFILLER_188_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19260_ _22066_/B _19254_/X _16869_/X _19259_/X VGND VGND VPWR VPWR _19260_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13684_ _13663_/Y _13667_/X _13680_/X _25296_/Q _13683_/Y VGND VGND VPWR VPWR _25296_/D
+ sky130_fd_sc_hd__a32o_4
X_16472_ _16472_/A VGND VGND VPWR VPWR _16472_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14214__B1 _13824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18211_ _17968_/X _18209_/X _18210_/X VGND VGND VPWR VPWR _18211_/X sky130_fd_sc_hd__and3_4
X_12635_ _12608_/X _12626_/D _12512_/Y VGND VGND VPWR VPWR _12636_/C sky130_fd_sc_hd__o21a_4
X_15423_ _15423_/A _15422_/Y VGND VGND VPWR VPWR _15424_/B sky130_fd_sc_hd__or2_4
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19191_ _19191_/A VGND VGND VPWR VPWR _19191_/X sky130_fd_sc_hd__buf_2
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15962__B1 _24760_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15354_ _15353_/X VGND VGND VPWR VPWR _24996_/D sky130_fd_sc_hd__inv_2
X_18142_ _18027_/A _23749_/Q VGND VGND VPWR VPWR _18144_/B sky130_fd_sc_hd__or2_4
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ _12566_/A _12561_/X _12563_/X _12566_/D VGND VGND VPWR VPWR _12587_/B sky130_fd_sc_hd__or4_4
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14305_ _14295_/X _14304_/X _25321_/Q _14300_/X VGND VGND VPWR VPWR _14305_/X sky130_fd_sc_hd__o22a_4
XFILLER_172_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15285_ _15285_/A VGND VGND VPWR VPWR _15285_/Y sky130_fd_sc_hd__inv_2
X_18073_ _17985_/X _18073_/B VGND VGND VPWR VPWR _18073_/X sky130_fd_sc_hd__or2_4
X_12497_ _12263_/A _12456_/X _12497_/C VGND VGND VPWR VPWR _25433_/D sky130_fd_sc_hd__and3_4
XFILLER_156_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14236_ _13929_/Y _13938_/X _13949_/Y _14236_/D VGND VGND VPWR VPWR _14236_/X sky130_fd_sc_hd__or4_4
X_17024_ _17024_/A VGND VGND VPWR VPWR _17045_/A sky130_fd_sc_hd__inv_2
XFILLER_125_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23249__C _23075_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24999__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14167_ _14162_/A _14161_/X _14162_/Y VGND VGND VPWR VPWR _14167_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__15329__A _15282_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13118_ _13118_/A _13117_/X VGND VGND VPWR VPWR _13119_/B sky130_fd_sc_hd__or2_4
XANTENNA__24928__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14098_ _14115_/A VGND VGND VPWR VPWR _14099_/A sky130_fd_sc_hd__inv_2
X_18975_ _19411_/A _19141_/B _13615_/A _13596_/A VGND VGND VPWR VPWR _18975_/X sky130_fd_sc_hd__or4_4
XFILLER_67_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13049_ _13046_/A _13046_/B VGND VGND VPWR VPWR _13050_/C sky130_fd_sc_hd__nand2_4
X_17926_ _17926_/A _17917_/B VGND VGND VPWR VPWR _17926_/X sky130_fd_sc_hd__or2_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22763__A1 _12801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18967__B1 _18965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24581__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17857_ _17747_/Y _17854_/X VGND VGND VPWR VPWR _17858_/C sky130_fd_sc_hd__or2_4
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__17176__A1_N _24633_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24510__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15064__A _15059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16808_ _16799_/A VGND VGND VPWR VPWR _16808_/X sky130_fd_sc_hd__buf_2
XFILLER_242_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17788_ _24285_/Q _17787_/Y VGND VGND VPWR VPWR _17790_/B sky130_fd_sc_hd__or2_4
XFILLER_226_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14453__B1 _14392_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19527_ _19521_/Y _19526_/X _19414_/X _19526_/X VGND VGND VPWR VPWR _19527_/X sky130_fd_sc_hd__a2bb2o_4
X_16739_ _16730_/A VGND VGND VPWR VPWR _16739_/X sky130_fd_sc_hd__buf_2
X_19458_ _19457_/Y VGND VGND VPWR VPWR _19458_/X sky130_fd_sc_hd__buf_2
XFILLER_50_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15548__A3 _15545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18409_ _18409_/A VGND VGND VPWR VPWR _18409_/Y sky130_fd_sc_hd__inv_2
X_19389_ _19388_/Y VGND VGND VPWR VPWR _19389_/X sky130_fd_sc_hd__buf_2
XFILLER_148_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14408__A _14408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_194_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21420_ _22466_/A VGND VGND VPWR VPWR _21421_/A sky130_fd_sc_hd__buf_2
XANTENNA__20829__B2 _20828_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21351_ _14209_/A VGND VGND VPWR VPWR _21351_/X sky130_fd_sc_hd__buf_2
XFILLER_163_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20302_ _20302_/A VGND VGND VPWR VPWR _21482_/B sky130_fd_sc_hd__inv_2
X_24070_ _25346_/CLK _24070_/D HRESETn VGND VGND VPWR VPWR HREADYOUT sky130_fd_sc_hd__dfstp_4
X_21282_ _21281_/B _21280_/X _21178_/X _21281_/Y VGND VGND VPWR VPWR _21282_/X sky130_fd_sc_hd__a211o_4
XANTENNA__17438__B _17438_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23243__A2 _22661_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15720__A3 _15719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23021_ _23021_/A VGND VGND VPWR VPWR _23021_/Y sky130_fd_sc_hd__inv_2
X_20233_ _13360_/B VGND VGND VPWR VPWR _20233_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24669__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20164_ _20158_/Y VGND VGND VPWR VPWR _20164_/X sky130_fd_sc_hd__buf_2
XFILLER_226_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16130__B1 _11735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20095_ _24411_/Q VGND VGND VPWR VPWR _20095_/X sky130_fd_sc_hd__buf_2
X_24972_ _24973_/CLK _15437_/X HRESETn VGND VGND VPWR VPWR _13922_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18958__B1 _17418_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23923_ _23927_/CLK _23923_/D HRESETn VGND VGND VPWR VPWR _20994_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_85_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_162_0_HCLK clkbuf_7_81_0_HCLK/X VGND VGND VPWR VPWR _24889_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__24251__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_5_0_HCLK clkbuf_7_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_5_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_23854_ _23735_/CLK _23854_/D VGND VGND VPWR VPWR _23854_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_242_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_19_0_HCLK clkbuf_7_9_0_HCLK/X VGND VGND VPWR VPWR _23675_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_217_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14444__B1 _14400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22805_ _22844_/A _22800_/X _22804_/X VGND VGND VPWR VPWR _22811_/C sky130_fd_sc_hd__and3_4
XFILLER_214_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21704__A _24751_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23785_ _23785_/CLK _23785_/D VGND VGND VPWR VPWR _23785_/Q sky130_fd_sc_hd__dfxtp_4
X_20997_ _20997_/A VGND VGND VPWR VPWR _20998_/B sky130_fd_sc_hd__inv_2
XFILLER_25_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__19383__B1 _19360_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22736_ _22515_/X _22734_/X _21956_/A _22735_/X VGND VGND VPWR VPWR _22736_/X sky130_fd_sc_hd__o22a_4
X_25524_ _25524_/CLK _11776_/X HRESETn VGND VGND VPWR VPWR _11772_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_213_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15702__A HWDATA[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25455_ _25453_/CLK _12416_/Y HRESETn VGND VGND VPWR VPWR _12240_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22667_ _22667_/A _22572_/X VGND VGND VPWR VPWR _22669_/B sky130_fd_sc_hd__or2_4
XFILLER_240_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12420_ _12274_/X _12428_/D VGND VGND VPWR VPWR _12420_/X sky130_fd_sc_hd__or2_4
X_24406_ _23859_/CLK _16886_/X HRESETn VGND VGND VPWR VPWR _19852_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13222__A _13199_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21618_ _14753_/X _21618_/B VGND VGND VPWR VPWR _21618_/X sky130_fd_sc_hd__or2_4
X_25386_ _25387_/CLK _25386_/D HRESETn VGND VGND VPWR VPWR _25386_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22598_ _21294_/X _22597_/X _21300_/A _24831_/Q _22490_/X VGND VGND VPWR VPWR _22598_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_224_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12351_ _12351_/A VGND VGND VPWR VPWR _13069_/A sky130_fd_sc_hd__inv_2
X_24337_ _24340_/CLK _24337_/D HRESETn VGND VGND VPWR VPWR _21000_/A sky130_fd_sc_hd__dfstp_4
X_21549_ _14474_/Y _14246_/A VGND VGND VPWR VPWR _21549_/X sky130_fd_sc_hd__or2_4
XFILLER_181_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15070_ _15070_/A VGND VGND VPWR VPWR _15070_/Y sky130_fd_sc_hd__inv_2
X_12282_ _12282_/A VGND VGND VPWR VPWR _12993_/A sky130_fd_sc_hd__inv_2
X_24268_ _24266_/CLK _24268_/D HRESETn VGND VGND VPWR VPWR _24268_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15711__A3 _15710_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14021_ _14012_/A VGND VGND VPWR VPWR _14021_/Y sky130_fd_sc_hd__inv_2
X_23219_ _23219_/A _23040_/X VGND VGND VPWR VPWR _23219_/X sky130_fd_sc_hd__or2_4
XANTENNA__11677__A _11700_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24199_ _24199_/CLK _24199_/D HRESETn VGND VGND VPWR VPWR _18354_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_134_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22993__B2 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16121__B1 _15953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23366__A _21013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22783__A1_N _17314_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18760_ _18760_/A _18764_/B VGND VGND VPWR VPWR _18761_/C sky130_fd_sc_hd__nand2_4
X_15972_ _15930_/Y VGND VGND VPWR VPWR _15972_/X sky130_fd_sc_hd__buf_2
XFILLER_95_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18949__B1 _18948_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17711_ _19455_/A VGND VGND VPWR VPWR _17711_/Y sky130_fd_sc_hd__inv_2
X_14923_ _25027_/Q _14922_/A _14921_/X _14922_/Y VGND VGND VPWR VPWR _14923_/X sky130_fd_sc_hd__o22a_4
X_18691_ _18689_/Y _18691_/B _18613_/A _18658_/Y VGND VGND VPWR VPWR _18694_/C sky130_fd_sc_hd__or4_4
X_17642_ _17648_/A _17648_/B VGND VGND VPWR VPWR _17643_/B sky130_fd_sc_hd__or2_4
X_14854_ _14854_/A VGND VGND VPWR VPWR _14854_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13805_ _13804_/Y VGND VGND VPWR VPWR _21642_/A sky130_fd_sc_hd__buf_2
XFILLER_223_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17573_ _24303_/Q VGND VGND VPWR VPWR _17582_/B sky130_fd_sc_hd__inv_2
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11997_ _13490_/A _11996_/Y _13490_/A _11996_/Y VGND VGND VPWR VPWR _11997_/X sky130_fd_sc_hd__a2bb2o_4
X_14785_ _18082_/A _14784_/Y _25078_/Q _14784_/A VGND VGND VPWR VPWR _14785_/X sky130_fd_sc_hd__o22a_4
XFILLER_189_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19312_ _18138_/B VGND VGND VPWR VPWR _19312_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15532__A1_N _12086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16524_ _24552_/Q VGND VGND VPWR VPWR _16524_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13736_ _13736_/A VGND VGND VPWR VPWR _13736_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16188__B1 _15554_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19243_ _19242_/Y _19238_/X _16878_/X _19238_/X VGND VGND VPWR VPWR _23806_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_231_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16455_ _16450_/Y _16454_/X _15545_/X _16454_/X VGND VGND VPWR VPWR _16455_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13667_ _13666_/Y VGND VGND VPWR VPWR _13667_/X sky130_fd_sc_hd__buf_2
XFILLER_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25127__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15406_ _15385_/X _15405_/X _15402_/X VGND VGND VPWR VPWR _24981_/D sky130_fd_sc_hd__and3_4
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12618_ _12610_/X _12626_/D _12580_/Y VGND VGND VPWR VPWR _12618_/X sky130_fd_sc_hd__o21a_4
X_19174_ _23830_/Q VGND VGND VPWR VPWR _19174_/Y sky130_fd_sc_hd__inv_2
X_13598_ _18057_/A VGND VGND VPWR VPWR _18016_/A sky130_fd_sc_hd__buf_2
X_16386_ HWDATA[24] VGND VGND VPWR VPWR _16386_/X sky130_fd_sc_hd__buf_2
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18125_ _18125_/A _23846_/Q VGND VGND VPWR VPWR _18127_/B sky130_fd_sc_hd__or2_4
X_12549_ _25418_/Q _12547_/Y _12692_/A _12551_/A VGND VGND VPWR VPWR _12549_/X sky130_fd_sc_hd__a2bb2o_4
X_15337_ _15333_/A _15333_/B VGND VGND VPWR VPWR _15337_/Y sky130_fd_sc_hd__nand2_4
XFILLER_247_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22681__B1 _22696_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12971__A _24781_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18056_ _18056_/A _18056_/B _18056_/C VGND VGND VPWR VPWR _18056_/X sky130_fd_sc_hd__and3_4
XFILLER_172_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15268_ _25013_/Q _15268_/B VGND VGND VPWR VPWR _15268_/X sky130_fd_sc_hd__or2_4
XANTENNA__17258__B _17231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17007_ _24738_/Q _17006_/Y _16022_/Y _24393_/Q VGND VGND VPWR VPWR _17008_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14219_ _14217_/Y _14213_/X _13829_/X _14218_/X VGND VGND VPWR VPWR _14219_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22433__B1 _16052_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19754__A _19740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15199_ _15165_/A _15188_/X _15199_/C VGND VGND VPWR VPWR _25031_/D sky130_fd_sc_hd__and3_4
XANTENNA__24762__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16112__B1 _16020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18958_ _18957_/Y _14654_/X _17418_/X _14654_/X VGND VGND VPWR VPWR _18958_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24009__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17909_ _17901_/Y _17908_/A _17907_/X _17893_/A _17908_/Y VGND VGND VPWR VPWR _24256_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_100_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18889_ _18871_/X _18885_/X _24123_/Q _20984_/A _18888_/X VGND VGND VPWR VPWR _18889_/X
+ sky130_fd_sc_hd__a32o_4
X_20920_ _24056_/Q VGND VGND VPWR VPWR _20920_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_235_0_HCLK clkbuf_8_234_0_HCLK/A VGND VGND VPWR VPWR _23986_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_212_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20851_ _20857_/B VGND VGND VPWR VPWR _20862_/B sky130_fd_sc_hd__inv_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23570_ _23559_/CLK _19921_/X VGND VGND VPWR VPWR _23570_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20782_ _20781_/A _13108_/B _20754_/X _13108_/D VGND VGND VPWR VPWR _20782_/X sky130_fd_sc_hd__or4_4
XANTENNA__21172__B1 _11701_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22521_ _22518_/X _22521_/B VGND VGND VPWR VPWR _22521_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__18427__A1_N _22814_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25240_ _25238_/CLK _14057_/X HRESETn VGND VGND VPWR VPWR _25240_/Q sky130_fd_sc_hd__dfrtp_4
X_22452_ _23075_/B VGND VGND VPWR VPWR _22452_/X sky130_fd_sc_hd__buf_2
XFILLER_148_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15941__A3 HWDATA[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21403_ _14681_/A _21401_/X _21403_/C VGND VGND VPWR VPWR _21403_/X sky130_fd_sc_hd__and3_4
X_25171_ _25171_/CLK _25171_/D HRESETn VGND VGND VPWR VPWR _25171_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22383_ _22383_/A _22381_/X _22383_/C VGND VGND VPWR VPWR _22383_/X sky130_fd_sc_hd__and3_4
XFILLER_148_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22672__B1 _21582_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18340__A1 _18900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16353__A _14392_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24122_ _23951_/CLK _24122_/D HRESETn VGND VGND VPWR VPWR _20984_/B sky130_fd_sc_hd__dfstp_4
X_21334_ _21323_/A VGND VGND VPWR VPWR _22701_/B sky130_fd_sc_hd__buf_2
XANTENNA__16351__B1 _16349_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24053_ _24501_/CLK _20909_/X HRESETn VGND VGND VPWR VPWR _24053_/Q sky130_fd_sc_hd__dfrtp_4
X_21265_ _21261_/X _21264_/X _21247_/X VGND VGND VPWR VPWR _21265_/X sky130_fd_sc_hd__o21a_4
XFILLER_190_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23004_ _24435_/Q _22807_/X _23001_/X _23003_/X VGND VGND VPWR VPWR _23005_/C sky130_fd_sc_hd__a211o_4
X_20216_ _20215_/Y _20213_/X _19711_/X _20213_/X VGND VGND VPWR VPWR _20216_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21196_ _18314_/A _21187_/X _21195_/X VGND VGND VPWR VPWR _21196_/X sky130_fd_sc_hd__or3_4
XANTENNA__24432__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20147_ _23486_/Q VGND VGND VPWR VPWR _20147_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_45_0_HCLK clkbuf_6_45_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_91_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20078_ _23509_/Q VGND VGND VPWR VPWR _21637_/B sky130_fd_sc_hd__inv_2
X_24955_ _24958_/CLK _15467_/X HRESETn VGND VGND VPWR VPWR _15465_/A sky130_fd_sc_hd__dfstp_4
XFILLER_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11920_ _19613_/A VGND VGND VPWR VPWR _11920_/X sky130_fd_sc_hd__buf_2
X_23906_ _23875_/CLK _23906_/D VGND VGND VPWR VPWR _17959_/B sky130_fd_sc_hd__dfxtp_4
X_24886_ _24886_/CLK _15708_/X HRESETn VGND VGND VPWR VPWR _24886_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11851_ _11934_/C _11850_/Y VGND VGND VPWR VPWR _11851_/X sky130_fd_sc_hd__or2_4
X_23837_ _23846_/CLK _19157_/X VGND VGND VPWR VPWR _18158_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_205_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16528__A _16453_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14570_/A _14570_/B VGND VGND VPWR VPWR _14570_/X sky130_fd_sc_hd__or2_4
XPHY_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _11777_/Y _11778_/X _11781_/X _11778_/X VGND VGND VPWR VPWR _25523_/D sky130_fd_sc_hd__a2bb2o_4
X_23768_ _24088_/CLK _19349_/X VGND VGND VPWR VPWR _23768_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_202_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21163__B1 _17438_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_HCLK clkbuf_3_0_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_1_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _14262_/A VGND VGND VPWR VPWR _13521_/X sky130_fd_sc_hd__buf_2
X_25507_ _23406_/CLK _11912_/X HRESETn VGND VGND VPWR VPWR _19974_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_198_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22719_ _22275_/X VGND VGND VPWR VPWR _22719_/X sky130_fd_sc_hd__buf_2
XPHY_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23699_ _23706_/CLK _23699_/D VGND VGND VPWR VPWR _23699_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__25220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13452_ _25325_/Q VGND VGND VPWR VPWR _13452_/Y sky130_fd_sc_hd__inv_2
X_16240_ _16240_/A VGND VGND VPWR VPWR _16240_/X sky130_fd_sc_hd__buf_2
X_25438_ _25450_/CLK _12483_/X HRESETn VGND VGND VPWR VPWR _12217_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__16590__B1 _16236_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22265__A _21954_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ _12232_/Y _12402_/X VGND VGND VPWR VPWR _12413_/B sky130_fd_sc_hd__or2_4
X_13383_ _13314_/X _13383_/B _13382_/X VGND VGND VPWR VPWR _13384_/C sky130_fd_sc_hd__and3_4
X_16171_ _14765_/A _14775_/A VGND VGND VPWR VPWR _16171_/X sky130_fd_sc_hd__and2_4
X_25369_ _25369_/CLK _12965_/X HRESETn VGND VGND VPWR VPWR _25369_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ _12982_/A _12332_/Y _25340_/Q _12333_/Y VGND VGND VPWR VPWR _12334_/X sky130_fd_sc_hd__a2bb2o_4
X_15122_ _15417_/A _15120_/Y _15405_/A _15121_/Y VGND VGND VPWR VPWR _15127_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16342__B1 _16055_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15053_ _14981_/A VGND VGND VPWR VPWR _15241_/A sky130_fd_sc_hd__buf_2
X_19930_ _19929_/Y _19925_/X _19613_/X _19925_/X VGND VGND VPWR VPWR _19930_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_182_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_7_127_0_HCLK clkbuf_6_63_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_255_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_12265_ _12172_/Y _12194_/Y VGND VGND VPWR VPWR _12265_/X sky130_fd_sc_hd__or2_4
XFILLER_147_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19574__A _13807_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16893__B2 _24274_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14004_ _13973_/X _13984_/X _13995_/X _14003_/X VGND VGND VPWR VPWR _14004_/X sky130_fd_sc_hd__a211o_4
XANTENNA_clkbuf_3_6_0_HCLK_A clkbuf_3_7_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19861_ _19861_/A VGND VGND VPWR VPWR _19861_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21609__A _22221_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12196_ _25457_/Q _24772_/Q _12194_/Y _12195_/Y VGND VGND VPWR VPWR _12196_/X sky130_fd_sc_hd__o22a_4
XANTENNA__24173__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18812_ _18793_/A _18812_/B _18811_/X VGND VGND VPWR VPWR _24131_/D sky130_fd_sc_hd__and3_4
X_19792_ _19791_/Y _19789_/X _19702_/X _19789_/X VGND VGND VPWR VPWR _23615_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24102__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18743_ _18743_/A VGND VGND VPWR VPWR _24148_/D sky130_fd_sc_hd__inv_2
X_15955_ _15783_/X VGND VGND VPWR VPWR _15955_/X sky130_fd_sc_hd__buf_2
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13772__D _13772_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19595__B1 _19408_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14906_ _25026_/Q VGND VGND VPWR VPWR _15062_/A sky130_fd_sc_hd__inv_2
X_18674_ _24152_/Q VGND VGND VPWR VPWR _18697_/A sky130_fd_sc_hd__inv_2
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15886_ _15879_/X _15880_/X _16236_/A _24797_/Q _15881_/X VGND VGND VPWR VPWR _24797_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_63_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25379__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17625_ _17625_/A _17621_/Y _17625_/C VGND VGND VPWR VPWR _17625_/X sky130_fd_sc_hd__or3_4
X_14837_ _14805_/X _14836_/X _25196_/Q _14830_/X VGND VGND VPWR VPWR _14837_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12966__A _21027_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17556_ _17555_/X VGND VGND VPWR VPWR _17602_/B sky130_fd_sc_hd__buf_2
Xclkbuf_8_65_0_HCLK clkbuf_7_32_0_HCLK/X VGND VGND VPWR VPWR _24263_/CLK sky130_fd_sc_hd__clkbuf_1
X_14768_ _14768_/A VGND VGND VPWR VPWR _14769_/C sky130_fd_sc_hd__inv_2
XANTENNA__13092__C1 _13019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16507_ _16507_/A VGND VGND VPWR VPWR _16507_/Y sky130_fd_sc_hd__inv_2
X_13719_ _13668_/X _13718_/X _13667_/X _13700_/X _11829_/A VGND VGND VPWR VPWR _25282_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_232_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17487_ _17487_/A _17487_/B _17483_/X _17486_/X VGND VGND VPWR VPWR _17487_/X sky130_fd_sc_hd__or4_4
X_14699_ _13731_/X _14699_/B VGND VGND VPWR VPWR _14699_/X sky130_fd_sc_hd__or2_4
X_19226_ _19226_/A VGND VGND VPWR VPWR _19226_/Y sky130_fd_sc_hd__inv_2
X_16438_ _24580_/Q VGND VGND VPWR VPWR _16438_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16581__B1 _16320_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13797__A _13797_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19157_ _19155_/Y _19156_/X _19063_/X _19156_/X VGND VGND VPWR VPWR _19157_/X sky130_fd_sc_hd__a2bb2o_4
X_16369_ _16375_/A VGND VGND VPWR VPWR _16370_/A sky130_fd_sc_hd__buf_2
X_18108_ _17981_/A _18108_/B _18107_/X VGND VGND VPWR VPWR _18108_/X sky130_fd_sc_hd__and3_4
XANTENNA__24943__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19088_ _19088_/A VGND VGND VPWR VPWR _19088_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16333__B1 _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18039_ _18182_/A _18039_/B VGND VGND VPWR VPWR _18039_/X sky130_fd_sc_hd__or2_4
XFILLER_160_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21050_ _21040_/X _21046_/X _21047_/X _21049_/X VGND VGND VPWR VPWR _21051_/C sky130_fd_sc_hd__a211o_4
XANTENNA__21519__A _21519_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22421__A3 _22296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20001_ _21799_/B _19996_/X _19977_/X _19996_/X VGND VGND VPWR VPWR _20001_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21952_ _21937_/A _21952_/B _21952_/C VGND VGND VPWR VPWR _21952_/X sky130_fd_sc_hd__and3_4
X_24740_ _24744_/CLK _16013_/X HRESETn VGND VGND VPWR VPWR _24740_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20903_ _20898_/Y _20894_/Y _20902_/Y VGND VGND VPWR VPWR _20903_/X sky130_fd_sc_hd__and3_4
X_24671_ _24678_/CLK _16204_/X HRESETn VGND VGND VPWR VPWR _23074_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_199_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21883_ _21902_/A _19816_/Y VGND VGND VPWR VPWR _21883_/X sky130_fd_sc_hd__or2_4
XFILLER_215_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12876__A _12759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25049__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11780__A _11780_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23622_ _23806_/CLK _19774_/X VGND VGND VPWR VPWR _19773_/A sky130_fd_sc_hd__dfxtp_4
X_20834_ _20827_/A VGND VGND VPWR VPWR _20834_/X sky130_fd_sc_hd__buf_2
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23553_ _23441_/CLK _23553_/D VGND VGND VPWR VPWR _23553_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21696__A1 _21689_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20765_ _13107_/A _20760_/X _20764_/X VGND VGND VPWR VPWR _20765_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_223_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22504_ _14929_/Y _22452_/X _21582_/X _22503_/X VGND VGND VPWR VPWR _22504_/X sky130_fd_sc_hd__o22a_4
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23484_ _23476_/CLK _23484_/D VGND VGND VPWR VPWR _23484_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__21701__B _23002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20696_ _20716_/A VGND VGND VPWR VPWR _20696_/X sky130_fd_sc_hd__buf_2
XFILLER_195_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22085__A _22365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_195_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25223_ _25100_/CLK _25223_/D HRESETn VGND VGND VPWR VPWR _25223_/Q sky130_fd_sc_hd__dfrtp_4
X_22435_ _22435_/A VGND VGND VPWR VPWR _22437_/A sky130_fd_sc_hd__buf_2
XANTENNA__24684__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25154_ _25158_/CLK _14361_/X HRESETn VGND VGND VPWR VPWR _25154_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22366_ _22383_/A _22366_/B _22365_/X VGND VGND VPWR VPWR _22366_/X sky130_fd_sc_hd__and3_4
XFILLER_108_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24105_ _24159_/CLK _20974_/X HRESETn VGND VGND VPWR VPWR _24105_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24613__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21317_ _21598_/A VGND VGND VPWR VPWR _21317_/X sky130_fd_sc_hd__buf_2
X_25085_ _25098_/CLK _25085_/D HRESETn VGND VGND VPWR VPWR _25085_/Q sky130_fd_sc_hd__dfrtp_4
X_22297_ _22294_/X _22295_/X _22296_/X _24861_/Q _22282_/A VGND VGND VPWR VPWR _22298_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_105_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22948__A1 _12248_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12050_ _12050_/A VGND VGND VPWR VPWR _13800_/B sky130_fd_sc_hd__buf_2
X_24036_ _24035_/CLK _20833_/Y HRESETn VGND VGND VPWR VPWR _24036_/Q sky130_fd_sc_hd__dfrtp_4
X_21248_ _21241_/X _21246_/X _21247_/X VGND VGND VPWR VPWR _21248_/X sky130_fd_sc_hd__o21a_4
XFILLER_104_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12361__B2 _12332_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21179_ _24212_/Q _21179_/B VGND VGND VPWR VPWR _21181_/B sky130_fd_sc_hd__or2_4
XANTENNA__11674__B _13765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19577__B1 _19414_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15740_ _15724_/X _15738_/X _15739_/X _24870_/Q _15736_/X VGND VGND VPWR VPWR _24870_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_133_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12358__A2_N _12356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12952_ _12952_/A _12952_/B _12951_/Y VGND VGND VPWR VPWR _12952_/X sky130_fd_sc_hd__and3_4
X_24938_ _23476_/CLK _15509_/X HRESETn VGND VGND VPWR VPWR _24938_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__25472__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11903_ _11901_/Y _11898_/X _11902_/X _11898_/X VGND VGND VPWR VPWR _11903_/X sky130_fd_sc_hd__a2bb2o_4
X_15671_ _15671_/A _15670_/X VGND VGND VPWR VPWR _15671_/X sky130_fd_sc_hd__or2_4
XFILLER_93_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12883_ _12875_/B VGND VGND VPWR VPWR _12884_/B sky130_fd_sc_hd__inv_2
X_24869_ _25403_/CLK _15742_/X HRESETn VGND VGND VPWR VPWR _24869_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25401__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17410_/A VGND VGND VPWR VPWR _21368_/A sky130_fd_sc_hd__buf_2
XPHY_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14610_/X _14606_/Y _14621_/X _21964_/A _14611_/Y VGND VGND VPWR VPWR _25080_/D
+ sky130_fd_sc_hd__a32o_4
X_11834_ _11832_/A _24234_/Q _11832_/Y _11833_/Y VGND VGND VPWR VPWR _11834_/X sky130_fd_sc_hd__o22a_4
X_18390_ _24109_/Q _18372_/X _24191_/Q _18386_/X VGND VGND VPWR VPWR _24191_/D sky130_fd_sc_hd__o22a_4
XPHY_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17341_/A VGND VGND VPWR VPWR _17351_/A sky130_fd_sc_hd__buf_2
XFILLER_214_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _13826_/A VGND VGND VPWR VPWR _11765_/X sky130_fd_sc_hd__buf_2
X_14553_ _14553_/A _14553_/B VGND VGND VPWR VPWR _14554_/B sky130_fd_sc_hd__or2_4
XFILLER_186_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13503_/Y _13499_/X _13459_/X _13499_/X VGND VGND VPWR VPWR _25307_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17272_ _17272_/A VGND VGND VPWR VPWR _17273_/B sky130_fd_sc_hd__inv_2
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _11694_/Y _11692_/X _11695_/X _11692_/X VGND VGND VPWR VPWR _25542_/D sky130_fd_sc_hd__a2bb2o_4
X_14484_ _20605_/A VGND VGND VPWR VPWR _14484_/X sky130_fd_sc_hd__buf_2
XANTENNA__16563__B1 _16301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19011_ _19011_/A VGND VGND VPWR VPWR _19011_/X sky130_fd_sc_hd__buf_2
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16223_ _16239_/A VGND VGND VPWR VPWR _16223_/X sky130_fd_sc_hd__buf_2
X_13435_ _13334_/A _13435_/B VGND VGND VPWR VPWR _13435_/X sky130_fd_sc_hd__or2_4
XFILLER_139_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22100__A2 _21863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13366_ _13252_/A _23917_/Q VGND VGND VPWR VPWR _13368_/B sky130_fd_sc_hd__or2_4
X_16154_ _16154_/A VGND VGND VPWR VPWR _16154_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24354__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15105_ _25005_/Q _15104_/A _15304_/C _15104_/Y VGND VGND VPWR VPWR _15105_/X sky130_fd_sc_hd__o22a_4
X_12317_ _12315_/A _24849_/Q _12315_/Y _12316_/Y VGND VGND VPWR VPWR _12317_/X sky130_fd_sc_hd__o22a_4
XFILLER_170_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13297_ _13334_/A _18920_/A VGND VGND VPWR VPWR _13297_/X sky130_fd_sc_hd__or2_4
X_16085_ _16084_/X VGND VGND VPWR VPWR _16086_/A sky130_fd_sc_hd__buf_2
XANTENNA__16721__A _16721_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14877__B1 _14876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12248_ _12248_/A VGND VGND VPWR VPWR _12248_/Y sky130_fd_sc_hd__inv_2
X_15036_ _25014_/Q _15023_/Y _15249_/A _16765_/A VGND VGND VPWR VPWR _15042_/A sky130_fd_sc_hd__a2bb2o_4
X_19913_ _19911_/Y _19912_/X _19824_/X _19912_/X VGND VGND VPWR VPWR _19913_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20243__A _20243_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19844_ _23598_/Q VGND VGND VPWR VPWR _21770_/B sky130_fd_sc_hd__inv_2
XANTENNA__16618__B2 _16541_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12179_ _25459_/Q VGND VGND VPWR VPWR _12278_/A sky130_fd_sc_hd__inv_2
XANTENNA__13783__C _13772_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19775_ _23621_/Q VGND VGND VPWR VPWR _21610_/B sky130_fd_sc_hd__inv_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15056__B _15261_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16987_ _16987_/A _16987_/B _16977_/X _16986_/X VGND VGND VPWR VPWR _16987_/X sky130_fd_sc_hd__or4_4
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18726_ _18724_/X _18720_/Y _18726_/C VGND VGND VPWR VPWR _18726_/X sky130_fd_sc_hd__or3_4
X_15938_ _15923_/X _15928_/X HWDATA[25] _23101_/A _15926_/X VGND VGND VPWR VPWR _15938_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21074__A _21056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18657_ _16610_/Y _24130_/Q _16550_/A _18665_/A VGND VGND VPWR VPWR _18662_/B sky130_fd_sc_hd__a2bb2o_4
X_15869_ _12760_/Y _15865_/X _11688_/X _15865_/X VGND VGND VPWR VPWR _15869_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17608_ _17494_/A _17607_/Y VGND VGND VPWR VPWR _17608_/X sky130_fd_sc_hd__or2_4
XFILLER_240_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18588_ _18420_/Y _18592_/B VGND VGND VPWR VPWR _18593_/A sky130_fd_sc_hd__or2_4
XANTENNA__13065__C1 _13019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_10_0_HCLK_A clkbuf_3_5_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21224__D _21223_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17539_ _17535_/X _17536_/X _17539_/C _17539_/D VGND VGND VPWR VPWR _17539_/X sky130_fd_sc_hd__or4_4
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22875__B1 _25386_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20550_ _14435_/Y _20543_/X _20600_/A _20549_/X VGND VGND VPWR VPWR _20550_/X sky130_fd_sc_hd__a211o_4
XFILLER_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21521__B _23002_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_6_9_0_HCLK clkbuf_5_4_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_9_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_220_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19209_ _19209_/A _19094_/B _20387_/C VGND VGND VPWR VPWR _19209_/X sky130_fd_sc_hd__or3_4
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20481_ _20478_/Y _20525_/C _20480_/X VGND VGND VPWR VPWR _20481_/X sky130_fd_sc_hd__a21o_4
X_22220_ _22205_/A _22220_/B _22219_/X VGND VGND VPWR VPWR _22228_/B sky130_fd_sc_hd__or3_4
XANTENNA__22633__A _24760_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24095__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22151_ _22149_/X _22150_/X _22134_/A _24825_/Q _23171_/A VGND VGND VPWR VPWR _22151_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_172_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24024__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21102_ _24612_/Q _22630_/B VGND VGND VPWR VPWR _21102_/X sky130_fd_sc_hd__or2_4
X_22082_ _22077_/X _22081_/X _14666_/X VGND VGND VPWR VPWR _22082_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__21249__A _21622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_110_0_HCLK clkbuf_6_55_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_110_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17446__B _21176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21033_ _21832_/A VGND VGND VPWR VPWR _22525_/A sky130_fd_sc_hd__buf_2
XANTENNA__11775__A _14380_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22984_ _22721_/A VGND VGND VPWR VPWR _22984_/X sky130_fd_sc_hd__buf_2
XFILLER_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25243__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24723_ _24725_/CLK _24723_/D HRESETn VGND VGND VPWR VPWR _24723_/Q sky130_fd_sc_hd__dfrtp_4
X_21935_ _21935_/A _19948_/Y VGND VGND VPWR VPWR _21937_/B sky130_fd_sc_hd__or2_4
XFILLER_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21866_ _23091_/A _21866_/B _21866_/C VGND VGND VPWR VPWR _21867_/D sky130_fd_sc_hd__and3_4
X_24654_ _24654_/CLK _16250_/X HRESETn VGND VGND VPWR VPWR _24654_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_215_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _13125_/C VGND VGND VPWR VPWR _20817_/Y sky130_fd_sc_hd__inv_2
X_23605_ _23494_/CLK _23605_/D VGND VGND VPWR VPWR _23605_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22866__B1 _24734_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21797_ _21793_/X _21796_/X _17725_/X VGND VGND VPWR VPWR _21797_/X sky130_fd_sc_hd__o21a_4
X_24585_ _24591_/CLK _24585_/D HRESETn VGND VGND VPWR VPWR _15121_/A sky130_fd_sc_hd__dfrtp_4
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22527__B _22686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24865__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15710__A HWDATA[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20748_ _13121_/D VGND VGND VPWR VPWR _20748_/Y sky130_fd_sc_hd__inv_2
X_23536_ _23534_/CLK _23536_/D VGND VGND VPWR VPWR _20017_/A sky130_fd_sc_hd__dfxtp_4
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16545__B1 _16373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15899__A2 _15887_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23467_ _23499_/CLK _23467_/D VGND VGND VPWR VPWR _20196_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20679_ _20673_/A _20676_/Y _20677_/Y _20510_/B _20678_/X VGND VGND VPWR VPWR _20679_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _13225_/A VGND VGND VPWR VPWR _13220_/X sky130_fd_sc_hd__buf_2
X_22418_ _22287_/X _22416_/X _22290_/X _22417_/X VGND VGND VPWR VPWR _22419_/B sky130_fd_sc_hd__o22a_4
X_25206_ _24146_/CLK _14197_/X HRESETn VGND VGND VPWR VPWR _20489_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22094__A1 _14940_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23398_ _23398_/CLK _23398_/D VGND VGND VPWR VPWR _20377_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_164_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22543__A _22543_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13151_ _13142_/X _13148_/X _13150_/X VGND VGND VPWR VPWR _13151_/X sky130_fd_sc_hd__o21a_4
XFILLER_128_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12582__B2 _24859_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22349_ _22345_/X _22348_/X _18301_/A VGND VGND VPWR VPWR _22349_/Y sky130_fd_sc_hd__o21ai_4
X_25137_ _25134_/CLK _25137_/D HRESETn VGND VGND VPWR VPWR _25137_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__21841__A1 _21315_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12102_ _12102_/A VGND VGND VPWR VPWR _12102_/X sky130_fd_sc_hd__buf_2
X_13082_ _13073_/A _13073_/B VGND VGND VPWR VPWR _13082_/Y sky130_fd_sc_hd__nand2_4
X_25068_ _24257_/CLK _14732_/X HRESETn VGND VGND VPWR VPWR _14729_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21159__A _21159_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15520__B2 _15519_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23077__C _23076_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12033_ _16366_/A VGND VGND VPWR VPWR _16181_/A sky130_fd_sc_hd__buf_2
X_16910_ _16910_/A _16905_/X _16910_/C _16909_/X VGND VGND VPWR VPWR _16910_/X sky130_fd_sc_hd__or4_4
X_24019_ _24051_/CLK _20762_/X HRESETn VGND VGND VPWR VPWR _13107_/C sky130_fd_sc_hd__dfrtp_4
XANTENNA__11685__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17890_ _17890_/A VGND VGND VPWR VPWR _21997_/A sky130_fd_sc_hd__inv_2
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16841_ _16841_/A VGND VGND VPWR VPWR _16841_/X sky130_fd_sc_hd__buf_2
XFILLER_238_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_15_0_HCLK clkbuf_4_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_6_31_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_19560_ _21816_/B _19555_/X _11920_/X _19555_/X VGND VGND VPWR VPWR _23694_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__12098__B1 _11765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16772_ _24453_/Q VGND VGND VPWR VPWR _16772_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13984_ _13975_/Y _13984_/B VGND VGND VPWR VPWR _13984_/X sky130_fd_sc_hd__and2_4
XFILLER_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21357__B1 SSn_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18511_ _18481_/A _18510_/X VGND VGND VPWR VPWR _18515_/B sky130_fd_sc_hd__or2_4
XFILLER_219_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15723_ _12527_/Y _15717_/X _11688_/X _15717_/X VGND VGND VPWR VPWR _24879_/D sky130_fd_sc_hd__a2bb2o_4
X_12935_ _12830_/A _12932_/X VGND VGND VPWR VPWR _12936_/C sky130_fd_sc_hd__or2_4
X_19491_ _19491_/A VGND VGND VPWR VPWR _21791_/B sky130_fd_sc_hd__inv_2
XFILLER_74_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15036__B1 _15249_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18442_ _24178_/Q VGND VGND VPWR VPWR _18442_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13405__A _13300_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15654_ _16270_/A VGND VGND VPWR VPWR _15773_/B sky130_fd_sc_hd__buf_2
XFILLER_233_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12866_ _12868_/B VGND VGND VPWR VPWR _12872_/B sky130_fd_sc_hd__inv_2
XFILLER_206_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16784__B1 _16783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22718__A _22416_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14605_ _14604_/Y _13625_/A _21964_/A _13623_/X VGND VGND VPWR VPWR _14605_/X sky130_fd_sc_hd__o22a_4
XANTENNA__21622__A _21622_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _13670_/A _24229_/Q _13670_/A _24229_/Q VGND VGND VPWR VPWR _11817_/X sky130_fd_sc_hd__a2bb2o_4
X_18373_ _18372_/X VGND VGND VPWR VPWR _18373_/Y sky130_fd_sc_hd__inv_2
XPHY_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _15583_/Y _15584_/X _11711_/X _15584_/X VGND VGND VPWR VPWR _15585_/X sky130_fd_sc_hd__a2bb2o_4
X_12797_ _12796_/Y _24808_/Q _12796_/Y _24808_/Q VGND VGND VPWR VPWR _12797_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17314_/C _17305_/X _17276_/X _17322_/B VGND VGND VPWR VPWR _17325_/A sky130_fd_sc_hd__a211o_4
XFILLER_30_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14536_ _14536_/A _14536_/B _14532_/X _14535_/X VGND VGND VPWR VPWR _14536_/X sky130_fd_sc_hd__or4_4
XFILLER_159_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _16240_/A VGND VGND VPWR VPWR _11748_/X sky130_fd_sc_hd__buf_2
XFILLER_239_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__24535__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_139_0_HCLK clkbuf_7_69_0_HCLK/X VGND VGND VPWR VPWR _23785_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17255_ _17255_/A _17254_/X VGND VGND VPWR VPWR _17256_/B sky130_fd_sc_hd__or2_4
X_14467_ _14467_/A VGND VGND VPWR VPWR _14467_/Y sky130_fd_sc_hd__inv_2
X_11679_ _11678_/X VGND VGND VPWR VPWR _22136_/B sky130_fd_sc_hd__buf_2
X_16206_ _16205_/Y _16203_/X _11691_/X _16203_/X VGND VGND VPWR VPWR _16206_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13140__A _13421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13418_ _11951_/A _13402_/X _13417_/X _25328_/Q _11950_/A VGND VGND VPWR VPWR _13418_/X
+ sky130_fd_sc_hd__o32a_4
X_17186_ _17185_/Y VGND VGND VPWR VPWR _17346_/A sky130_fd_sc_hd__buf_2
X_14398_ _14408_/A VGND VGND VPWR VPWR _14398_/X sky130_fd_sc_hd__buf_2
X_16137_ _16135_/Y _16136_/X _11748_/X _16136_/X VGND VGND VPWR VPWR _16137_/X sky130_fd_sc_hd__a2bb2o_4
X_13349_ _13445_/A _23630_/Q VGND VGND VPWR VPWR _13351_/B sky130_fd_sc_hd__or2_4
XFILLER_115_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16451__A _15855_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16068_ _16067_/Y _16065_/X _15469_/X _16065_/X VGND VGND VPWR VPWR _24719_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17266__B _17231_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13522__B1 _13521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15019_ _25013_/Q _14986_/Y _15026_/A _15018_/Y VGND VGND VPWR VPWR _15028_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_229_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25394__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19827_ _19827_/A VGND VGND VPWR VPWR _19827_/X sky130_fd_sc_hd__buf_2
XANTENNA__25323__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17282__A _17175_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19758_ _19758_/A VGND VGND VPWR VPWR _19758_/Y sky130_fd_sc_hd__inv_2
X_18709_ _18735_/A VGND VGND VPWR VPWR _18709_/X sky130_fd_sc_hd__buf_2
X_19689_ _13436_/B VGND VGND VPWR VPWR _19689_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15027__B1 _15246_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21720_ _21720_/A _21719_/X VGND VGND VPWR VPWR _21720_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__13315__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16775__B1 _16522_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21651_ _18274_/A _21648_/X _21510_/A _21650_/Y VGND VGND VPWR VPWR _21652_/A sky130_fd_sc_hd__a211o_4
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_35_0_HCLK clkbuf_7_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_70_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20602_ _14391_/Y _20450_/X VGND VGND VPWR VPWR _20602_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15530__A _15530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24370_ _24365_/CLK _17275_/X HRESETn VGND VGND VPWR VPWR _17273_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_33_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9_0_HCLK_A clkbuf_3_4_0_HCLK/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21582_ _21582_/A VGND VGND VPWR VPWR _21582_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_98_0_HCLK clkbuf_7_99_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_98_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_23321_ _17261_/Y _22485_/X _25399_/Q _22444_/X VGND VGND VPWR VPWR _23321_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__24276__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20533_ _20478_/Y _20532_/X _20479_/B VGND VGND VPWR VPWR _20533_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23935__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24205__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23252_ _17273_/A _22423_/A VGND VGND VPWR VPWR _23252_/X sky130_fd_sc_hd__or2_4
X_20464_ _20444_/A _20449_/X _20464_/C VGND VGND VPWR VPWR _20465_/B sky130_fd_sc_hd__and3_4
X_22203_ _22210_/A _22203_/B VGND VGND VPWR VPWR _22204_/C sky130_fd_sc_hd__or2_4
X_23183_ _23160_/X _23163_/X _23167_/Y _23182_/X VGND VGND VPWR VPWR HRDATA[26] sky130_fd_sc_hd__a211o_4
XFILLER_145_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20395_ _20393_/Y _20389_/X _13829_/A _20394_/X VGND VGND VPWR VPWR _23390_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_3_4_0_HCLK clkbuf_3_5_0_HCLK/A VGND VGND VPWR VPWR clkbuf_3_4_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22134_ _22134_/A VGND VGND VPWR VPWR _22135_/C sky130_fd_sc_hd__buf_2
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22065_ _22059_/X _22064_/X _21773_/X VGND VGND VPWR VPWR _22065_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21016_ _21016_/A _24819_/Q VGND VGND VPWR VPWR _21016_/X sky130_fd_sc_hd__and2_4
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21707__A _24615_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25064__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15705__A _16539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16614__A1_N _16613_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22967_ _21439_/X VGND VGND VPWR VPWR _23103_/A sky130_fd_sc_hd__buf_2
XFILLER_83_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12720_ _12718_/Y _12719_/X _12722_/C VGND VGND VPWR VPWR _12720_/X sky130_fd_sc_hd__and3_4
X_24706_ _24681_/CLK _16102_/X HRESETn VGND VGND VPWR VPWR _23112_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__13225__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21918_ _17707_/X VGND VGND VPWR VPWR _21937_/A sky130_fd_sc_hd__buf_2
XFILLER_203_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22898_ _22898_/A _22897_/X VGND VGND VPWR VPWR _22898_/X sky130_fd_sc_hd__or2_4
X_12651_ _12651_/A VGND VGND VPWR VPWR _12651_/Y sky130_fd_sc_hd__inv_2
X_24637_ _24639_/CLK _24637_/D HRESETn VGND VGND VPWR VPWR _24637_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21849_ _14182_/A VGND VGND VPWR VPWR _21849_/X sky130_fd_sc_hd__buf_2
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22303__A2 _22293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _25429_/Q _12570_/Y _12569_/Y _24859_/Q VGND VGND VPWR VPWR _12582_/X sky130_fd_sc_hd__a2bb2o_4
X_15370_ _15352_/A _15370_/B _15370_/C VGND VGND VPWR VPWR _24991_/D sky130_fd_sc_hd__and3_4
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24568_ _24540_/CLK _24568_/D HRESETn VGND VGND VPWR VPWR _24568_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ _25168_/Q _14314_/X _14320_/Y VGND VGND VPWR VPWR _25168_/D sky130_fd_sc_hd__o21a_4
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23519_ _23912_/CLK _23519_/D VGND VGND VPWR VPWR _13299_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_157_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19847__A _19835_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24499_ _24460_/CLK _24499_/D HRESETn VGND VGND VPWR VPWR _24499_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__18751__A _18613_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ _17040_/A VGND VGND VPWR VPWR _17040_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14252_ _14247_/A VGND VGND VPWR VPWR _14252_/X sky130_fd_sc_hd__buf_2
XANTENNA__23264__B1 _22098_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23369__A _21016_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22273__A _21289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13203_ _13433_/A VGND VGND VPWR VPWR _13369_/A sky130_fd_sc_hd__buf_2
X_14183_ _14182_/X VGND VGND VPWR VPWR _14183_/X sky130_fd_sc_hd__buf_2
XANTENNA__23999__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13134_ _13189_/A VGND VGND VPWR VPWR _13225_/A sky130_fd_sc_hd__buf_2
XANTENNA__23016__B1 _16940_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23928__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18991_ _18990_/Y _18986_/X _18965_/X _18986_/X VGND VGND VPWR VPWR _23894_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13504__B1 _13459_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12307__B2 _12306_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13065_ _12985_/B _13059_/X _13062_/B _13019_/X VGND VGND VPWR VPWR _13065_/X sky130_fd_sc_hd__a211o_4
X_17942_ _17942_/A _17940_/X _17942_/C VGND VGND VPWR VPWR _17942_/X sky130_fd_sc_hd__and3_4
XFILLER_79_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12016_ _11975_/Y _12015_/X _25494_/Q _12015_/X VGND VGND VPWR VPWR _25495_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21617__A _14678_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17873_ _16889_/Y _17873_/B VGND VGND VPWR VPWR _17873_/Y sky130_fd_sc_hd__nand2_4
XFILLER_66_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16824_ _24429_/Q VGND VGND VPWR VPWR _16824_/Y sky130_fd_sc_hd__inv_2
X_19612_ _19612_/A VGND VGND VPWR VPWR _21817_/B sky130_fd_sc_hd__inv_2
XFILLER_120_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19543_ _19360_/A VGND VGND VPWR VPWR _19543_/X sky130_fd_sc_hd__buf_2
X_16755_ _16766_/A VGND VGND VPWR VPWR _16755_/X sky130_fd_sc_hd__buf_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13967_ _14007_/A VGND VGND VPWR VPWR _13967_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15706_ _15736_/A VGND VGND VPWR VPWR _15706_/X sky130_fd_sc_hd__buf_2
XFILLER_207_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13135__A _13225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24787__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12918_ _12917_/X VGND VGND VPWR VPWR _25382_/D sky130_fd_sc_hd__inv_2
X_19474_ _23723_/Q VGND VGND VPWR VPWR _21188_/B sky130_fd_sc_hd__inv_2
XFILLER_234_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16686_ _22684_/A _16680_/X _15743_/X _16685_/X VGND VGND VPWR VPWR _24492_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13898_ _13888_/A _13898_/B _13892_/A _13935_/B VGND VGND VPWR VPWR _13917_/B sky130_fd_sc_hd__or4_4
XANTENNA__21750__B1 _21596_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22448__A _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18425_ _18398_/X _18406_/X _18415_/X _18424_/X VGND VGND VPWR VPWR _18425_/X sky130_fd_sc_hd__or4_4
XANTENNA__24716__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15637_ _22111_/A VGND VGND VPWR VPWR _22829_/A sky130_fd_sc_hd__buf_2
X_12849_ _12861_/A _12847_/X _12848_/X VGND VGND VPWR VPWR _25399_/D sky130_fd_sc_hd__and3_4
XANTENNA__22167__B _21849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_5_2_0_HCLK_A clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18356_ _17476_/X _18356_/B VGND VGND VPWR VPWR _18356_/X sky130_fd_sc_hd__or2_4
X_15568_ _15566_/Y _15561_/X _15567_/X _15561_/X VGND VGND VPWR VPWR _15568_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__16509__B1 _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21502__B1 _21501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17307_ _17249_/D _17307_/B VGND VGND VPWR VPWR _17310_/B sky130_fd_sc_hd__or2_4
X_14519_ _21347_/A _14499_/X _25102_/Q _14494_/X VGND VGND VPWR VPWR _14519_/X sky130_fd_sc_hd__o22a_4
XFILLER_230_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18287_ _18283_/X _17728_/X _18279_/X _17706_/X VGND VGND VPWR VPWR _24218_/D sky130_fd_sc_hd__o22a_4
X_15499_ _15489_/A VGND VGND VPWR VPWR _15499_/X sky130_fd_sc_hd__buf_2
XANTENNA__17182__B1 _16339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17238_ _21856_/A VGND VGND VPWR VPWR _17345_/A sky130_fd_sc_hd__inv_2
XFILLER_163_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17169_ _17169_/A _17164_/X _17167_/X _17168_/X VGND VGND VPWR VPWR _17169_/X sky130_fd_sc_hd__or4_4
XFILLER_190_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16181__A _16181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23270__A3 _22849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23007__B1 _22991_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20180_ _20180_/A VGND VGND VPWR VPWR _20180_/X sky130_fd_sc_hd__buf_2
XFILLER_116_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25504__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12742__A2_N _24801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23870_ _25171_/CLK _23870_/D VGND VGND VPWR VPWR _23870_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16996__B1 _16040_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22821_ _22821_/A _22821_/B _22505_/B VGND VGND VPWR VPWR _22821_/X sky130_fd_sc_hd__and3_4
XFILLER_72_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25540_ _24310_/CLK _25540_/D HRESETn VGND VGND VPWR VPWR _11710_/A sky130_fd_sc_hd__dfrtp_4
X_22752_ _21077_/A _22749_/X _22712_/A _22751_/X VGND VGND VPWR VPWR _22752_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_37_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24457__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21703_ _22716_/A _21703_/B VGND VGND VPWR VPWR _21703_/X sky130_fd_sc_hd__and2_4
X_22683_ _22683_/A _22730_/A VGND VGND VPWR VPWR _22683_/X sky130_fd_sc_hd__and2_4
X_25471_ _25471_/CLK _25471_/D HRESETn VGND VGND VPWR VPWR _25471_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12884__A _12796_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21634_ _21771_/A _21634_/B VGND VGND VPWR VPWR _21635_/C sky130_fd_sc_hd__or2_4
X_24422_ _24073_/CLK _16839_/X HRESETn VGND VGND VPWR VPWR _24422_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__22297__A1 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22297__B2 _22282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21565_ _15662_/A VGND VGND VPWR VPWR _21730_/A sky130_fd_sc_hd__buf_2
X_24353_ _24346_/CLK _17340_/Y HRESETn VGND VGND VPWR VPWR _24353_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__18571__A _18400_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20516_ _20516_/A _14271_/X _20510_/B VGND VGND VPWR VPWR _20516_/X sky130_fd_sc_hd__and3_4
X_23304_ _23213_/A _23304_/B _23304_/C VGND VGND VPWR VPWR _23305_/D sky130_fd_sc_hd__and3_4
Xclkbuf_8_122_0_HCLK clkbuf_7_61_0_HCLK/X VGND VGND VPWR VPWR _24907_/CLK sky130_fd_sc_hd__clkbuf_1
X_24284_ _24275_/CLK _17794_/Y HRESETn VGND VGND VPWR VPWR _24284_/Q sky130_fd_sc_hd__dfrtp_4
X_21496_ _21817_/A _21496_/B VGND VGND VPWR VPWR _21496_/X sky130_fd_sc_hd__or2_4
XFILLER_119_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_8_185_0_HCLK clkbuf_7_92_0_HCLK/X VGND VGND VPWR VPWR _25224_/CLK sky130_fd_sc_hd__clkbuf_1
X_23235_ _23235_/A _23235_/B VGND VGND VPWR VPWR _23235_/Y sky130_fd_sc_hd__nor2_4
X_20447_ _20461_/A _20444_/X _20447_/C _20446_/X VGND VGND VPWR VPWR _20447_/X sky130_fd_sc_hd__or4_4
XFILLER_118_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23166_ _23120_/X _23164_/X _23123_/X _23165_/X VGND VGND VPWR VPWR _23167_/B sky130_fd_sc_hd__o22a_4
X_20378_ _20377_/Y _20375_/Y _15762_/X _20375_/Y VGND VGND VPWR VPWR _23398_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15487__B1 HWRITE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22117_ _21569_/X _22115_/X _21575_/X _22116_/X VGND VGND VPWR VPWR _22117_/X sky130_fd_sc_hd__o22a_4
X_23097_ _22761_/X _23095_/X _22691_/X _23096_/X VGND VGND VPWR VPWR _23097_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22048_ _22048_/A _19585_/X VGND VGND VPWR VPWR _22048_/X sky130_fd_sc_hd__and2_4
XANTENNA__21437__A _21232_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20232__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14870_ _14869_/X VGND VGND VPWR VPWR _14870_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13821_ _13820_/Y _13817_/X _11753_/X _13817_/X VGND VGND VPWR VPWR _13821_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23999_ _25226_/CLK _20460_/X HRESETn VGND VGND VPWR VPWR _23999_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16540_ _16792_/A _16540_/B VGND VGND VPWR VPWR _16547_/A sky130_fd_sc_hd__nor2_4
XANTENNA__24880__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13752_ _13743_/X _13748_/Y _19898_/D _14697_/A VGND VGND VPWR VPWR _13752_/X sky130_fd_sc_hd__o22a_4
XFILLER_44_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24198__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12703_ _12686_/A _12697_/B _12703_/C VGND VGND VPWR VPWR _25410_/D sky130_fd_sc_hd__and3_4
X_16471_ _16469_/Y _16470_/X _16382_/X _16470_/X VGND VGND VPWR VPWR _16471_/X sky130_fd_sc_hd__a2bb2o_4
X_13683_ _13683_/A VGND VGND VPWR VPWR _13683_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18210_ _18146_/A _18210_/B VGND VGND VPWR VPWR _18210_/X sky130_fd_sc_hd__or2_4
XANTENNA__24127__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15422_ _15422_/A VGND VGND VPWR VPWR _15422_/Y sky130_fd_sc_hd__inv_2
X_12634_ _12648_/A _12634_/B _12634_/C VGND VGND VPWR VPWR _12634_/X sky130_fd_sc_hd__and3_4
X_19190_ _19190_/A VGND VGND VPWR VPWR _19190_/Y sky130_fd_sc_hd__inv_2
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18141_ _18044_/A _18141_/B _18140_/X VGND VGND VPWR VPWR _18141_/X sky130_fd_sc_hd__or3_4
XANTENNA__12820__A1_N _12828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15353_ _15293_/B _15347_/X _15313_/A _15349_/Y VGND VGND VPWR VPWR _15353_/X sky130_fd_sc_hd__a211o_4
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _12564_/Y _24870_/Q _12564_/Y _24870_/Q VGND VGND VPWR VPWR _12566_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_7_81_0_HCLK clkbuf_7_81_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_81_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ _25175_/Q _14291_/X _25174_/Q _14296_/X VGND VGND VPWR VPWR _14304_/X sky130_fd_sc_hd__o22a_4
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18072_ _18220_/A _18072_/B _18071_/X VGND VGND VPWR VPWR _18072_/X sky130_fd_sc_hd__or3_4
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15284_ _15281_/A VGND VGND VPWR VPWR _15338_/A sky130_fd_sc_hd__buf_2
XFILLER_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _21078_/A _13028_/A VGND VGND VPWR VPWR _12497_/C sky130_fd_sc_hd__or2_4
XFILLER_172_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17023_ _17023_/A VGND VGND VPWR VPWR _17023_/Y sky130_fd_sc_hd__inv_2
X_14235_ _13956_/A _15436_/A _13962_/A VGND VGND VPWR VPWR _14235_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14166_ _25131_/Q VGND VGND VPWR VPWR _14166_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13117_ _13117_/A _13117_/B _20727_/A _20722_/A VGND VGND VPWR VPWR _13117_/X sky130_fd_sc_hd__or4_4
X_14097_ _14097_/A VGND VGND VPWR VPWR _14115_/A sky130_fd_sc_hd__buf_2
X_18974_ _17937_/B VGND VGND VPWR VPWR _18974_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12034__A _16181_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13048_ _13048_/A _13048_/B _13047_/Y VGND VGND VPWR VPWR _13048_/X sky130_fd_sc_hd__and3_4
X_17925_ _13528_/C _17924_/Y _17919_/X VGND VGND VPWR VPWR _24252_/D sky130_fd_sc_hd__o21a_4
XFILLER_67_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23265__C _23264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20223__B1 _18250_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24968__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17856_ _17747_/A _17856_/B VGND VGND VPWR VPWR _17858_/B sky130_fd_sc_hd__or2_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21971__B1 _13772_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16807_ _16806_/Y _16804_/X _15721_/X _16804_/X VGND VGND VPWR VPWR _16807_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17787_ _17787_/A VGND VGND VPWR VPWR _17787_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14999_ _14892_/A _14998_/A _15214_/C _14998_/Y VGND VGND VPWR VPWR _14999_/X sky130_fd_sc_hd__o22a_4
XFILLER_207_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__17560__A _17559_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16738_ _16737_/Y _16735_/X _15721_/X _16735_/X VGND VGND VPWR VPWR _16738_/X sky130_fd_sc_hd__a2bb2o_4
X_19526_ _19526_/A VGND VGND VPWR VPWR _19526_/X sky130_fd_sc_hd__buf_2
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21082__A _22523_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24550__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19457_ _19456_/X VGND VGND VPWR VPWR _19457_/Y sky130_fd_sc_hd__inv_2
X_16669_ _16667_/Y _16668_/X _16395_/X _16668_/X VGND VGND VPWR VPWR _24499_/D sky130_fd_sc_hd__a2bb2o_4
X_18408_ _22927_/A _18407_/A _16214_/Y _18407_/Y VGND VGND VPWR VPWR _18408_/X sky130_fd_sc_hd__o22a_4
X_19388_ _19388_/A VGND VGND VPWR VPWR _19388_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18339_ _18326_/C _18326_/B _18932_/B VGND VGND VPWR VPWR _24207_/D sky130_fd_sc_hd__o21a_4
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21350_ _14166_/Y _22327_/B _23926_/Q _21364_/B VGND VGND VPWR VPWR _21356_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20301_ _21672_/B _20300_/X _19981_/X _20300_/X VGND VGND VPWR VPWR _20301_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21281_ _25057_/Q _21281_/B VGND VGND VPWR VPWR _21281_/Y sky130_fd_sc_hd__nor2_4
XFILLER_135_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14424__A _22327_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23020_ _21421_/A _23018_/Y _22831_/X _23019_/X VGND VGND VPWR VPWR _23021_/A sky130_fd_sc_hd__o22a_4
X_20232_ _20231_/Y _20227_/X _19728_/X _20227_/X VGND VGND VPWR VPWR _20232_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__17458__B2 _13157_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18655__B1 _24525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22641__A _16687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20163_ _20163_/A VGND VGND VPWR VPWR _22085_/B sky130_fd_sc_hd__inv_2
XANTENNA__18657__A1_N _16610_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20094_ _23504_/Q VGND VGND VPWR VPWR _22072_/B sky130_fd_sc_hd__inv_2
X_24971_ _24973_/CLK _24971_/D HRESETn VGND VGND VPWR VPWR _13914_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21545__A1_N _12211_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23175__C _23174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20214__B1 _19708_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11783__A _25522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23922_ _23391_/CLK _23922_/D VGND VGND VPWR VPWR _18909_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_45_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24638__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23853_ _23853_/CLK _23853_/D VGND VGND VPWR VPWR _23853_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22506__A2 _22452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22804_ _16820_/A _21871_/X _22801_/X _22803_/X VGND VGND VPWR VPWR _22804_/X sky130_fd_sc_hd__a211o_4
XFILLER_55_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21704__B _23172_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20996_ _14203_/Y _14185_/X VGND VGND VPWR VPWR _23965_/D sky130_fd_sc_hd__and2_4
X_23784_ _24252_/CLK _23784_/D VGND VGND VPWR VPWR _18032_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_214_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24291__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25523_ _24236_/CLK _25523_/D HRESETn VGND VGND VPWR VPWR _25523_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_225_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22735_ _22735_/A _22735_/B VGND VGND VPWR VPWR _22735_/X sky130_fd_sc_hd__and2_4
XANTENNA__24220__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_240_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25454_ _25453_/CLK _12425_/X HRESETn VGND VGND VPWR VPWR _25454_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_197_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22666_ _17245_/Y _22543_/X VGND VGND VPWR VPWR _22669_/A sky130_fd_sc_hd__or2_4
XFILLER_185_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22816__A _22816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24405_ _24645_/CLK _16954_/X HRESETn VGND VGND VPWR VPWR _21014_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_40_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21617_ _14678_/X _21617_/B VGND VGND VPWR VPWR _21617_/X sky130_fd_sc_hd__or2_4
X_25385_ _25387_/CLK _25385_/D HRESETn VGND VGND VPWR VPWR _25385_/Q sky130_fd_sc_hd__dfrtp_4
X_22597_ _22597_/A _21441_/X VGND VGND VPWR VPWR _22597_/X sky130_fd_sc_hd__or2_4
XFILLER_138_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25497__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12350_ _12349_/Y _24842_/Q _12980_/A _12293_/Y VGND VGND VPWR VPWR _12350_/X sky130_fd_sc_hd__a2bb2o_4
X_24336_ _24340_/CLK _17406_/X HRESETn VGND VGND VPWR VPWR _24336_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_139_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21548_ _21289_/X _21525_/X _21530_/X _21544_/X _21547_/X VGND VGND VPWR VPWR _21548_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_217_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12281_ _12981_/C _24831_/Q _12981_/C _24831_/Q VGND VGND VPWR VPWR _12281_/X sky130_fd_sc_hd__a2bb2o_4
X_21479_ _22261_/A VGND VGND VPWR VPWR _21809_/A sky130_fd_sc_hd__buf_2
X_24267_ _24686_/CLK _17866_/X HRESETn VGND VGND VPWR VPWR _16915_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14020_ _14020_/A VGND VGND VPWR VPWR _14020_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23218_ _23277_/A _23217_/X VGND VGND VPWR VPWR _23218_/X sky130_fd_sc_hd__and2_4
XANTENNA__18646__B1 _16584_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24198_ _24159_/CLK _24198_/D HRESETn VGND VGND VPWR VPWR _18371_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_150_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23149_ _22971_/X _23148_/X _22973_/X _24881_/Q _22974_/X VGND VGND VPWR VPWR _23150_/B
+ sky130_fd_sc_hd__a32o_4
XFILLER_150_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15971_ _12169_/Y _15968_/X _15619_/X _15968_/X VGND VGND VPWR VPWR _24754_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12789__A _22713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17710_ _24217_/Q VGND VGND VPWR VPWR _19455_/A sky130_fd_sc_hd__buf_2
X_14922_ _14922_/A VGND VGND VPWR VPWR _14922_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15165__A _15165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18690_ _24140_/Q VGND VGND VPWR VPWR _18691_/B sky130_fd_sc_hd__inv_2
XFILLER_248_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17641_ _17569_/A _17645_/B _17640_/Y VGND VGND VPWR VPWR _24310_/D sky130_fd_sc_hd__o21a_4
XANTENNA__24379__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14853_ _14809_/A _14809_/B _14809_/A _14809_/B VGND VGND VPWR VPWR _14854_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24308__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ _21958_/B VGND VGND VPWR VPWR _13804_/Y sky130_fd_sc_hd__inv_2
X_17572_ _17659_/A VGND VGND VPWR VPWR _17660_/A sky130_fd_sc_hd__inv_2
XFILLER_205_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14784_ _14784_/A VGND VGND VPWR VPWR _14784_/Y sky130_fd_sc_hd__inv_2
X_11996_ _11995_/X VGND VGND VPWR VPWR _11996_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17811__C _17555_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21705__B1 _24823_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19311_ _19310_/Y _19306_/X _19221_/X _19306_/X VGND VGND VPWR VPWR _19311_/X sky130_fd_sc_hd__a2bb2o_4
X_16523_ _16520_/Y _16521_/X _16522_/X _16521_/X VGND VGND VPWR VPWR _24553_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13735_ _14683_/A VGND VGND VPWR VPWR _13745_/A sky130_fd_sc_hd__inv_2
XFILLER_16_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21333__C _21333_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19242_ _19242_/A VGND VGND VPWR VPWR _19242_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16454_ _16454_/A VGND VGND VPWR VPWR _16454_/X sky130_fd_sc_hd__buf_2
X_13666_ _13681_/B VGND VGND VPWR VPWR _13666_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15405_ _15405_/A _15405_/B VGND VGND VPWR VPWR _15405_/X sky130_fd_sc_hd__or2_4
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12617_ _12681_/A _12617_/B VGND VGND VPWR VPWR _12626_/D sky130_fd_sc_hd__and2_4
X_19173_ _19172_/Y _19170_/X _19057_/X _19170_/X VGND VGND VPWR VPWR _23831_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16385_ _16384_/Y _16381_/X _16295_/X _16381_/X VGND VGND VPWR VPWR _24605_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13597_ _13597_/A VGND VGND VPWR VPWR _18057_/A sky130_fd_sc_hd__buf_2
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16724__A _16724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18124_ _18124_/A _18120_/X _18124_/C VGND VGND VPWR VPWR _18132_/B sky130_fd_sc_hd__or3_4
X_15336_ _15075_/Y _15338_/B _15335_/Y VGND VGND VPWR VPWR _15336_/X sky130_fd_sc_hd__o21a_4
X_12548_ _25406_/Q VGND VGND VPWR VPWR _12692_/A sky130_fd_sc_hd__inv_2
XFILLER_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22681__A1 _21111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23943__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15529__A2_N _15524_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22681__B2 _22680_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18055_ _18126_/A _19148_/A VGND VGND VPWR VPWR _18056_/C sky130_fd_sc_hd__or2_4
X_15267_ _15261_/B VGND VGND VPWR VPWR _15268_/B sky130_fd_sc_hd__inv_2
X_12479_ _12257_/Y _12476_/B VGND VGND VPWR VPWR _12479_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__17258__C _17232_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17006_ _24395_/Q VGND VGND VPWR VPWR _17006_/Y sky130_fd_sc_hd__inv_2
X_14218_ _14213_/A VGND VGND VPWR VPWR _14218_/X sky130_fd_sc_hd__buf_2
XANTENNA__22433__A1 _16339_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21236__A2 _21119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15198_ _25031_/Q _15201_/B VGND VGND VPWR VPWR _15199_/C sky130_fd_sc_hd__or2_4
Xclkbuf_8_25_0_HCLK clkbuf_7_12_0_HCLK/X VGND VGND VPWR VPWR _24302_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_153_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14149_ _14149_/A VGND VGND VPWR VPWR _14149_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_88_0_HCLK clkbuf_7_44_0_HCLK/X VGND VGND VPWR VPWR _24766_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__20995__A1 _20496_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17860__A1 _16895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18957_ _23905_/Q VGND VGND VPWR VPWR _18957_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14674__A1 _14666_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15871__B1 _11695_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17908_ _17908_/A VGND VGND VPWR VPWR _17908_/Y sky130_fd_sc_hd__inv_2
X_18888_ _18888_/A VGND VGND VPWR VPWR _18888_/X sky130_fd_sc_hd__buf_2
XFILLER_94_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24731__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17839_ _17838_/X VGND VGND VPWR VPWR _24272_/D sky130_fd_sc_hd__inv_2
XFILLER_94_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24049__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20850_ _20850_/A VGND VGND VPWR VPWR _24040_/D sky130_fd_sc_hd__inv_2
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19509_ _22027_/B _19503_/X _11911_/X _19508_/X VGND VGND VPWR VPWR _19509_/X sky130_fd_sc_hd__a2bb2o_4
X_20781_ _20781_/A VGND VGND VPWR VPWR _20781_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21172__A1 _16789_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17915__A2 _14764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14419__A _25138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22520_ _22520_/A VGND VGND VPWR VPWR _22521_/B sky130_fd_sc_hd__buf_2
XFILLER_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22451_ _22451_/A VGND VGND VPWR VPWR _23075_/B sky130_fd_sc_hd__buf_2
XFILLER_194_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21402_ _21385_/X _21402_/B VGND VGND VPWR VPWR _21403_/C sky130_fd_sc_hd__or2_4
X_22382_ _22379_/A _20065_/Y VGND VGND VPWR VPWR _22383_/C sky130_fd_sc_hd__or2_4
X_25170_ _25164_/CLK _14313_/X HRESETn VGND VGND VPWR VPWR _25170_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21333_ _23176_/A _21333_/B _21333_/C VGND VGND VPWR VPWR _21419_/A sky130_fd_sc_hd__and3_4
X_24121_ _25211_/CLK _18892_/X HRESETn VGND VGND VPWR VPWR _24121_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__11778__A _11682_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21264_ _14688_/A _21262_/X _21263_/X VGND VGND VPWR VPWR _21264_/X sky130_fd_sc_hd__and3_4
X_24052_ _24501_/CLK _24052_/D HRESETn VGND VGND VPWR VPWR _24052_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22424__B2 _21317_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20215_ _18171_/B VGND VGND VPWR VPWR _20215_/Y sky130_fd_sc_hd__inv_2
X_23003_ _15020_/A _23002_/X _22891_/X VGND VGND VPWR VPWR _23003_/X sky130_fd_sc_hd__o21a_4
X_21195_ _21191_/X _21194_/X _24214_/Q VGND VGND VPWR VPWR _21195_/X sky130_fd_sc_hd__o21a_4
XFILLER_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20146_ _20145_/Y _20143_/X _20099_/X _20143_/X VGND VGND VPWR VPWR _23487_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24819__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22188__B1 _22176_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20077_ _20076_/Y _20072_/X _19820_/X _20072_/X VGND VGND VPWR VPWR _23510_/D sky130_fd_sc_hd__a2bb2o_4
X_24954_ _24958_/CLK _15470_/X HRESETn VGND VGND VPWR VPWR _15468_/A sky130_fd_sc_hd__dfstp_4
XFILLER_100_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12402__A _12240_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24472__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23905_ _23875_/CLK _18958_/X VGND VGND VPWR VPWR _23905_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_85_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24885_ _24834_/CLK _15711_/X HRESETn VGND VGND VPWR VPWR _24885_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15614__B1 _11757_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24401__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11850_ _25514_/Q _11856_/B VGND VGND VPWR VPWR _11850_/Y sky130_fd_sc_hd__nand2_4
X_23836_ _23844_/CLK _23836_/D VGND VGND VPWR VPWR _19158_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_45_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _14392_/A VGND VGND VPWR VPWR _11781_/X sky130_fd_sc_hd__buf_2
X_23767_ _23767_/CLK _23767_/D VGND VGND VPWR VPWR _19350_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21163__A1 _21343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20979_ _23372_/Q VGND VGND VPWR VPWR _20979_/Y sky130_fd_sc_hd__inv_2
XPHY_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _13520_/A VGND VGND VPWR VPWR _13520_/Y sky130_fd_sc_hd__inv_2
X_25506_ _23437_/CLK _11916_/X HRESETn VGND VGND VPWR VPWR _19977_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22718_ _22416_/B VGND VGND VPWR VPWR _22718_/X sky130_fd_sc_hd__buf_2
XFILLER_14_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23698_ _23406_/CLK _19551_/X VGND VGND VPWR VPWR _19547_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_202_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13451_ _13186_/A _13450_/X _25326_/Q _13184_/A VGND VGND VPWR VPWR _25326_/D sky130_fd_sc_hd__o22a_4
X_25437_ _25450_/CLK _12485_/Y HRESETn VGND VGND VPWR VPWR _25437_/Q sky130_fd_sc_hd__dfrtp_4
X_22649_ _22648_/X VGND VGND VPWR VPWR _22649_/Y sky130_fd_sc_hd__inv_2
X_12402_ _12240_/Y _12402_/B _12370_/X VGND VGND VPWR VPWR _12402_/X sky130_fd_sc_hd__or3_4
X_16170_ _14764_/X _16170_/B VGND VGND VPWR VPWR _16170_/X sky130_fd_sc_hd__and2_4
XANTENNA__22663__A1 _16539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13382_ _13350_/A _13382_/B VGND VGND VPWR VPWR _13382_/X sky130_fd_sc_hd__or2_4
X_25368_ _25373_/CLK _25368_/D HRESETn VGND VGND VPWR VPWR _21027_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_127_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22663__B2 _21833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25130__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15121_ _15121_/A VGND VGND VPWR VPWR _15121_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11688__A HWDATA[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12333_ _24825_/Q VGND VGND VPWR VPWR _12333_/Y sky130_fd_sc_hd__inv_2
X_24319_ _23411_/CLK _24319_/D HRESETn VGND VGND VPWR VPWR _17561_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__25193__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25299_ _24907_/CLK _25299_/D HRESETn VGND VGND VPWR VPWR _25299_/Q sky130_fd_sc_hd__dfrtp_4
X_15052_ _15051_/X VGND VGND VPWR VPWR _15052_/Y sky130_fd_sc_hd__inv_2
X_12264_ _12264_/A VGND VGND VPWR VPWR _12264_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19574__B _13807_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22281__A _24618_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_241_0_HCLK clkbuf_8_241_0_HCLK/A VGND VGND VPWR VPWR _24574_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_147_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14003_ _13999_/X _14536_/A _13999_/X _14536_/A VGND VGND VPWR VPWR _14003_/X sky130_fd_sc_hd__a2bb2o_4
X_12195_ _24772_/Q VGND VGND VPWR VPWR _12195_/Y sky130_fd_sc_hd__inv_2
X_19860_ _19859_/Y _19857_/X _19603_/X _19857_/X VGND VGND VPWR VPWR _19860_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18811_ _24131_/Q _18811_/B VGND VGND VPWR VPWR _18811_/X sky130_fd_sc_hd__or2_4
XFILLER_96_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19791_ _19791_/A VGND VGND VPWR VPWR _19791_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15954_ _12216_/Y _15949_/X _15953_/X _15949_/X VGND VGND VPWR VPWR _24765_/D sky130_fd_sc_hd__a2bb2o_4
X_18742_ _18735_/A _18738_/Y _18741_/X VGND VGND VPWR VPWR _18743_/A sky130_fd_sc_hd__or3_4
XANTENNA__12312__A _24827_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14905_ _14894_/X _14897_/X _14901_/X _14905_/D VGND VGND VPWR VPWR _14905_/X sky130_fd_sc_hd__or4_4
XFILLER_237_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18673_ _24156_/Q VGND VGND VPWR VPWR _18700_/C sky130_fd_sc_hd__inv_2
XFILLER_236_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21625__A _22379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15885_ _15879_/X _15880_/X _16233_/A _24798_/Q _15881_/X VGND VGND VPWR VPWR _15885_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24142__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15623__A _14407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14836_ _25051_/Q _14796_/X _25051_/Q _14796_/X VGND VGND VPWR VPWR _14836_/X sky130_fd_sc_hd__a2bb2o_4
X_17624_ _17583_/X _17602_/X _17545_/Y VGND VGND VPWR VPWR _17625_/C sky130_fd_sc_hd__o21a_4
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12966__B _12650_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17555_ _17555_/A _17555_/B VGND VGND VPWR VPWR _17555_/X sky130_fd_sc_hd__or2_4
X_14767_ _14758_/B _14763_/Y _14764_/X _14766_/X VGND VGND VPWR VPWR _14768_/A sky130_fd_sc_hd__or4_4
X_11979_ _11979_/A _11990_/A VGND VGND VPWR VPWR _11979_/X sky130_fd_sc_hd__and2_4
XFILLER_17_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18934__A _18947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16506_ _16505_/Y _16501_/X _16236_/X _16501_/X VGND VGND VPWR VPWR _16506_/X sky130_fd_sc_hd__a2bb2o_4
X_13718_ _11829_/A _11836_/A VGND VGND VPWR VPWR _13718_/X sky130_fd_sc_hd__or2_4
X_17486_ _13162_/X _17485_/A _13150_/X _17485_/Y VGND VGND VPWR VPWR _17486_/X sky130_fd_sc_hd__o22a_4
X_14698_ _14664_/X VGND VGND VPWR VPWR _14699_/B sky130_fd_sc_hd__inv_2
XANTENNA__16030__B1 _15953_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25348__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16437_ _15120_/Y _16370_/A _16358_/X _16370_/A VGND VGND VPWR VPWR _24581_/D sky130_fd_sc_hd__a2bb2o_4
X_19225_ _19223_/Y _19224_/X _19200_/X _19224_/X VGND VGND VPWR VPWR _23813_/D sky130_fd_sc_hd__a2bb2o_4
X_13649_ _24047_/Q _13648_/X VGND VGND VPWR VPWR _13649_/X sky130_fd_sc_hd__or2_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19156_ _19149_/A VGND VGND VPWR VPWR _19156_/X sky130_fd_sc_hd__buf_2
XFILLER_192_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16368_ _16368_/A _16792_/B VGND VGND VPWR VPWR _16375_/A sky130_fd_sc_hd__nor2_4
XANTENNA__18858__B1 _24571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18107_ _17979_/X _18107_/B VGND VGND VPWR VPWR _18107_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_51_0_HCLK clkbuf_6_51_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_51_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15319_ _15338_/A _15317_/X _15318_/X VGND VGND VPWR VPWR _25005_/D sky130_fd_sc_hd__and3_4
XFILLER_157_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19087_ _21615_/B _19086_/X _16882_/X _19086_/X VGND VGND VPWR VPWR _19087_/X sky130_fd_sc_hd__a2bb2o_4
X_16299_ _16297_/Y _16292_/X _15939_/X _16298_/X VGND VGND VPWR VPWR _16299_/X sky130_fd_sc_hd__a2bb2o_4
X_18038_ _17984_/X _18036_/X _18038_/C VGND VGND VPWR VPWR _18038_/X sky130_fd_sc_hd__and3_4
XFILLER_105_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22191__A _22191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22957__A2 _22948_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24983__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20000_ _23542_/Q VGND VGND VPWR VPWR _21799_/B sky130_fd_sc_hd__inv_2
XANTENNA__16097__B1 _16004_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24912__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19989_ _18285_/A _18285_/B _18280_/A _18289_/X VGND VGND VPWR VPWR _19989_/X sky130_fd_sc_hd__or4_4
XFILLER_143_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21917__B1 _21284_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21951_ _21936_/A _21951_/B VGND VGND VPWR VPWR _21952_/C sky130_fd_sc_hd__or2_4
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20902_ _24052_/Q VGND VGND VPWR VPWR _20902_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15533__A _15530_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19005__A HWDATA[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24670_ _24678_/CLK _16206_/X HRESETn VGND VGND VPWR VPWR _23064_/A sky130_fd_sc_hd__dfrtp_4
X_21882_ _21882_/A _21881_/X VGND VGND VPWR VPWR _21882_/X sky130_fd_sc_hd__and2_4
XFILLER_199_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _23859_/CLK _23621_/D VGND VGND VPWR VPWR _23621_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833_ _20833_/A VGND VGND VPWR VPWR _20833_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16967__A1_N _16073_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23552_ _23534_/CLK _23552_/D VGND VGND VPWR VPWR _19969_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_211_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20764_ _20759_/Y _20755_/Y _20764_/C VGND VGND VPWR VPWR _20764_/X sky130_fd_sc_hd__and3_4
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16021__B1 _16020_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19894__A1_N _19893_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25089__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22503_ _15008_/Y _22505_/B VGND VGND VPWR VPWR _22503_/X sky130_fd_sc_hd__and2_4
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20695_ _20695_/A VGND VGND VPWR VPWR _20695_/Y sky130_fd_sc_hd__inv_2
X_23483_ _23499_/CLK _23483_/D VGND VGND VPWR VPWR _23483_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_210_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25018__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25222_ _25113_/CLK _14127_/X HRESETn VGND VGND VPWR VPWR _14092_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_210_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22434_ _22430_/X _22433_/X VGND VGND VPWR VPWR _22443_/B sky130_fd_sc_hd__nor2_4
XANTENNA__18849__B1 _16520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16083__B _22505_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25153_ _23926_/CLK _25153_/D HRESETn VGND VGND VPWR VPWR _20469_/A sky130_fd_sc_hd__dfrtp_4
X_22365_ _22365_/A _22365_/B VGND VGND VPWR VPWR _22365_/X sky130_fd_sc_hd__or2_4
XFILLER_164_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24104_ _24159_/CLK _20973_/X HRESETn VGND VGND VPWR VPWR _12115_/A sky130_fd_sc_hd__dfrtp_4
X_21316_ _22429_/A VGND VGND VPWR VPWR _22543_/A sky130_fd_sc_hd__buf_2
X_22296_ _21311_/X VGND VGND VPWR VPWR _22296_/X sky130_fd_sc_hd__buf_2
X_25084_ _25098_/CLK _14600_/X HRESETn VGND VGND VPWR VPWR _25084_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21247_ _14706_/A VGND VGND VPWR VPWR _21247_/X sky130_fd_sc_hd__buf_2
X_24035_ _24035_/CLK _20830_/Y HRESETn VGND VGND VPWR VPWR _24035_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24653__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21178_ _21178_/A VGND VGND VPWR VPWR _21178_/X sky130_fd_sc_hd__buf_2
XFILLER_77_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_71_0_HCLK clkbuf_8_70_0_HCLK/A VGND VGND VPWR VPWR _25450_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA__15835__B1 _24820_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20129_ _21636_/B _20128_/X _20106_/X _20128_/X VGND VGND VPWR VPWR _20129_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11674__C _15640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21908__B1 _22205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21445__A _21034_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12951_ _12948_/A _12948_/B VGND VGND VPWR VPWR _12951_/Y sky130_fd_sc_hd__nand2_4
X_24937_ _23476_/CLK _15513_/X HRESETn VGND VGND VPWR VPWR _24937_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16539__A _16539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11902_ _19600_/A VGND VGND VPWR VPWR _11902_/X sky130_fd_sc_hd__buf_2
XFILLER_234_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15670_ _16368_/A VGND VGND VPWR VPWR _15670_/X sky130_fd_sc_hd__buf_2
X_12882_ _12881_/X VGND VGND VPWR VPWR _25392_/D sky130_fd_sc_hd__inv_2
X_24868_ _24866_/CLK _24868_/D HRESETn VGND VGND VPWR VPWR _24868_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16260__B1 _15469_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14606_/A _14605_/X VGND VGND VPWR VPWR _14621_/X sky130_fd_sc_hd__or2_4
XPHY_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _24234_/Q VGND VGND VPWR VPWR _11833_/Y sky130_fd_sc_hd__inv_2
X_23819_ _23827_/CLK _23819_/D VGND VGND VPWR VPWR _23819_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _24800_/CLK _15884_/X HRESETn VGND VGND VPWR VPWR _22714_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__21136__B2 _21368_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17340_/A VGND VGND VPWR VPWR _17340_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14552_/A _14551_/X VGND VGND VPWR VPWR _14553_/B sky130_fd_sc_hd__or2_4
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ HWDATA[6] VGND VGND VPWR VPWR _13826_/A sky130_fd_sc_hd__buf_2
XPHY_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13503_/A VGND VGND VPWR VPWR _13503_/Y sky130_fd_sc_hd__inv_2
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _17231_/X _17271_/B VGND VGND VPWR VPWR _17272_/A sky130_fd_sc_hd__or2_4
XPHY_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _13965_/X VGND VGND VPWR VPWR _14530_/A sky130_fd_sc_hd__buf_2
XFILLER_158_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ HWDATA[22] VGND VGND VPWR VPWR _11695_/X sky130_fd_sc_hd__buf_2
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19010_ _18045_/B VGND VGND VPWR VPWR _19010_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16222_ _16183_/Y VGND VGND VPWR VPWR _16239_/A sky130_fd_sc_hd__buf_2
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13434_ _13434_/A _13434_/B _13434_/C VGND VGND VPWR VPWR _13434_/X sky130_fd_sc_hd__and3_4
XANTENNA__22636__A1 _21305_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16153_ _16152_/Y _16150_/X _16062_/X _16150_/X VGND VGND VPWR VPWR _24686_/D sky130_fd_sc_hd__a2bb2o_4
X_13365_ _13365_/A _13365_/B _13365_/C VGND VGND VPWR VPWR _13365_/X sky130_fd_sc_hd__and3_4
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17512__B1 _11687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15104_ _15104_/A VGND VGND VPWR VPWR _15104_/Y sky130_fd_sc_hd__inv_2
X_12316_ _24849_/Q VGND VGND VPWR VPWR _12316_/Y sky130_fd_sc_hd__inv_2
X_16084_ _16084_/A VGND VGND VPWR VPWR _16084_/X sky130_fd_sc_hd__buf_2
X_13296_ _13365_/A _13294_/X _13296_/C VGND VGND VPWR VPWR _13296_/X sky130_fd_sc_hd__and3_4
XFILLER_114_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16721__B _16721_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15035_ _15029_/X _15035_/B _15035_/C _15034_/X VGND VGND VPWR VPWR _15035_/X sky130_fd_sc_hd__or4_4
X_19912_ _19900_/A VGND VGND VPWR VPWR _19912_/X sky130_fd_sc_hd__buf_2
X_12247_ _12247_/A VGND VGND VPWR VPWR _12247_/Y sky130_fd_sc_hd__inv_2
XANTENNA__23061__B2 _21227_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24394__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19843_ _19842_/Y _19840_/X _19817_/X _19840_/X VGND VGND VPWR VPWR _19843_/X sky130_fd_sc_hd__a2bb2o_4
X_12178_ _22558_/A VGND VGND VPWR VPWR _12178_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__13783__D _13783_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15826__B1 _15619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24323__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19774_ _21755_/B _19769_/X _16878_/X _19769_/X VGND VGND VPWR VPWR _19774_/X sky130_fd_sc_hd__a2bb2o_4
X_16986_ _16979_/X _16981_/X _16983_/X _16986_/D VGND VGND VPWR VPWR _16986_/X sky130_fd_sc_hd__or4_4
XFILLER_96_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18725_ _18696_/X _18705_/X _18697_/A VGND VGND VPWR VPWR _18726_/C sky130_fd_sc_hd__o21a_4
X_15937_ _15923_/X _15928_/X _15719_/X _23144_/A _15926_/X VGND VGND VPWR VPWR _24774_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_237_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15868_ _15843_/X _15850_/X _15721_/X _24810_/Q _15857_/X VGND VGND VPWR VPWR _15868_/X
+ sky130_fd_sc_hd__a32o_4
X_18656_ _24154_/Q VGND VGND VPWR VPWR _18665_/A sky130_fd_sc_hd__inv_2
XFILLER_25_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24088__D _20962_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25529__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14819_ _14818_/X VGND VGND VPWR VPWR _14838_/A sky130_fd_sc_hd__buf_2
X_17607_ _17597_/B VGND VGND VPWR VPWR _17607_/Y sky130_fd_sc_hd__inv_2
X_15799_ _15777_/X _15789_/X _15721_/X _24845_/Q _15787_/X VGND VGND VPWR VPWR _15799_/X
+ sky130_fd_sc_hd__a32o_4
X_18587_ _18561_/C _18587_/B VGND VGND VPWR VPWR _18592_/B sky130_fd_sc_hd__or2_4
XFILLER_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17538_ _11728_/Y _24306_/Q _11728_/Y _24306_/Q VGND VGND VPWR VPWR _17539_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__25182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17469_ _17487_/B VGND VGND VPWR VPWR _17469_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__25111__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19208_ _20220_/A _19208_/B _18910_/B VGND VGND VPWR VPWR _20387_/C sky130_fd_sc_hd__or3_4
XFILLER_177_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20480_ _14266_/Y _20502_/B _20525_/B VGND VGND VPWR VPWR _20480_/X sky130_fd_sc_hd__and3_4
XFILLER_165_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22914__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19139_ _19137_/Y _19133_/X _19138_/X _19133_/A VGND VGND VPWR VPWR _19139_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22150_ _22150_/A _21101_/A VGND VGND VPWR VPWR _22150_/X sky130_fd_sc_hd__or2_4
XANTENNA__17005__A1_N _16006_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21850__A2 _21849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21101_ _21101_/A VGND VGND VPWR VPWR _22630_/B sky130_fd_sc_hd__buf_2
XFILLER_133_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22081_ _22383_/A _22079_/X _22081_/C VGND VGND VPWR VPWR _22081_/X sky130_fd_sc_hd__and3_4
X_21032_ _21024_/X VGND VGND VPWR VPWR _21832_/A sky130_fd_sc_hd__inv_2
XANTENNA__15817__B1 _24832_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_7_58_0_HCLK clkbuf_7_59_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_58_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24064__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_219_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17743__A _24284_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15832__A3 _15764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22983_ _23160_/A _22970_/X _22983_/C _22982_/X VGND VGND VPWR VPWR _22983_/X sky130_fd_sc_hd__or4_4
XANTENNA__11791__A HWDATA[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24722_ _24266_/CLK _24722_/D HRESETn VGND VGND VPWR VPWR _24722_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_216_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21934_ _21924_/A VGND VGND VPWR VPWR _21935_/A sky130_fd_sc_hd__buf_2
XFILLER_103_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24653_ _24654_/CLK _16253_/X HRESETn VGND VGND VPWR VPWR _22163_/A sky130_fd_sc_hd__dfrtp_4
X_21865_ _24418_/Q _21863_/X _21730_/A _21864_/X VGND VGND VPWR VPWR _21866_/C sky130_fd_sc_hd__a211o_4
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23604_ _23499_/CLK _23604_/D VGND VGND VPWR VPWR _19826_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ _20690_/X _20815_/X _15556_/A _20735_/X VGND VGND VPWR VPWR _20816_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24584_ _24591_/CLK _16431_/X HRESETn VGND VGND VPWR VPWR _24584_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21796_ _21484_/X _21796_/B _21795_/X VGND VGND VPWR VPWR _21796_/X sky130_fd_sc_hd__and3_4
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23535_ _23678_/CLK _20021_/X VGND VGND VPWR VPWR _20020_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20747_ _20731_/X _20746_/X _15600_/A _20736_/X VGND VGND VPWR VPWR _20747_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23466_ _23754_/CLK _20202_/X VGND VGND VPWR VPWR _17952_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_149_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15899__A3 _15764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20678_ _20678_/A _14271_/X VGND VGND VPWR VPWR _20678_/X sky130_fd_sc_hd__or2_4
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22824__A _21289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25205_ _24958_/CLK _25205_/D HRESETn VGND VGND VPWR VPWR _25205_/Q sky130_fd_sc_hd__dfrtp_4
X_22417_ _15615_/Y _22417_/B VGND VGND VPWR VPWR _22417_/X sky130_fd_sc_hd__and2_4
XFILLER_136_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12031__A1 _24099_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22094__A2 _22417_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23397_ _23398_/CLK _20379_/X VGND VGND VPWR VPWR _23397_/Q sky130_fd_sc_hd__dfxtp_4
X_13150_ _13433_/A VGND VGND VPWR VPWR _13150_/X sky130_fd_sc_hd__buf_2
X_25136_ _23958_/CLK _25136_/D HRESETn VGND VGND VPWR VPWR _14428_/A sky130_fd_sc_hd__dfstp_4
XANTENNA__24834__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22348_ _21937_/A _22348_/B _22348_/C VGND VGND VPWR VPWR _22348_/X sky130_fd_sc_hd__and3_4
XFILLER_152_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15470__A1_N _15468_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12101_ _25473_/Q VGND VGND VPWR VPWR _12101_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18855__A2_N _24138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13081_ _13085_/A _13074_/X _13081_/C VGND VGND VPWR VPWR _13081_/X sky130_fd_sc_hd__and3_4
X_25067_ _24257_/CLK _25067_/D HRESETn VGND VGND VPWR VPWR _14720_/A sky130_fd_sc_hd__dfrtp_4
X_22279_ _22279_/A VGND VGND VPWR VPWR _22279_/X sky130_fd_sc_hd__buf_2
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12032_ _23350_/A VGND VGND VPWR VPWR _12032_/Y sky130_fd_sc_hd__inv_2
X_24018_ _24051_/CLK _24018_/D HRESETn VGND VGND VPWR VPWR _13121_/C sky130_fd_sc_hd__dfrtp_4
XFILLER_105_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15808__B1 _11718_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16840_ _14917_/Y _16837_/X _16518_/X _16837_/X VGND VGND VPWR VPWR _16840_/X sky130_fd_sc_hd__a2bb2o_4
X_16771_ _15003_/Y _16769_/X _16601_/X _16769_/X VGND VGND VPWR VPWR _16771_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_93_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13983_ _13982_/X VGND VGND VPWR VPWR _13984_/B sky130_fd_sc_hd__inv_2
XANTENNA__21357__A1 SSn_S3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15722_ _15540_/X _15709_/X _15721_/X _24880_/Q _15707_/X VGND VGND VPWR VPWR _24880_/D
+ sky130_fd_sc_hd__a32o_4
X_18510_ _18560_/A _18479_/X _18510_/C _18510_/D VGND VGND VPWR VPWR _18510_/X sky130_fd_sc_hd__or4_4
X_12934_ _12934_/A _12934_/B VGND VGND VPWR VPWR _12936_/B sky130_fd_sc_hd__or2_4
XFILLER_218_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19490_ _21919_/B _19487_/X _11915_/X _19487_/X VGND VGND VPWR VPWR _23719_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15036__B2 _16765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15653_ _21089_/B VGND VGND VPWR VPWR _16270_/A sky130_fd_sc_hd__buf_2
X_18441_ _16256_/Y _24162_/Q _23238_/A _18440_/Y VGND VGND VPWR VPWR _18446_/B sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21903__A _22225_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12865_ _12617_/B _12842_/X VGND VGND VPWR VPWR _12868_/B sky130_fd_sc_hd__or2_4
XPHY_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _21964_/A VGND VGND VPWR VPWR _14604_/Y sky130_fd_sc_hd__inv_2
XPHY_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11816_/A VGND VGND VPWR VPWR _13670_/A sky130_fd_sc_hd__inv_2
X_18372_ _18372_/A _18372_/B _12148_/C _18372_/D VGND VGND VPWR VPWR _18372_/X sky130_fd_sc_hd__or4_4
XFILLER_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15901__A _18951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15576_/A VGND VGND VPWR VPWR _15584_/X sky130_fd_sc_hd__buf_2
XPHY_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12796_/A VGND VGND VPWR VPWR _12796_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17338_/A _17319_/B _17323_/C VGND VGND VPWR VPWR _24358_/D sky130_fd_sc_hd__and3_4
XFILLER_159_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__20868__B1 _20855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _23959_/Q _14535_/B VGND VGND VPWR VPWR _14535_/X sky130_fd_sc_hd__and2_4
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ HWDATA[11] VGND VGND VPWR VPWR _16240_/A sky130_fd_sc_hd__buf_2
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13421__A _13421_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17254_ _17234_/Y _17219_/Y _17236_/X _17253_/X VGND VGND VPWR VPWR _17254_/X sky130_fd_sc_hd__or4_4
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ _14465_/Y _14463_/X _14403_/X _14463_/X VGND VGND VPWR VPWR _25120_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _21519_/A VGND VGND VPWR VPWR _11678_/X sky130_fd_sc_hd__buf_2
XFILLER_128_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16205_ _23064_/A VGND VGND VPWR VPWR _16205_/Y sky130_fd_sc_hd__inv_2
X_13417_ _13385_/A _13409_/X _13416_/X VGND VGND VPWR VPWR _13417_/X sky130_fd_sc_hd__and3_4
X_17185_ _24348_/Q VGND VGND VPWR VPWR _17185_/Y sky130_fd_sc_hd__inv_2
X_14397_ _11676_/A _14442_/B VGND VGND VPWR VPWR _14408_/A sky130_fd_sc_hd__nor2_4
XANTENNA__16732__A _24474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16136_ _16124_/A VGND VGND VPWR VPWR _16136_/X sky130_fd_sc_hd__buf_2
XANTENNA__24575__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13348_ _13231_/X _13346_/X _13347_/X VGND VGND VPWR VPWR _13348_/X sky130_fd_sc_hd__and3_4
XFILLER_182_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__24504__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16067_ _24719_/Q VGND VGND VPWR VPWR _16067_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13279_ _13169_/A _13277_/X _13278_/X VGND VGND VPWR VPWR _13280_/C sky130_fd_sc_hd__and3_4
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15018_ _15018_/A VGND VGND VPWR VPWR _15018_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19826_ _19826_/A VGND VGND VPWR VPWR _21384_/B sky130_fd_sc_hd__inv_2
XFILLER_96_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21085__A _22451_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19757_ _19756_/Y _19754_/X _19711_/X _19754_/X VGND VGND VPWR VPWR _19757_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16969_ _24392_/Q VGND VGND VPWR VPWR _16969_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24919__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16179__A _16179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22545__B1 _22544_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18708_ _18705_/B VGND VGND VPWR VPWR _18735_/A sky130_fd_sc_hd__inv_2
X_19688_ _19687_/Y _19685_/X _19543_/X _19685_/X VGND VGND VPWR VPWR _23652_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16224__B1 _11726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15027__B2 _15018_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25363__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18639_ _24143_/Q VGND VGND VPWR VPWR _18755_/B sky130_fd_sc_hd__inv_2
XFILLER_213_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15811__A _15811_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21650_ _13726_/A _21649_/X VGND VGND VPWR VPWR _21650_/Y sky130_fd_sc_hd__nor2_4
XFILLER_178_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20601_ _20601_/A _20450_/X VGND VGND VPWR VPWR _20603_/B sky130_fd_sc_hd__or2_4
XANTENNA__20859__B1 _20855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21581_ _11678_/X VGND VGND VPWR VPWR _21581_/X sky130_fd_sc_hd__buf_2
XFILLER_221_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23320_ _23320_/A _21525_/A VGND VGND VPWR VPWR _23320_/X sky130_fd_sc_hd__and2_4
XFILLER_138_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14538__B1 sda_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20532_ _15451_/A _24072_/Q _20515_/B VGND VGND VPWR VPWR _20532_/X sky130_fd_sc_hd__and3_4
XFILLER_229_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20463_ _20454_/X _20463_/B VGND VGND VPWR VPWR _20523_/B sky130_fd_sc_hd__and2_4
X_23251_ _23251_/A _23251_/B _23250_/X VGND VGND VPWR VPWR _23251_/X sky130_fd_sc_hd__and3_4
XFILLER_229_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22202_ _22202_/A VGND VGND VPWR VPWR _22210_/A sky130_fd_sc_hd__buf_2
XFILLER_146_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_21_0_HCLK clkbuf_5_21_0_HCLK/A VGND VGND VPWR VPWR clkbuf_6_43_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20394_ _20389_/A VGND VGND VPWR VPWR _20394_/X sky130_fd_sc_hd__buf_2
X_23182_ _23182_/A _23169_/Y _23175_/X _23182_/D VGND VGND VPWR VPWR _23182_/X sky130_fd_sc_hd__or4_4
XANTENNA__20164__A _20158_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24245__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22133_ _21297_/Y VGND VGND VPWR VPWR _22134_/A sky130_fd_sc_hd__buf_2
XANTENNA__19229__B1 _19138_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22064_ _22373_/A _22061_/X _22063_/X VGND VGND VPWR VPWR _22064_/X sky130_fd_sc_hd__and3_4
XFILLER_248_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21015_ _21015_/A _21015_/B VGND VGND VPWR VPWR _23368_/A sky130_fd_sc_hd__and2_4
XANTENNA__21707__B _22130_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__18288__B _17704_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19401__B1 _19377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_145_0_HCLK clkbuf_7_72_0_HCLK/X VGND VGND VPWR VPWR _25325_/CLK sky130_fd_sc_hd__clkbuf_1
X_22966_ _21099_/X VGND VGND VPWR VPWR _23160_/A sky130_fd_sc_hd__buf_2
XFILLER_216_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24705_ _24704_/CLK _24705_/D HRESETn VGND VGND VPWR VPWR _24705_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21917_ _21901_/X _21916_/X _21284_/X VGND VGND VPWR VPWR _21917_/X sky130_fd_sc_hd__a21o_4
X_22897_ _21087_/A VGND VGND VPWR VPWR _22897_/X sky130_fd_sc_hd__buf_2
XANTENNA__17963__B1 _14608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25033__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15721__A HWDATA[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12650_ _12650_/A _12650_/B _12649_/X VGND VGND VPWR VPWR _12651_/A sky130_fd_sc_hd__or3_4
X_24636_ _24634_/CLK _16299_/X HRESETn VGND VGND VPWR VPWR _24636_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21442__B _21441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21848_ _14410_/Y _14212_/A _14433_/Y _22327_/B VGND VGND VPWR VPWR _21851_/C sky130_fd_sc_hd__o22a_4
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _12580_/Y _24885_/Q _12580_/Y _24885_/Q VGND VGND VPWR VPWR _12581_/X sky130_fd_sc_hd__a2bb2o_4
X_24567_ _24573_/CLK _24567_/D HRESETn VGND VGND VPWR VPWR _16485_/A sky130_fd_sc_hd__dfrtp_4
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21779_ _21756_/A _20076_/Y VGND VGND VPWR VPWR _21779_/X sky130_fd_sc_hd__or2_4
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14320_ _25168_/Q _14349_/A _14315_/X VGND VGND VPWR VPWR _14320_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__13241__A _13150_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23518_ _23912_/CLK _23518_/D VGND VGND VPWR VPWR _13335_/B sky130_fd_sc_hd__dfxtp_4
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24498_ _24460_/CLK _24498_/D HRESETn VGND VGND VPWR VPWR _16670_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_168_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _14251_/A VGND VGND VPWR VPWR _14251_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23449_ _24413_/CLK _20246_/X VGND VGND VPWR VPWR _20245_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_109_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23264__A1 _24443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ _13293_/A _13202_/B _13202_/C VGND VGND VPWR VPWR _13217_/B sky130_fd_sc_hd__or3_4
X_14182_ _14182_/A VGND VGND VPWR VPWR _14182_/X sky130_fd_sc_hd__buf_2
X_13133_ _13422_/A VGND VGND VPWR VPWR _13169_/A sky130_fd_sc_hd__buf_2
X_25119_ _25117_/CLK _14469_/X HRESETn VGND VGND VPWR VPWR _14467_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_151_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__23016__A1 _12804_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18990_ _18122_/B VGND VGND VPWR VPWR _18990_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13064_ _13085_/A _13064_/B _13064_/C VGND VGND VPWR VPWR _25348_/D sky130_fd_sc_hd__and3_4
X_17941_ _17944_/A _19140_/A VGND VGND VPWR VPWR _17942_/C sky130_fd_sc_hd__or2_4
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21578__A1 _21556_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12015_ _12014_/Y VGND VGND VPWR VPWR _12015_/X sky130_fd_sc_hd__buf_2
XFILLER_238_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17872_ _16908_/Y _17874_/B _17871_/Y VGND VGND VPWR VPWR _17872_/X sky130_fd_sc_hd__o21a_4
XANTENNA__23968__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19611_ _21951_/B _19607_/X _19610_/X _19607_/X VGND VGND VPWR VPWR _23679_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_41_0_HCLK clkbuf_7_41_0_HCLK/A VGND VGND VPWR VPWR clkbuf_8_83_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_16823_ _16820_/Y _16822_/X _15735_/X _16822_/X VGND VGND VPWR VPWR _16823_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19542_ _23700_/Q VGND VGND VPWR VPWR _19542_/Y sky130_fd_sc_hd__inv_2
X_13966_ _25233_/Q VGND VGND VPWR VPWR _14007_/A sky130_fd_sc_hd__buf_2
X_16754_ _16725_/A VGND VGND VPWR VPWR _16766_/A sky130_fd_sc_hd__buf_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15009__B2 _15008_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16206__B1 _11691_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22729__A _24595_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12917_ _12912_/A _12890_/X _12862_/X _12914_/B VGND VGND VPWR VPWR _12917_/X sky130_fd_sc_hd__a211o_4
X_15705_ _16539_/A _15836_/B VGND VGND VPWR VPWR _15736_/A sky130_fd_sc_hd__or2_4
X_16685_ _16668_/A VGND VGND VPWR VPWR _16685_/X sky130_fd_sc_hd__buf_2
X_19473_ _19472_/Y _19470_/X _11927_/X _19470_/X VGND VGND VPWR VPWR _23724_/D sky130_fd_sc_hd__a2bb2o_4
X_13897_ _13958_/B _13896_/Y VGND VGND VPWR VPWR _13897_/X sky130_fd_sc_hd__or2_4
XFILLER_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17954__B1 _18020_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21750__A1 _21119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18424_ _18424_/A _18424_/B _18424_/C _18423_/X VGND VGND VPWR VPWR _18424_/X sky130_fd_sc_hd__or4_4
XFILLER_222_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12848_ _12732_/Y _12848_/B VGND VGND VPWR VPWR _12848_/X sky130_fd_sc_hd__or2_4
X_15636_ _15636_/A _15636_/B _15636_/C _15636_/D VGND VGND VPWR VPWR _22111_/A sky130_fd_sc_hd__or4_4
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15567_ HWDATA[26] VGND VGND VPWR VPWR _15567_/X sky130_fd_sc_hd__buf_2
X_18355_ _18352_/Y _17476_/X _18354_/Y VGND VGND VPWR VPWR _18365_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__15992__A1_N _15980_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12779_ _12779_/A _12751_/X _12779_/C _12778_/X VGND VGND VPWR VPWR _12779_/X sky130_fd_sc_hd__or4_4
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14518_ _14510_/X _14517_/X _25116_/Q _14495_/Y VGND VGND VPWR VPWR _14518_/X sky130_fd_sc_hd__o22a_4
X_17306_ _17252_/D _17305_/X VGND VGND VPWR VPWR _17307_/B sky130_fd_sc_hd__or2_4
XFILLER_187_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24756__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15498_ _24942_/Q VGND VGND VPWR VPWR _15498_/Y sky130_fd_sc_hd__inv_2
X_18286_ _19597_/A _18280_/X _18285_/X VGND VGND VPWR VPWR _24219_/D sky130_fd_sc_hd__o21a_4
XFILLER_147_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14449_ _14447_/Y _14443_/X _14407_/X _14448_/X VGND VGND VPWR VPWR _25127_/D sky130_fd_sc_hd__a2bb2o_4
X_17237_ _24352_/Q VGND VGND VPWR VPWR _17237_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17168_ _16294_/Y _17292_/A _16294_/Y _17292_/A VGND VGND VPWR VPWR _17168_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11754__B1 _11753_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16119_ _16118_/Y _16116_/X _15951_/X _16116_/X VGND VGND VPWR VPWR _16119_/X sky130_fd_sc_hd__a2bb2o_4
X_17099_ _16984_/Y _17103_/A _17099_/C _17099_/D VGND VGND VPWR VPWR _17099_/X sky130_fd_sc_hd__or4_4
XANTENNA__16693__B1 _16420_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17293__A _17236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14710__A _14710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25544__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19809_ _23609_/Q VGND VGND VPWR VPWR _19809_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15799__A2 _15789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22820_ _17200_/A _21058_/X VGND VGND VPWR VPWR _22820_/X sky130_fd_sc_hd__or2_4
XFILLER_244_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__23191__B1 _24743_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_218_0_HCLK clkbuf_8_219_0_HCLK/A VGND VGND VPWR VPWR _24573_/CLK sky130_fd_sc_hd__clkbuf_1
X_22751_ _21305_/B _22750_/X _21312_/X _16035_/A _21708_/X VGND VGND VPWR VPWR _22751_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16637__A _16637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_225_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21702_ _21520_/X _21701_/X _21522_/X _24858_/Q _22522_/B VGND VGND VPWR VPWR _21703_/B
+ sky130_fd_sc_hd__a32o_4
XANTENNA__12281__A2_N _24831_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25470_ _25109_/CLK _12110_/X HRESETn VGND VGND VPWR VPWR _12109_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_197_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22682_ _22681_/X VGND VGND VPWR VPWR _22682_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20159__A _20158_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24421_ _24073_/CLK _16840_/X HRESETn VGND VGND VPWR VPWR _14917_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_240_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21633_ _21775_/A _21633_/B VGND VGND VPWR VPWR _21633_/X sky130_fd_sc_hd__or2_4
XFILLER_139_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24497__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24352_ _24667_/CLK _24352_/D HRESETn VGND VGND VPWR VPWR _24352_/Q sky130_fd_sc_hd__dfrtp_4
X_21564_ _21557_/Y _21558_/Y _21564_/C _21564_/D VGND VGND VPWR VPWR _21564_/X sky130_fd_sc_hd__or4_4
XFILLER_138_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23303_ _16796_/A _23138_/X _22801_/X _23302_/X VGND VGND VPWR VPWR _23304_/C sky130_fd_sc_hd__a211o_4
XANTENNA__24426__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20515_ _14266_/Y _20515_/B _24077_/Q VGND VGND VPWR VPWR _20519_/A sky130_fd_sc_hd__and3_4
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22805__C _22804_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24283_ _24275_/CLK _17801_/X HRESETn VGND VGND VPWR VPWR _24283_/Q sky130_fd_sc_hd__dfrtp_4
X_21495_ _21657_/A _21495_/B VGND VGND VPWR VPWR _21495_/X sky130_fd_sc_hd__or2_4
XFILLER_166_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21257__B1 _14672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23234_ _23120_/X _23232_/X _23123_/X _23233_/X VGND VGND VPWR VPWR _23235_/B sky130_fd_sc_hd__o22a_4
X_20446_ _20605_/A _20437_/C _20444_/B VGND VGND VPWR VPWR _20446_/X sky130_fd_sc_hd__o21a_4
XFILLER_106_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11745__B1 _11743_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23165_ _15566_/Y _23292_/B VGND VGND VPWR VPWR _23165_/X sky130_fd_sc_hd__and2_4
X_20377_ _20377_/A VGND VGND VPWR VPWR _20377_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__19870__B1 _19617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22821__B _22821_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22116_ _12099_/Y _21570_/X _18378_/Y _21571_/X VGND VGND VPWR VPWR _22116_/X sky130_fd_sc_hd__o22a_4
XFILLER_161_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23096_ _16103_/Y _22559_/X _22849_/X _11687_/Y _21051_/A VGND VGND VPWR VPWR _23096_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22047_ _14720_/Y _23685_/Q _22048_/A _19585_/X VGND VGND VPWR VPWR _22047_/X sky130_fd_sc_hd__o22a_4
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16436__B1 _16435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_28_0_HCLK clkbuf_6_29_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_57_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13820_ _13820_/A VGND VGND VPWR VPWR _13820_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23998_ _24074_/CLK _23998_/D HRESETn VGND VGND VPWR VPWR _23998_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13751_ _13733_/Y VGND VGND VPWR VPWR _14697_/A sky130_fd_sc_hd__buf_2
XFILLER_244_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22949_ _20916_/A _22829_/X _20776_/Y _22290_/A VGND VGND VPWR VPWR _22949_/X sky130_fd_sc_hd__o22a_4
XFILLER_90_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12473__A1 _12191_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12702_ _12696_/A _12696_/B VGND VGND VPWR VPWR _12703_/C sky130_fd_sc_hd__nand2_4
XFILLER_232_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16470_ _16470_/A VGND VGND VPWR VPWR _16470_/X sky130_fd_sc_hd__buf_2
XFILLER_216_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13682_ _13682_/A _13681_/X VGND VGND VPWR VPWR _13683_/A sky130_fd_sc_hd__and2_4
X_15421_ _13924_/A _15421_/B _13923_/D VGND VGND VPWR VPWR _15422_/A sky130_fd_sc_hd__or3_4
X_12633_ _12503_/Y _12633_/B VGND VGND VPWR VPWR _12634_/C sky130_fd_sc_hd__or2_4
X_24619_ _24618_/CLK _16342_/X HRESETn VGND VGND VPWR VPWR _24619_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15352_ _15352_/A _15350_/X _15352_/C VGND VGND VPWR VPWR _15352_/X sky130_fd_sc_hd__and3_4
X_18140_ _17981_/A _18138_/X _18139_/X VGND VGND VPWR VPWR _18140_/X sky130_fd_sc_hd__and3_4
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _12676_/A VGND VGND VPWR VPWR _12564_/Y sky130_fd_sc_hd__inv_2
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12802__A2_N _24800_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ _14295_/X _14302_/X _13468_/A _14300_/X VGND VGND VPWR VPWR _14303_/X sky130_fd_sc_hd__o22a_4
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18071_ _17981_/A _18069_/X _18070_/X VGND VGND VPWR VPWR _18071_/X sky130_fd_sc_hd__and3_4
XANTENNA__24167__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15283_ _15241_/A _15243_/B _15282_/X VGND VGND VPWR VPWR _25008_/D sky130_fd_sc_hd__and3_4
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ _13087_/A VGND VGND VPWR VPWR _13028_/A sky130_fd_sc_hd__inv_2
XFILLER_200_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17022_ _17022_/A _16965_/Y VGND VGND VPWR VPWR _17047_/C sky130_fd_sc_hd__or2_4
X_14234_ _14234_/A _14234_/B VGND VGND VPWR VPWR _15436_/A sky130_fd_sc_hd__or2_4
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21248__B1 _21247_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11736__B1 _11735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14165_ _14164_/X VGND VGND VPWR VPWR _14165_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13116_ _13116_/A _13116_/B VGND VGND VPWR VPWR _13117_/B sky130_fd_sc_hd__or2_4
XFILLER_125_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11751__A3 _15965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21628__A _22381_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14096_ _14096_/A _14096_/B _14095_/X VGND VGND VPWR VPWR _14097_/A sky130_fd_sc_hd__or3_4
X_18973_ _18972_/Y _14654_/A _17440_/X _14654_/A VGND VGND VPWR VPWR _23899_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__13489__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13047_ _12324_/Y _13046_/X VGND VGND VPWR VPWR _13047_/Y sky130_fd_sc_hd__nand2_4
X_17924_ _17924_/A VGND VGND VPWR VPWR _17924_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21347__B _22181_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16427__B1 _16059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17419__A1_N _17417_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17855_ _17854_/X VGND VGND VPWR VPWR _17856_/B sky130_fd_sc_hd__inv_2
XFILLER_227_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21971__A1 _21649_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20774__A2 _20708_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21971__B2 _21970_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16806_ _16806_/A VGND VGND VPWR VPWR _16806_/Y sky130_fd_sc_hd__inv_2
X_17786_ _17602_/B _17786_/B VGND VGND VPWR VPWR _17787_/A sky130_fd_sc_hd__or2_4
XFILLER_208_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14998_ _14998_/A VGND VGND VPWR VPWR _14998_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22459__A _16272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23173__B1 _23133_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19525_ _19524_/X VGND VGND VPWR VPWR _19526_/A sky130_fd_sc_hd__buf_2
XFILLER_35_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21363__A _14179_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16737_ _16737_/A VGND VGND VPWR VPWR _16737_/Y sky130_fd_sc_hd__inv_2
X_13949_ _13949_/A VGND VGND VPWR VPWR _13949_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_191_0_HCLK clkbuf_7_95_0_HCLK/X VGND VGND VPWR VPWR _25238_/CLK sky130_fd_sc_hd__clkbuf_1
X_19456_ _19597_/A _19939_/B _19455_/X VGND VGND VPWR VPWR _19456_/X sky130_fd_sc_hd__or3_4
XANTENNA__24937__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16668_ _16668_/A VGND VGND VPWR VPWR _16668_/X sky130_fd_sc_hd__buf_2
X_18407_ _18407_/A VGND VGND VPWR VPWR _18407_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_48_0_HCLK clkbuf_8_49_0_HCLK/A VGND VGND VPWR VPWR _25285_/CLK sky130_fd_sc_hd__clkbuf_1
X_15619_ _14403_/A VGND VGND VPWR VPWR _15619_/X sky130_fd_sc_hd__buf_2
X_19387_ _19387_/A _19163_/B _19320_/C VGND VGND VPWR VPWR _19388_/A sky130_fd_sc_hd__or3_4
XFILLER_201_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16599_ _16596_/Y _16592_/X _16597_/X _16598_/X VGND VGND VPWR VPWR _16599_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA_clkbuf_5_29_0_HCLK_A clkbuf_5_29_0_HCLK/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24590__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18338_ _19716_/C _18932_/B _19716_/C _18932_/B VGND VGND VPWR VPWR _18338_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22194__A _22194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_18269_ _18268_/Y _18265_/Y _16849_/X _18265_/Y VGND VGND VPWR VPWR _24223_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20300_ _20287_/Y VGND VGND VPWR VPWR _20300_/X sky130_fd_sc_hd__buf_2
XFILLER_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21280_ _22582_/A _21279_/X _13837_/Y _22582_/A VGND VGND VPWR VPWR _21280_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11727__B1 _11726_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20231_ _20231_/A VGND VGND VPWR VPWR _20231_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16666__B1 _16483_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20162_ _20161_/Y _20159_/X _20092_/X _20159_/X VGND VGND VPWR VPWR _20162_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21538__A _21537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22739__B1 _22423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20093_ _22218_/B _20088_/X _20092_/X _20088_/X VGND VGND VPWR VPWR _23505_/D sky130_fd_sc_hd__a2bb2o_4
X_24970_ _24959_/CLK _15440_/X HRESETn VGND VGND VPWR VPWR _13908_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_130_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23921_ _23912_/CLK _18916_/X VGND VGND VPWR VPWR _23921_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22754__A3 _22146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__17751__A _24261_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23852_ _25171_/CLK _19112_/X VGND VGND VPWR VPWR _23852_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22803_ _14998_/A _22661_/X _22802_/X VGND VGND VPWR VPWR _22803_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21273__A _14710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23783_ _24252_/CLK _19309_/X VGND VGND VPWR VPWR _19308_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20995_ _20496_/A _23962_/Q _13962_/A VGND VGND VPWR VPWR _23962_/D sky130_fd_sc_hd__a21o_4
XFILLER_26_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21714__A1 _21289_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12895__A _12895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25522_ _24236_/CLK _25522_/D HRESETn VGND VGND VPWR VPWR _25522_/Q sky130_fd_sc_hd__dfrtp_4
X_22734_ _22734_/A _22619_/B VGND VGND VPWR VPWR _22734_/X sky130_fd_sc_hd__and2_4
XFILLER_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24678__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25453_ _25453_/CLK _25453_/D HRESETn VGND VGND VPWR VPWR _12248_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_186_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24607__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22665_ _22725_/A _22665_/B _22665_/C _22665_/D VGND VGND VPWR VPWR _22665_/X sky130_fd_sc_hd__or4_4
XFILLER_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24404_ _24377_/CLK _24404_/D HRESETn VGND VGND VPWR VPWR _17050_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_71_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21616_ _21757_/A _21614_/X _21615_/X VGND VGND VPWR VPWR _21616_/X sky130_fd_sc_hd__and3_4
X_25384_ _25382_/CLK _25384_/D HRESETn VGND VGND VPWR VPWR _12740_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_200_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21720__B _21719_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22596_ _22632_/A _22595_/X VGND VGND VPWR VPWR _22596_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__24260__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24335_ _24340_/CLK _17407_/X HRESETn VGND VGND VPWR VPWR _21000_/B sky130_fd_sc_hd__dfstp_4
XFILLER_166_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21547_ _21545_/X _21546_/X _21111_/X VGND VGND VPWR VPWR _21547_/X sky130_fd_sc_hd__or3_4
XFILLER_154_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12280_ _12280_/A VGND VGND VPWR VPWR _12981_/C sky130_fd_sc_hd__inv_2
X_24266_ _24266_/CLK _17868_/Y HRESETn VGND VGND VPWR VPWR _24266_/Q sky130_fd_sc_hd__dfrtp_4
X_21478_ _17709_/A VGND VGND VPWR VPWR _21656_/A sky130_fd_sc_hd__buf_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22978__B1 _24737_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23217_ _23035_/X _23216_/X _23145_/X _24848_/Q _23037_/X VGND VGND VPWR VPWR _23217_/X
+ sky130_fd_sc_hd__a32o_4
X_20429_ _24069_/D _20429_/B VGND VGND VPWR VPWR _24068_/D sky130_fd_sc_hd__or2_4
XFILLER_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24197_ _25474_/CLK _24197_/D HRESETn VGND VGND VPWR VPWR _18376_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_106_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18646__B2 _24140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12391__B1 _12390_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23148_ _24811_/Q _23040_/X VGND VGND VPWR VPWR _23148_/X sky130_fd_sc_hd__or2_4
XANTENNA__21448__A _15780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15970_ _12198_/Y _15968_/X _15616_/X _15968_/X VGND VGND VPWR VPWR _24755_/D sky130_fd_sc_hd__a2bb2o_4
X_23079_ _24636_/Q _22817_/B _22817_/C VGND VGND VPWR VPWR _23079_/X sky130_fd_sc_hd__and3_4
XFILLER_0_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16409__B1 _16226_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14921_ _14921_/A VGND VGND VPWR VPWR _14921_/X sky130_fd_sc_hd__buf_2
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25412__CLK _24032_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17640_ _17569_/A _17645_/B _17593_/X VGND VGND VPWR VPWR _17640_/Y sky130_fd_sc_hd__a21oi_4
X_14852_ _14838_/X _14851_/Y _25047_/Q _14838_/X VGND VGND VPWR VPWR _25047_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13803_ _19570_/A _17410_/A VGND VGND VPWR VPWR _21958_/B sky130_fd_sc_hd__or2_4
X_14783_ _18020_/A _14656_/X _18020_/A _14656_/X VGND VGND VPWR VPWR _14783_/X sky130_fd_sc_hd__a2bb2o_4
X_17571_ _17502_/Y _17543_/Y _17570_/X VGND VGND VPWR VPWR _17571_/X sky130_fd_sc_hd__or3_4
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11995_ _11979_/A _11990_/A _11994_/Y VGND VGND VPWR VPWR _11995_/X sky130_fd_sc_hd__o21a_4
XANTENNA__21705__A1 _21581_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21705__B2 _21336_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19310_ _19310_/A VGND VGND VPWR VPWR _19310_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_8_201_0_HCLK clkbuf_8_201_0_HCLK/A VGND VGND VPWR VPWR _24591_/CLK sky130_fd_sc_hd__clkbuf_1
X_13734_ _13724_/X _13733_/Y _14683_/A _25279_/Q VGND VGND VPWR VPWR _13734_/X sky130_fd_sc_hd__and4_4
X_16522_ _14403_/A VGND VGND VPWR VPWR _16522_/X sky130_fd_sc_hd__buf_2
XFILLER_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_8_7_0_HCLK clkbuf_8_7_0_HCLK/A VGND VGND VPWR VPWR _23441_/CLK sky130_fd_sc_hd__clkbuf_1
X_19241_ _19240_/Y _19238_/X _16873_/X _19238_/X VGND VGND VPWR VPWR _23807_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__24348__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13665_ _13664_/Y _11853_/X VGND VGND VPWR VPWR _13681_/B sky130_fd_sc_hd__or2_4
X_16453_ _16453_/A VGND VGND VPWR VPWR _16454_/A sky130_fd_sc_hd__buf_2
XFILLER_188_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12616_ _12680_/A VGND VGND VPWR VPWR _12650_/A sky130_fd_sc_hd__inv_2
X_15404_ _15384_/X VGND VGND VPWR VPWR _15405_/B sky130_fd_sc_hd__inv_2
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__21469__B1 _17725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16384_ _24605_/Q VGND VGND VPWR VPWR _16384_/Y sky130_fd_sc_hd__inv_2
X_19172_ _23831_/Q VGND VGND VPWR VPWR _19172_/Y sky130_fd_sc_hd__inv_2
X_13596_ _13596_/A _13596_/B VGND VGND VPWR VPWR _13614_/A sky130_fd_sc_hd__and2_4
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16724__B _16792_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15335_ _15075_/Y _15338_/B _15334_/X VGND VGND VPWR VPWR _15335_/Y sky130_fd_sc_hd__a21oi_4
X_18123_ _18123_/A _18123_/B _18123_/C VGND VGND VPWR VPWR _18124_/C sky130_fd_sc_hd__and3_4
X_12547_ _24872_/Q VGND VGND VPWR VPWR _12547_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22681__A2 _22679_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15266_ _15269_/A _15266_/B _15265_/Y VGND VGND VPWR VPWR _25014_/D sky130_fd_sc_hd__and3_4
X_18054_ _18054_/A VGND VGND VPWR VPWR _18126_/A sky130_fd_sc_hd__buf_2
XFILLER_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12478_ _12197_/Y _12480_/B _12477_/Y VGND VGND VPWR VPWR _12478_/X sky130_fd_sc_hd__o21a_4
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__11709__B1 _25541_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14217_ _20664_/A VGND VGND VPWR VPWR _14217_/Y sky130_fd_sc_hd__inv_2
X_17005_ _16006_/Y _17023_/A _24736_/Q _17004_/Y VGND VGND VPWR VPWR _17005_/X sky130_fd_sc_hd__a2bb2o_4
X_15197_ _15187_/X VGND VGND VPWR VPWR _15201_/B sky130_fd_sc_hd__inv_2
XANTENNA__22433__A2 _21833_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23983__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14148_ _14088_/C _14102_/X _14088_/C _14102_/X VGND VGND VPWR VPWR _14149_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21641__B1 _21501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20995__A2 _23962_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14079_ _20541_/B _14536_/B _14058_/X _14005_/B _14073_/X VGND VGND VPWR VPWR _25228_/D
+ sky130_fd_sc_hd__a32o_4
X_18956_ _18955_/Y _14654_/X _17415_/X _14654_/X VGND VGND VPWR VPWR _23906_/D sky130_fd_sc_hd__a2bb2o_4
X_17907_ _17907_/A _17899_/Y VGND VGND VPWR VPWR _17907_/X sky130_fd_sc_hd__or2_4
XFILLER_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18887_ _18886_/X VGND VGND VPWR VPWR _18888_/A sky130_fd_sc_hd__buf_2
XFILLER_227_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17838_ _17758_/Y _17833_/B _17783_/X _17835_/B VGND VGND VPWR VPWR _17838_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_6_11_0_HCLK clkbuf_5_5_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_23_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17769_ _17769_/A VGND VGND VPWR VPWR _17769_/Y sky130_fd_sc_hd__inv_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19508_ _19502_/Y VGND VGND VPWR VPWR _19508_/X sky130_fd_sc_hd__buf_2
XANTENNA__24771__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20780_ _20780_/A VGND VGND VPWR VPWR _20780_/X sky130_fd_sc_hd__buf_2
XANTENNA__17376__A1 _17241_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24700__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19439_ _18039_/B VGND VGND VPWR VPWR _19439_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16915__A _16915_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24018__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22450_ _16366_/B VGND VGND VPWR VPWR _22450_/X sky130_fd_sc_hd__buf_2
XFILLER_22_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__21540__B _22130_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21401_ _14668_/X _21401_/B VGND VGND VPWR VPWR _21401_/X sky130_fd_sc_hd__or2_4
X_22381_ _22381_/A _20113_/Y VGND VGND VPWR VPWR _22381_/X sky130_fd_sc_hd__or2_4
XFILLER_136_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22672__A2 _22294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24120_ _25211_/CLK _24120_/D HRESETn VGND VGND VPWR VPWR _24120_/Q sky130_fd_sc_hd__dfstp_4
X_21332_ _24415_/Q _21325_/X _23001_/A _21331_/X VGND VGND VPWR VPWR _21333_/C sky130_fd_sc_hd__a211o_4
XFILLER_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21880__B1 _24262_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24051_ _24051_/CLK _24051_/D HRESETn VGND VGND VPWR VPWR _24051_/Q sky130_fd_sc_hd__dfrtp_4
X_21263_ _21884_/A _21263_/B VGND VGND VPWR VPWR _21263_/X sky130_fd_sc_hd__or2_4
XFILLER_237_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23002_ _23002_/A VGND VGND VPWR VPWR _23002_/X sky130_fd_sc_hd__buf_2
X_20214_ _20212_/Y _20213_/X _19708_/X _20213_/X VGND VGND VPWR VPWR _20214_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21194_ _24213_/Q _21192_/X _21193_/X VGND VGND VPWR VPWR _21194_/X sky130_fd_sc_hd__and3_4
XANTENNA__11794__A _11682_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20145_ _23487_/Q VGND VGND VPWR VPWR _20145_/Y sky130_fd_sc_hd__inv_2
XANTENNA__22188__A1 _21345_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24953_ _24953_/CLK _15473_/X HRESETn VGND VGND VPWR VPWR _24953_/Q sky130_fd_sc_hd__dfstp_4
X_20076_ _23510_/Q VGND VGND VPWR VPWR _20076_/Y sky130_fd_sc_hd__inv_2
XFILLER_246_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23904_ _25171_/CLK _23904_/D VGND VGND VPWR VPWR _18040_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_73_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24859__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24884_ _25428_/CLK _15715_/X HRESETn VGND VGND VPWR VPWR _24884_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16811__B1 _15725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23835_ _23827_/CLK _23835_/D VGND VGND VPWR VPWR _23835_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_122_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21699__B1 _25523_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11780_/A VGND VGND VPWR VPWR _14392_/A sky130_fd_sc_hd__buf_2
X_23766_ _24088_/CLK _19354_/X VGND VGND VPWR VPWR _18103_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22896__C1 _22895_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20978_ _14388_/Y _14369_/X VGND VGND VPWR VPWR _23927_/D sky130_fd_sc_hd__and2_4
XFILLER_26_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22360__A1 _21935_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22717_ _22704_/X _22708_/X _22712_/X _22716_/X VGND VGND VPWR VPWR _22717_/X sky130_fd_sc_hd__or4_4
X_25505_ _23691_/CLK _11921_/X HRESETn VGND VGND VPWR VPWR _19981_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__24441__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23697_ _23406_/CLK _19553_/X VGND VGND VPWR VPWR _19552_/A sky130_fd_sc_hd__dfxtp_4
XPHY_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ _11951_/A _13434_/X _13449_/X _25327_/Q _11950_/A VGND VGND VPWR VPWR _13450_/X
+ sky130_fd_sc_hd__o32a_4
X_25436_ _25444_/CLK _12489_/X HRESETn VGND VGND VPWR VPWR _12251_/A sky130_fd_sc_hd__dfrtp_4
Xclkbuf_8_31_0_HCLK clkbuf_8_31_0_HCLK/A VGND VGND VPWR VPWR _24310_/CLK sky130_fd_sc_hd__clkbuf_1
X_22648_ _22632_/Y _22637_/Y _22645_/Y _21445_/X _22647_/X VGND VGND VPWR VPWR _22648_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__22112__A1 _12781_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12401_ _12401_/A VGND VGND VPWR VPWR _12401_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_94_0_HCLK clkbuf_8_95_0_HCLK/A VGND VGND VPWR VPWR _24804_/CLK sky130_fd_sc_hd__clkbuf_1
X_13381_ _13445_/A _19753_/A VGND VGND VPWR VPWR _13383_/B sky130_fd_sc_hd__or2_4
X_25367_ _24819_/CLK _12969_/X HRESETn VGND VGND VPWR VPWR _21016_/A sky130_fd_sc_hd__dfrtp_4
X_22579_ _16765_/A _22534_/X _22535_/X VGND VGND VPWR VPWR _22579_/X sky130_fd_sc_hd__o21a_4
XFILLER_166_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21320__C1 _21319_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15120_ _15120_/A VGND VGND VPWR VPWR _15120_/Y sky130_fd_sc_hd__inv_2
X_12332_ _24821_/Q VGND VGND VPWR VPWR _12332_/Y sky130_fd_sc_hd__inv_2
X_24318_ _24390_/CLK _24318_/D HRESETn VGND VGND VPWR VPWR _17494_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_166_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25298_ _25308_/CLK _25298_/D HRESETn VGND VGND VPWR VPWR _25298_/Q sky130_fd_sc_hd__dfrtp_4
X_15051_ _14879_/Y _15185_/A _15017_/X _15050_/X VGND VGND VPWR VPWR _15051_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12263_ _12263_/A VGND VGND VPWR VPWR _12413_/A sky130_fd_sc_hd__buf_2
X_24249_ _23890_/CLK _24249_/D HRESETn VGND VGND VPWR VPWR _24249_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__23073__C1 _23072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14002_ _14019_/D _14002_/B VGND VGND VPWR VPWR _14536_/A sky130_fd_sc_hd__nor2_4
XANTENNA__22281__B _22280_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12194_ _25457_/Q VGND VGND VPWR VPWR _12194_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18810_ _18810_/A VGND VGND VPWR VPWR _18811_/B sky130_fd_sc_hd__inv_2
XANTENNA__15176__A _15165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19790_ _19788_/Y _19784_/X _19746_/X _19789_/X VGND VGND VPWR VPWR _23616_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18741_ _18695_/X _18705_/X _18728_/A VGND VGND VPWR VPWR _18741_/X sky130_fd_sc_hd__o21a_4
XFILLER_95_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15953_ HWDATA[17] VGND VGND VPWR VPWR _15953_/X sky130_fd_sc_hd__buf_2
XFILLER_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11854__D _11853_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14904_ _14903_/X _16852_/A _14903_/X _16852_/A VGND VGND VPWR VPWR _14905_/D sky130_fd_sc_hd__a2bb2o_4
X_18672_ _18744_/A VGND VGND VPWR VPWR _18734_/A sky130_fd_sc_hd__buf_2
X_15884_ _15879_/X _15880_/X _16229_/A _22714_/A _15881_/X VGND VGND VPWR VPWR _15884_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16802__B1 _16467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17623_ _17620_/A _17615_/X _17622_/X VGND VGND VPWR VPWR _24314_/D sky130_fd_sc_hd__and3_4
XANTENNA__24529__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14835_ _23993_/D _14834_/Y _25197_/Q _23993_/D VGND VGND VPWR VPWR _14835_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17554_ _17554_/A _17539_/X _17547_/X _17553_/X VGND VGND VPWR VPWR _17555_/B sky130_fd_sc_hd__or4_4
X_11978_ _24093_/Q _11977_/X VGND VGND VPWR VPWR _11990_/A sky130_fd_sc_hd__and2_4
X_14766_ _14775_/A _14757_/X _14776_/B VGND VGND VPWR VPWR _14766_/X sky130_fd_sc_hd__o21a_4
XFILLER_205_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16505_ _24559_/Q VGND VGND VPWR VPWR _16505_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24182__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13717_ _13669_/X _13716_/Y _13667_/X _13700_/X _11840_/A VGND VGND VPWR VPWR _25283_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_60_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14697_ _14697_/A _14664_/X _14692_/X _14696_/X VGND VGND VPWR VPWR _14697_/X sky130_fd_sc_hd__or4_4
X_17485_ _17485_/A VGND VGND VPWR VPWR _17485_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19224_ _19224_/A VGND VGND VPWR VPWR _19224_/X sky130_fd_sc_hd__buf_2
XANTENNA__22918__A1_N _17251_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24111__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16436_ _15110_/Y _16430_/X _16435_/X _16430_/X VGND VGND VPWR VPWR _24582_/D sky130_fd_sc_hd__a2bb2o_4
X_13648_ _24046_/Q _13648_/B VGND VGND VPWR VPWR _13648_/X sky130_fd_sc_hd__or2_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21544__A1_N _21532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19155_ _18158_/B VGND VGND VPWR VPWR _19155_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18372__D _18372_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13579_ _14608_/A _13579_/B VGND VGND VPWR VPWR _13579_/X sky130_fd_sc_hd__or2_4
X_16367_ _16366_/X VGND VGND VPWR VPWR _16792_/B sky130_fd_sc_hd__buf_2
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_2_0_HCLK clkbuf_5_3_0_HCLK/A VGND VGND VPWR VPWR clkbuf_5_2_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_18106_ _18032_/A _19310_/A VGND VGND VPWR VPWR _18108_/B sky130_fd_sc_hd__or2_4
XANTENNA__25388__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15318_ _15304_/C _15315_/X VGND VGND VPWR VPWR _15318_/X sky130_fd_sc_hd__or2_4
XFILLER_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16298_ _16284_/X VGND VGND VPWR VPWR _16298_/X sky130_fd_sc_hd__buf_2
X_19086_ _19074_/A VGND VGND VPWR VPWR _19086_/X sky130_fd_sc_hd__buf_2
XFILLER_172_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18037_ _17987_/X _18037_/B VGND VGND VPWR VPWR _18038_/C sky130_fd_sc_hd__or2_4
XFILLER_172_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15249_ _15249_/A _15247_/A VGND VGND VPWR VPWR _15249_/X sky130_fd_sc_hd__or2_4
XFILLER_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__21088__A _21088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21090__A1 _24781_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19988_ _19988_/A VGND VGND VPWR VPWR _22344_/B sky130_fd_sc_hd__inv_2
XFILLER_86_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18939_ _18947_/A VGND VGND VPWR VPWR _18939_/X sky130_fd_sc_hd__buf_2
XANTENNA__21917__A1 _21901_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21950_ _22343_/A _21950_/B VGND VGND VPWR VPWR _21952_/B sky130_fd_sc_hd__or2_4
XFILLER_227_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20901_ _20892_/X _20900_/X _24495_/Q _20896_/X VGND VGND VPWR VPWR _24051_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21881_ _25437_/Q _23277_/A _21880_/X _21111_/X VGND VGND VPWR VPWR _21881_/X sky130_fd_sc_hd__a211o_4
X_23620_ _23859_/CLK _23620_/D VGND VGND VPWR VPWR _23620_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13334__A _13334_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20832_ _16713_/Y _20825_/X _20828_/X _20831_/Y VGND VGND VPWR VPWR _20833_/A sky130_fd_sc_hd__o22a_4
XFILLER_199_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23551_ _23534_/CLK _19975_/X VGND VGND VPWR VPWR _19973_/A sky130_fd_sc_hd__dfxtp_4
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20763_ _13107_/A VGND VGND VPWR VPWR _20764_/C sky130_fd_sc_hd__inv_2
XANTENNA__20353__B1 _19603_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22502_ _22500_/X _22502_/B _22876_/C VGND VGND VPWR VPWR _22502_/X sky130_fd_sc_hd__or3_4
XFILLER_210_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23482_ _23497_/CLK _23482_/D VGND VGND VPWR VPWR _20156_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_18_0_HCLK clkbuf_6_9_0_HCLK/X VGND VGND VPWR VPWR clkbuf_8_37_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20694_ _15632_/Y _20687_/X _20690_/X _20693_/Y VGND VGND VPWR VPWR _20695_/A sky130_fd_sc_hd__o22a_4
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25221_ _25113_/CLK _25221_/D HRESETn VGND VGND VPWR VPWR _14106_/A sky130_fd_sc_hd__dfrtp_4
X_22433_ _16339_/Y _21833_/X _22432_/X _16052_/Y _22274_/X VGND VGND VPWR VPWR _22433_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_183_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25152_ _23926_/CLK _14376_/X HRESETn VGND VGND VPWR VPWR _25152_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22364_ _22385_/A _22364_/B VGND VGND VPWR VPWR _22366_/B sky130_fd_sc_hd__or2_4
XANTENNA__22382__A _22379_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24103_ _24325_/CLK _20972_/X HRESETn VGND VGND VPWR VPWR _24103_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__25058__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21315_ _21303_/X VGND VGND VPWR VPWR _21315_/X sky130_fd_sc_hd__buf_2
XFILLER_164_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25083_ _25098_/CLK _14601_/X HRESETn VGND VGND VPWR VPWR _25083_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15532__B1 HADDR[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22295_ _22295_/A _22420_/B VGND VGND VPWR VPWR _22295_/X sky130_fd_sc_hd__or2_4
XFILLER_191_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24034_ _24910_/CLK _24034_/D HRESETn VGND VGND VPWR VPWR _13126_/A sky130_fd_sc_hd__dfrtp_4
X_21246_ _21627_/A _21243_/X _21245_/X VGND VGND VPWR VPWR _21246_/X sky130_fd_sc_hd__and3_4
XFILLER_104_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17285__B1 _17255_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21177_ _21177_/A VGND VGND VPWR VPWR _21178_/A sky130_fd_sc_hd__inv_2
XFILLER_238_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15835__B2 _15786_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20128_ _20116_/A VGND VGND VPWR VPWR _20128_/X sky130_fd_sc_hd__buf_2
XFILLER_58_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11674__D _15640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12950_ _12762_/Y _12952_/B _12949_/Y VGND VGND VPWR VPWR _12950_/X sky130_fd_sc_hd__o21a_4
XFILLER_46_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15724__A _15724_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24693__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20059_ _20053_/X _18328_/X _15830_/X _13299_/B _20055_/X VGND VGND VPWR VPWR _23519_/D
+ sky130_fd_sc_hd__a32o_4
X_24936_ _23476_/CLK _15515_/X HRESETn VGND VGND VPWR VPWR _11673_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_246_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11901_ _19603_/A VGND VGND VPWR VPWR _11901_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24622__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12881_ _12759_/Y _12885_/B _12862_/X _12878_/B VGND VGND VPWR VPWR _12881_/X sky130_fd_sc_hd__a211o_4
XANTENNA__15599__B1 _11735_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24867_ _24866_/CLK _15747_/X HRESETn VGND VGND VPWR VPWR _24867_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _11832_/A VGND VGND VPWR VPWR _11832_/Y sky130_fd_sc_hd__inv_2
X_14620_ _14612_/X _14619_/Y _25081_/Q _14611_/Y VGND VGND VPWR VPWR _25081_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_45_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23818_ _23754_/CLK _23818_/D VGND VGND VPWR VPWR _19207_/A sky130_fd_sc_hd__dfxtp_4
X_24798_ _24800_/CLK _15885_/X HRESETn VGND VGND VPWR VPWR _24798_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_199_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21136__A2 _14182_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _13560_/Y _14550_/X VGND VGND VPWR VPWR _14551_/X sky130_fd_sc_hd__or2_4
XFILLER_202_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _25526_/Q VGND VGND VPWR VPWR _11763_/Y sky130_fd_sc_hd__inv_2
X_23749_ _24889_/CLK _19404_/X VGND VGND VPWR VPWR _23749_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_187_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__20344__B1 _19620_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19569__C _13765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13501_/Y _13499_/X _12076_/X _13499_/X VGND VGND VPWR VPWR _13502_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12788__A1_N _12920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14481_/Y _14475_/X _14389_/X _14468_/A VGND VGND VPWR VPWR _25114_/D sky130_fd_sc_hd__a2bb2o_4
X_17270_ _17270_/A VGND VGND VPWR VPWR _24371_/D sky130_fd_sc_hd__inv_2
XPHY_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _25542_/Q VGND VGND VPWR VPWR _11694_/Y sky130_fd_sc_hd__inv_2
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13433_ _13433_/A _13429_/X _13432_/X VGND VGND VPWR VPWR _13434_/C sky130_fd_sc_hd__or3_4
X_16221_ _22806_/A VGND VGND VPWR VPWR _16221_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25419_ _25409_/CLK _25419_/D HRESETn VGND VGND VPWR VPWR _25419_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25481__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16152_ _22153_/A VGND VGND VPWR VPWR _16152_/Y sky130_fd_sc_hd__inv_2
X_13364_ _13396_/A _23909_/Q VGND VGND VPWR VPWR _13365_/C sky130_fd_sc_hd__or2_4
XFILLER_127_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__25410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12315_ _12315_/A VGND VGND VPWR VPWR _12315_/Y sky130_fd_sc_hd__inv_2
X_15103_ _25005_/Q VGND VGND VPWR VPWR _15304_/C sky130_fd_sc_hd__inv_2
XFILLER_6_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16083_ _11697_/Y _22505_/B VGND VGND VPWR VPWR _16084_/A sky130_fd_sc_hd__and2_4
X_13295_ _13392_/A _23911_/Q VGND VGND VPWR VPWR _13296_/C sky130_fd_sc_hd__or2_4
XFILLER_170_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15034_ _15204_/B _16763_/A _15204_/B _16763_/A VGND VGND VPWR VPWR _15034_/X sky130_fd_sc_hd__a2bb2o_4
X_19911_ _23573_/Q VGND VGND VPWR VPWR _19911_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16721__C _22539_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12246_ _12278_/A _23144_/A _12248_/A _12245_/Y VGND VGND VPWR VPWR _12246_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19842_ _19842_/A VGND VGND VPWR VPWR _19842_/Y sky130_fd_sc_hd__inv_2
X_12177_ _12428_/C _24764_/Q _12176_/A _24764_/Q VGND VGND VPWR VPWR _12186_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19773_ _19773_/A VGND VGND VPWR VPWR _21755_/B sky130_fd_sc_hd__inv_2
X_16985_ _24734_/Q _24391_/Q _16027_/Y _16984_/Y VGND VGND VPWR VPWR _16986_/D sky130_fd_sc_hd__o22a_4
XFILLER_209_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18724_ _18735_/A VGND VGND VPWR VPWR _18724_/X sky130_fd_sc_hd__buf_2
XFILLER_49_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15936_ _12182_/Y _15932_/X _15564_/X _15935_/X VGND VGND VPWR VPWR _15936_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18010__A _18090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24363__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18655_ _16564_/Y _24148_/Q _24525_/Q _18789_/C VGND VGND VPWR VPWR _18655_/X sky130_fd_sc_hd__a2bb2o_4
X_15867_ _15843_/X _15850_/X _15719_/X _24811_/Q _15857_/X VGND VGND VPWR VPWR _15867_/X
+ sky130_fd_sc_hd__a32o_4
X_17606_ _17606_/A VGND VGND VPWR VPWR _24319_/D sky130_fd_sc_hd__inv_2
XANTENNA__24123__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14818_ _14817_/X _14805_/A VGND VGND VPWR VPWR _14818_/X sky130_fd_sc_hd__and2_4
X_18586_ _18585_/X VGND VGND VPWR VPWR _24162_/D sky130_fd_sc_hd__inv_2
X_15798_ _15777_/X _15789_/X _15719_/X _24846_/Q _15787_/X VGND VGND VPWR VPWR _24846_/D
+ sky130_fd_sc_hd__a32o_4
XFILLER_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17537_ _11720_/Y _24308_/Q _25541_/Q _17502_/Y VGND VGND VPWR VPWR _17539_/C sky130_fd_sc_hd__a2bb2o_4
X_14749_ _21764_/A _14747_/X _14748_/Y VGND VGND VPWR VPWR _25062_/D sky130_fd_sc_hd__o21a_4
XANTENNA__20335__B1 _19606_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17468_ _13179_/A _17467_/X _13179_/A _17467_/X VGND VGND VPWR VPWR _17487_/B sky130_fd_sc_hd__a2bb2o_4
X_19207_ _19207_/A VGND VGND VPWR VPWR _19207_/Y sky130_fd_sc_hd__inv_2
X_16419_ _16417_/Y _16418_/X _16240_/X _16418_/X VGND VGND VPWR VPWR _24591_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__22088__B1 _14710_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22627__A2 _22432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19776__A _19764_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17399_ _17399_/A _17399_/B VGND VGND VPWR VPWR _17399_/X sky130_fd_sc_hd__or2_4
XFILLER_158_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19138_ _17440_/A VGND VGND VPWR VPWR _19138_/X sky130_fd_sc_hd__buf_2
XANTENNA__25151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19069_ _23867_/Q VGND VGND VPWR VPWR _19069_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21100_ _15851_/X VGND VGND VPWR VPWR _21101_/A sky130_fd_sc_hd__buf_2
X_22080_ _22379_/A _20071_/Y VGND VGND VPWR VPWR _22081_/C sky130_fd_sc_hd__or2_4
XFILLER_160_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21031_ _22730_/A VGND VGND VPWR VPWR _21031_/X sky130_fd_sc_hd__buf_2
XFILLER_113_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22982_ _22774_/X _22979_/Y _22868_/X _22981_/X VGND VGND VPWR VPWR _22982_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21933_ _21933_/A _21933_/B _21933_/C VGND VGND VPWR VPWR _21933_/X sky130_fd_sc_hd__and3_4
X_24721_ _24737_/CLK _24721_/D HRESETn VGND VGND VPWR VPWR _24721_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13064__A _13085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24033__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24652_ _24654_/CLK _24652_/D HRESETn VGND VGND VPWR VPWR _22097_/A sky130_fd_sc_hd__dfrtp_4
X_21864_ _15022_/A _21864_/B _21864_/C VGND VGND VPWR VPWR _21864_/X sky130_fd_sc_hd__and3_4
XANTENNA__16888__A2_N _23320_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_231_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14253__B1 _13829_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23603_ _23494_/CLK _19830_/X VGND VGND VPWR VPWR _19829_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_70_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__21281__A _25057_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20815_ _20813_/Y _20810_/X _20814_/X VGND VGND VPWR VPWR _20815_/X sky130_fd_sc_hd__o21a_4
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24583_ _24980_/CLK _24583_/D HRESETn VGND VGND VPWR VPWR _16432_/A sky130_fd_sc_hd__dfrtp_4
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21795_ _21662_/A _20022_/Y VGND VGND VPWR VPWR _21795_/X sky130_fd_sc_hd__or2_4
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19192__B1 _19125_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23534_ _23534_/CLK _23534_/D VGND VGND VPWR VPWR _20022_/A sky130_fd_sc_hd__dfxtp_4
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20746_ _20744_/Y _20741_/Y _20749_/A VGND VGND VPWR VPWR _20746_/X sky130_fd_sc_hd__o21a_4
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25239__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23465_ _23754_/CLK _23465_/D VGND VGND VPWR VPWR _17980_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__15753__B1 _15752_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20677_ _20495_/C VGND VGND VPWR VPWR _20677_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25204_ _25204_/CLK _14202_/X HRESETn VGND VGND VPWR VPWR _14201_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_7_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22416_ _16699_/Y _22416_/B VGND VGND VPWR VPWR _22416_/X sky130_fd_sc_hd__and2_4
XFILLER_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23396_ _23425_/CLK _23396_/D VGND VGND VPWR VPWR _23396_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_148_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_8_105_0_HCLK clkbuf_7_52_0_HCLK/X VGND VGND VPWR VPWR _24618_/CLK sky130_fd_sc_hd__clkbuf_1
X_25135_ _25134_/CLK _14432_/X HRESETn VGND VGND VPWR VPWR _25135_/Q sky130_fd_sc_hd__dfstp_4
X_22347_ _21936_/A _19918_/Y VGND VGND VPWR VPWR _22348_/C sky130_fd_sc_hd__or2_4
XANTENNA__15719__A HWDATA[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_168_0_HCLK clkbuf_7_84_0_HCLK/X VGND VGND VPWR VPWR _23767_/CLK sky130_fd_sc_hd__clkbuf_1
X_12100_ _12099_/Y _12095_/X _11770_/X _12095_/X VGND VGND VPWR VPWR _12100_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13080_ _13074_/A _13074_/B VGND VGND VPWR VPWR _13081_/C sky130_fd_sc_hd__nand2_4
X_25066_ _25070_/CLK _14736_/X HRESETn VGND VGND VPWR VPWR _22043_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_163_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22278_ _22141_/X VGND VGND VPWR VPWR _22946_/A sky130_fd_sc_hd__buf_2
XANTENNA__22840__A _22840_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12031_ _24099_/Q _12014_/A _25488_/Q _12027_/X VGND VGND VPWR VPWR _12031_/X sky130_fd_sc_hd__o22a_4
X_24017_ _24049_/CLK _24017_/D HRESETn VGND VGND VPWR VPWR _13121_/D sky130_fd_sc_hd__dfrtp_4
X_21229_ _16715_/Y _21124_/B VGND VGND VPWR VPWR _21235_/B sky130_fd_sc_hd__or2_4
XANTENNA__24874__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__21456__A _21463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24803__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13819__B1 _13818_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16770_ _15008_/Y _16766_/X _16597_/X _16769_/X VGND VGND VPWR VPWR _16770_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13982_ _14001_/A _14022_/B _14012_/A _13981_/X VGND VGND VPWR VPWR _13982_/X sky130_fd_sc_hd__or4_4
X_15721_ HWDATA[25] VGND VGND VPWR VPWR _15721_/X sky130_fd_sc_hd__buf_2
XFILLER_218_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12933_ _12932_/X VGND VGND VPWR VPWR _12934_/B sky130_fd_sc_hd__inv_2
X_24919_ _24032_/CLK _15568_/X HRESETn VGND VGND VPWR VPWR _15566_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_218_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18440_ _24186_/Q VGND VGND VPWR VPWR _18440_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__17430__B1 _16849_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15652_ _15648_/X VGND VGND VPWR VPWR _21089_/B sky130_fd_sc_hd__buf_2
X_12864_ _12864_/A VGND VGND VPWR VPWR _25396_/D sky130_fd_sc_hd__inv_2
XPHY_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22287__A _21597_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14602_/Y _14610_/A _25081_/Q _13623_/X VGND VGND VPWR VPWR _14619_/A sky130_fd_sc_hd__o22a_4
X_11815_ _11814_/Y _24233_/Q _11814_/Y _24233_/Q VGND VGND VPWR VPWR _11815_/X sky130_fd_sc_hd__a2bb2o_4
X_18371_ _18371_/A VGND VGND VPWR VPWR _18371_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20317__B1 _15762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _22667_/A _24798_/Q _22667_/A _24798_/Q VGND VGND VPWR VPWR _12803_/A sky130_fd_sc_hd__a2bb2o_4
X_15583_ _15583_/A VGND VGND VPWR VPWR _15583_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15992__B1 _15991_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17200_/A _17322_/B VGND VGND VPWR VPWR _17323_/C sky130_fd_sc_hd__or2_4
XFILLER_187_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__20868__A1 _16694_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _25531_/Q VGND VGND VPWR VPWR _11746_/Y sky130_fd_sc_hd__inv_2
X_14534_ _14030_/Y _14038_/X _14534_/C _14043_/Y VGND VGND VPWR VPWR _14535_/B sky130_fd_sc_hd__or4_4
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18930__B1 _17440_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _17244_/X _17252_/X VGND VGND VPWR VPWR _17253_/X sky130_fd_sc_hd__or2_4
XFILLER_147_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _11700_/A VGND VGND VPWR VPWR _21519_/A sky130_fd_sc_hd__buf_2
X_14465_ _25120_/Q VGND VGND VPWR VPWR _14465_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15744__B1 _24868_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16204_ _16202_/Y _16198_/X _15939_/X _16203_/X VGND VGND VPWR VPWR _16204_/X sky130_fd_sc_hd__a2bb2o_4
X_13416_ _13310_/X _13412_/X _13416_/C VGND VGND VPWR VPWR _13416_/X sky130_fd_sc_hd__or3_4
Xclkbuf_7_64_0_HCLK clkbuf_7_65_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_64_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14396_ _14395_/X VGND VGND VPWR VPWR _14442_/B sky130_fd_sc_hd__buf_2
X_17184_ _24636_/Q _23078_/A _16297_/Y _17183_/Y VGND VGND VPWR VPWR _17184_/X sky130_fd_sc_hd__o22a_4
X_13347_ _13312_/A _19727_/A VGND VGND VPWR VPWR _13347_/X sky130_fd_sc_hd__or2_4
X_16135_ _22602_/A VGND VGND VPWR VPWR _16135_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13278_ _13350_/A _23616_/Q VGND VGND VPWR VPWR _13278_/X sky130_fd_sc_hd__or2_4
X_16066_ _16064_/Y _16058_/X _15466_/X _16065_/X VGND VGND VPWR VPWR _16066_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__16966__A1_N _24737_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12229_ _12229_/A VGND VGND VPWR VPWR _12275_/A sky130_fd_sc_hd__inv_2
X_15017_ _15017_/A _14997_/X _15017_/C _15017_/D VGND VGND VPWR VPWR _15017_/X sky130_fd_sc_hd__or4_4
XANTENNA__17844__A _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19825_ _21605_/B _19823_/X _19824_/X _19823_/X VGND VGND VPWR VPWR _23605_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24544__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19756_ _19756_/A VGND VGND VPWR VPWR _19756_/Y sky130_fd_sc_hd__inv_2
X_16968_ _16968_/A _16963_/X _16966_/X _16967_/X VGND VGND VPWR VPWR _16987_/B sky130_fd_sc_hd__or4_4
XANTENNA__24099__D MSI_S2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22545__A1 _17347_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18707_ _18707_/A _18707_/B _18707_/C VGND VGND VPWR VPWR _18707_/X sky130_fd_sc_hd__or3_4
X_15919_ _15651_/X _15829_/X _15838_/X _24781_/Q _15918_/X VGND VGND VPWR VPWR _15919_/X
+ sky130_fd_sc_hd__a32o_4
X_19687_ _13404_/B VGND VGND VPWR VPWR _19687_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16899_ _22980_/A _17817_/A _23193_/A _16898_/Y VGND VGND VPWR VPWR _16899_/X sky130_fd_sc_hd__a2bb2o_4
X_18638_ _18638_/A _18638_/B _18627_/X _18637_/X VGND VGND VPWR VPWR _18638_/X sky130_fd_sc_hd__or4_4
XFILLER_80_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22197__A _22197_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18569_ _18473_/Y _18568_/X _18489_/X VGND VGND VPWR VPWR _18569_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20600_ _20600_/A _20600_/B VGND VGND VPWR VPWR _20600_/Y sky130_fd_sc_hd__nor2_4
XFILLER_178_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21580_ _14932_/Y _15704_/A _21582_/A _21579_/X VGND VGND VPWR VPWR _21580_/X sky130_fd_sc_hd__o22a_4
XANTENNA__18921__B1 _16778_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25332__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20531_ _24075_/Q _20535_/B _20503_/X VGND VGND VPWR VPWR _20531_/X sky130_fd_sc_hd__a21o_4
XFILLER_221_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23250_ _24544_/Q _22282_/X _15663_/X _23249_/X VGND VGND VPWR VPWR _23250_/X sky130_fd_sc_hd__a211o_4
X_20462_ _20462_/A _14052_/A VGND VGND VPWR VPWR _20463_/B sky130_fd_sc_hd__and2_4
X_22201_ _22209_/A _20118_/Y VGND VGND VPWR VPWR _22204_/B sky130_fd_sc_hd__or2_4
XFILLER_180_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23181_ _23213_/A _23181_/B _23181_/C VGND VGND VPWR VPWR _23182_/D sky130_fd_sc_hd__and3_4
XFILLER_146_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15539__A _11706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20393_ _13256_/B VGND VGND VPWR VPWR _20393_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14443__A _14455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22132_ _24484_/Q _22132_/B VGND VGND VPWR VPWR _22135_/B sky130_fd_sc_hd__or2_4
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16160__B1 _15976_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22063_ _22365_/A _22063_/B VGND VGND VPWR VPWR _22063_/X sky130_fd_sc_hd__or2_4
XFILLER_245_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22233__B1 _22231_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21014_ _21066_/A _21014_/B VGND VGND VPWR VPWR _21014_/X sky130_fd_sc_hd__and2_4
XFILLER_114_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__24285__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__20180__A _20180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24214__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_247_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22965_ _22942_/X _22965_/B _22957_/X _22965_/D VGND VGND VPWR VPWR HRDATA[20] sky130_fd_sc_hd__or4_4
XFILLER_56_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24704_ _24704_/CLK _16107_/X HRESETn VGND VGND VPWR VPWR _23049_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_83_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21916_ _22228_/A _21908_/X _21915_/X VGND VGND VPWR VPWR _21916_/X sky130_fd_sc_hd__or3_4
X_22896_ _22873_/X _22876_/X _22880_/Y _22895_/X VGND VGND VPWR VPWR HRDATA[18] sky130_fd_sc_hd__a211o_4
XANTENNA__14226__B1 _13791_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21847_ _21847_/A _22119_/B VGND VGND VPWR VPWR _21847_/Y sky130_fd_sc_hd__nand2_4
X_24635_ _24634_/CLK _24635_/D HRESETn VGND VGND VPWR VPWR _24635_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__15974__B1 _24752_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _25431_/Q VGND VGND VPWR VPWR _12580_/Y sky130_fd_sc_hd__inv_2
X_24566_ _24540_/CLK _24566_/D HRESETn VGND VGND VPWR VPWR _24566_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21778_ _21775_/A _21778_/B VGND VGND VPWR VPWR _21778_/X sky130_fd_sc_hd__or2_4
XFILLER_196_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25073__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14529__A1 scl_oen_o_S4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20729_ _15610_/Y _20708_/X _20716_/X _20728_/X VGND VGND VPWR VPWR _20729_/X sky130_fd_sc_hd__o22a_4
X_23517_ _23388_/CLK _20062_/X VGND VGND VPWR VPWR _13367_/B sky130_fd_sc_hd__dfxtp_4
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15726__B1 _24878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24497_ _24427_/CLK _16674_/X HRESETn VGND VGND VPWR VPWR _24497_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_196_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16833__A _24425_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__25002__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _14249_/Y _14247_/X _13826_/X _14247_/X VGND VGND VPWR VPWR _14250_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23448_ _23490_/CLK _20249_/X VGND VGND VPWR VPWR _20247_/A sky130_fd_sc_hd__dfxtp_4
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__23264__A2 _21542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _13254_/A _13201_/B _13201_/C VGND VGND VPWR VPWR _13202_/C sky130_fd_sc_hd__and3_4
XANTENNA__21275__A1 _21258_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14181_ _14181_/A VGND VGND VPWR VPWR _14182_/A sky130_fd_sc_hd__buf_2
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23379_ _23859_/CLK _23379_/D VGND VGND VPWR VPWR _23379_/Q sky130_fd_sc_hd__dfxtp_4
X_13132_ _13247_/A VGND VGND VPWR VPWR _13422_/A sky130_fd_sc_hd__buf_2
XANTENNA__12960__B1 _12854_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25118_ _25117_/CLK _25118_/D HRESETn VGND VGND VPWR VPWR _25118_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16151__B1 _16059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13063_ _12340_/Y _13063_/B VGND VGND VPWR VPWR _13064_/C sky130_fd_sc_hd__or2_4
X_17940_ _17940_/A _23850_/Q VGND VGND VPWR VPWR _17940_/X sky130_fd_sc_hd__or2_4
X_25049_ _25052_/CLK _14846_/X HRESETn VGND VGND VPWR VPWR _14796_/A sky130_fd_sc_hd__dfrtp_4
XANTENNA__17664__A _17559_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21578__A2 _21564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12014_ _12014_/A VGND VGND VPWR VPWR _12014_/Y sky130_fd_sc_hd__inv_2
X_17871_ _16908_/Y _17874_/B _16952_/X VGND VGND VPWR VPWR _17871_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_239_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_6_0_HCLK clkbuf_4_6_0_HCLK/A VGND VGND VPWR VPWR clkbuf_4_6_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19610_ _19610_/A VGND VGND VPWR VPWR _19610_/X sky130_fd_sc_hd__buf_2
X_16822_ _16841_/A VGND VGND VPWR VPWR _16822_/X sky130_fd_sc_hd__buf_2
XFILLER_48_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__12601__A _25411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19541_ _19538_/Y _19539_/X _19540_/X _19539_/X VGND VGND VPWR VPWR _19541_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16753_ _15025_/Y _16749_/X _16402_/X _16749_/X VGND VGND VPWR VPWR _24463_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_247_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13965_ _23929_/Q VGND VGND VPWR VPWR _13965_/X sky130_fd_sc_hd__buf_2
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15704_ _15704_/A VGND VGND VPWR VPWR _16539_/A sky130_fd_sc_hd__buf_2
X_12916_ _12889_/X _12914_/X _12915_/X VGND VGND VPWR VPWR _25383_/D sky130_fd_sc_hd__and3_4
X_19472_ _23724_/Q VGND VGND VPWR VPWR _19472_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16684_ _16684_/A VGND VGND VPWR VPWR _22684_/A sky130_fd_sc_hd__inv_2
XFILLER_74_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__23937__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13896_ _13895_/X VGND VGND VPWR VPWR _13896_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18423_ _22883_/A _24176_/Q _16217_/Y _18467_/A VGND VGND VPWR VPWR _18423_/X sky130_fd_sc_hd__o22a_4
X_15635_ _21124_/A _15553_/A _15475_/X _15553_/A VGND VGND VPWR VPWR _15635_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_221_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12847_ _25399_/Q _12847_/B VGND VGND VPWR VPWR _12847_/X sky130_fd_sc_hd__or2_4
X_18354_ _18354_/A _18353_/X VGND VGND VPWR VPWR _18354_/Y sky130_fd_sc_hd__nand2_4
X_15566_ _15566_/A VGND VGND VPWR VPWR _15566_/Y sky130_fd_sc_hd__inv_2
X_12778_ _12768_/X _12771_/X _12778_/C _12778_/D VGND VGND VPWR VPWR _12778_/X sky130_fd_sc_hd__or4_4
XFILLER_15_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22745__A _24800_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17329_/A _17248_/Y _17304_/X VGND VGND VPWR VPWR _17305_/X sky130_fd_sc_hd__or3_4
X_14517_ _25104_/Q _14499_/X _21347_/A _14494_/X VGND VGND VPWR VPWR _14517_/X sky130_fd_sc_hd__o22a_4
XANTENNA__16890__A1_N _22191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11729_ HWDATA[15] VGND VGND VPWR VPWR _16226_/A sky130_fd_sc_hd__buf_2
X_18285_ _18285_/A _18285_/B _18284_/X VGND VGND VPWR VPWR _18285_/X sky130_fd_sc_hd__or3_4
X_15497_ _15496_/Y _15494_/X HADDR[18] _15494_/X VGND VGND VPWR VPWR _15497_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17236_ _17236_/A _17183_/Y VGND VGND VPWR VPWR _17236_/X sky130_fd_sc_hd__or2_4
XFILLER_30_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14448_ _14455_/A VGND VGND VPWR VPWR _14448_/X sky130_fd_sc_hd__buf_2
XFILLER_80_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16390__B1 _16301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_196_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17167_ _24618_/Q _17366_/A _16289_/Y _24368_/Q VGND VGND VPWR VPWR _17167_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22463__B1 _13800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24796__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14379_ _20467_/C VGND VGND VPWR VPWR _20506_/D sky130_fd_sc_hd__inv_2
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16118_ _22870_/A VGND VGND VPWR VPWR _16118_/Y sky130_fd_sc_hd__inv_2
XANTENNA__24725__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17098_ _17030_/C _17098_/B VGND VGND VPWR VPWR _17099_/D sky130_fd_sc_hd__or2_4
XFILLER_131_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_8_151_0_HCLK clkbuf_7_75_0_HCLK/X VGND VGND VPWR VPWR _24159_/CLK sky130_fd_sc_hd__clkbuf_1
X_16049_ _24725_/Q VGND VGND VPWR VPWR _16049_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21096__A _21085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19808_ _22364_/B _19806_/X _19807_/X _19806_/X VGND VGND VPWR VPWR _23610_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12511__A _12511_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14456__B1 _14384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15799__A3 _15721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19739_ _19738_/X VGND VGND VPWR VPWR _19740_/A sky130_fd_sc_hd__inv_2
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22750_ _24627_/Q _21337_/X VGND VGND VPWR VPWR _22750_/X sky130_fd_sc_hd__or2_4
XFILLER_71_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21701_ _24788_/Q _23002_/A VGND VGND VPWR VPWR _21701_/X sky130_fd_sc_hd__or2_4
XFILLER_240_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__25513__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22681_ _21111_/X _22679_/X _22696_/B _22680_/X VGND VGND VPWR VPWR _22681_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__19147__B1 _19122_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24420_ _24419_/CLK _16842_/X HRESETn VGND VGND VPWR VPWR _14885_/A sky130_fd_sc_hd__dfrtp_4
X_21632_ _21626_/X _21631_/X _14707_/X VGND VGND VPWR VPWR _21632_/X sky130_fd_sc_hd__o21a_4
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__22297__A3 _22296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24351_ _24667_/CLK _17354_/Y HRESETn VGND VGND VPWR VPWR _17171_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_221_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21563_ _21563_/A VGND VGND VPWR VPWR _21564_/D sky130_fd_sc_hd__inv_2
XFILLER_178_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__17749__A _21059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15708__B1 _24886_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23302_ _24476_/Q _22661_/X _23178_/X VGND VGND VPWR VPWR _23302_/X sky130_fd_sc_hd__o21a_4
XFILLER_178_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20514_ _13962_/A _20514_/B _20514_/C VGND VGND VPWR VPWR _20514_/X sky130_fd_sc_hd__or3_4
X_24282_ _24263_/CLK _17803_/Y HRESETn VGND VGND VPWR VPWR _16906_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21494_ _21463_/A VGND VGND VPWR VPWR _21657_/A sky130_fd_sc_hd__buf_2
X_23233_ _15559_/Y _23292_/B VGND VGND VPWR VPWR _23233_/X sky130_fd_sc_hd__and2_4
X_20445_ _20445_/A _20444_/B VGND VGND VPWR VPWR _20447_/C sky130_fd_sc_hd__and2_4
X_23164_ _16652_/Y _23291_/B VGND VGND VPWR VPWR _23164_/X sky130_fd_sc_hd__and2_4
XFILLER_180_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24466__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20376_ _20374_/Y _20375_/Y _19746_/X _20375_/Y VGND VGND VPWR VPWR _23399_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21009__A1 _23968_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22115_ _13492_/Y _12086_/A _12019_/Y _21571_/X VGND VGND VPWR VPWR _22115_/X sky130_fd_sc_hd__o22a_4
XANTENNA__22821__C _22505_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23095_ _12760_/Y _21437_/X _22280_/X _12527_/Y _21085_/X VGND VGND VPWR VPWR _23095_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_121_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22046_ _22045_/X VGND VGND VPWR VPWR _22046_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12421__A _12248_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23997_ _24973_/CLK _20680_/X HRESETn VGND VGND VPWR VPWR _23997_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13750_ _20157_/D VGND VGND VPWR VPWR _19898_/D sky130_fd_sc_hd__buf_2
XFILLER_44_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22948_ _12248_/Y _23268_/A _22947_/X VGND VGND VPWR VPWR _22948_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__25254__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12701_ _12686_/A _12701_/B _12701_/C VGND VGND VPWR VPWR _12701_/X sky130_fd_sc_hd__and3_4
X_13681_ _13680_/X _13681_/B VGND VGND VPWR VPWR _13681_/X sky130_fd_sc_hd__or2_4
XANTENNA__15947__B1 _15946_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22879_ _22786_/X _22877_/X _22789_/X _22878_/X VGND VGND VPWR VPWR _22880_/B sky130_fd_sc_hd__o22a_4
Xclkbuf_4_14_0_HCLK clkbuf_3_7_0_HCLK/X VGND VGND VPWR VPWR clkbuf_5_29_0_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_15420_ _15419_/X VGND VGND VPWR VPWR _24976_/D sky130_fd_sc_hd__inv_2
XFILLER_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12632_ _12503_/A _12632_/B VGND VGND VPWR VPWR _12634_/B sky130_fd_sc_hd__or2_4
X_24618_ _24618_/CLK _24618_/D HRESETn VGND VGND VPWR VPWR _24618_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15962__A3 _16236_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _12671_/A _24872_/Q _12657_/A _12514_/Y VGND VGND VPWR VPWR _12563_/X sky130_fd_sc_hd__a2bb2o_4
X_15351_ _15351_/A _15349_/A VGND VGND VPWR VPWR _15352_/C sky130_fd_sc_hd__or2_4
X_24549_ _24520_/CLK _24549_/D HRESETn VGND VGND VPWR VPWR _24549_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22693__B1 _23062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14302_ _25176_/Q _14291_/X _25175_/Q _14296_/X VGND VGND VPWR VPWR _14302_/X sky130_fd_sc_hd__o22a_4
X_18070_ _17979_/X _18070_/B VGND VGND VPWR VPWR _18070_/X sky130_fd_sc_hd__or2_4
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _12494_/A VGND VGND VPWR VPWR _13087_/A sky130_fd_sc_hd__buf_2
X_15282_ _14902_/A _15282_/B VGND VGND VPWR VPWR _15282_/X sky130_fd_sc_hd__or2_4
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17021_ _17020_/Y VGND VGND VPWR VPWR _17062_/A sky130_fd_sc_hd__buf_2
XFILLER_156_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14233_ _13954_/A _14233_/B VGND VGND VPWR VPWR _14234_/B sky130_fd_sc_hd__or2_4
XFILLER_184_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14083__A _14083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14164_ _14158_/Y _14099_/X _14100_/X _14163_/X VGND VGND VPWR VPWR _14164_/X sky130_fd_sc_hd__o22a_4
XFILLER_125_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13115_ _20709_/A _20704_/A VGND VGND VPWR VPWR _13116_/B sky130_fd_sc_hd__or2_4
XFILLER_180_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__24136__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_8_224_0_HCLK clkbuf_7_112_0_HCLK/X VGND VGND VPWR VPWR _24326_/CLK sky130_fd_sc_hd__clkbuf_1
X_14095_ _14095_/A _14093_/Y _14094_/Y VGND VGND VPWR VPWR _14095_/X sky130_fd_sc_hd__and3_4
X_18972_ _18210_/B VGND VGND VPWR VPWR _18972_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13046_ _13046_/A _13046_/B VGND VGND VPWR VPWR _13046_/X sky130_fd_sc_hd__or2_4
X_17923_ _17921_/Y _17926_/A _17917_/B VGND VGND VPWR VPWR _17924_/A sky130_fd_sc_hd__or3_4
XFILLER_239_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12341__A2_N _24833_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13427__A _13285_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17854_ _16915_/Y _17849_/X _16895_/X _17862_/B VGND VGND VPWR VPWR _17854_/X sky130_fd_sc_hd__or4_4
XFILLER_66_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14438__B1 _14384_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16805_ _16803_/Y _16804_/X _15719_/X _16804_/X VGND VGND VPWR VPWR _16805_/X sky130_fd_sc_hd__a2bb2o_4
X_17785_ _17784_/X VGND VGND VPWR VPWR _24286_/D sky130_fd_sc_hd__inv_2
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14997_ _14992_/X _14997_/B _14997_/C _14996_/X VGND VGND VPWR VPWR _14997_/X sky130_fd_sc_hd__or4_4
X_19524_ _16721_/A _16721_/B _13763_/X _19523_/Y VGND VGND VPWR VPWR _19524_/X sky130_fd_sc_hd__and4_4
XFILLER_235_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16736_ _15046_/Y _16735_/X _16382_/X _16735_/X VGND VGND VPWR VPWR _24472_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__21363__B _21343_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13948_ _13947_/X VGND VGND VPWR VPWR _13948_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0_HCLK clkbuf_0_HCLK/X VGND VGND VPWR VPWR clkbuf_1_1_0_HCLK/X sky130_fd_sc_hd__clkbuf_1
X_19455_ _19455_/A _19455_/B _18283_/X VGND VGND VPWR VPWR _19455_/X sky130_fd_sc_hd__or3_4
XFILLER_222_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16667_ _24499_/Q VGND VGND VPWR VPWR _16667_/Y sky130_fd_sc_hd__inv_2
X_13879_ _24974_/Q _24973_/Q _13879_/C VGND VGND VPWR VPWR _13879_/X sky130_fd_sc_hd__or3_4
XANTENNA__19129__B1 _19057_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18406_ _18399_/X _18401_/X _18404_/X _18406_/D VGND VGND VPWR VPWR _18406_/X sky130_fd_sc_hd__or4_4
X_15618_ _15618_/A VGND VGND VPWR VPWR _22291_/A sky130_fd_sc_hd__inv_2
XFILLER_179_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19386_ _17955_/B VGND VGND VPWR VPWR _19386_/Y sky130_fd_sc_hd__inv_2
X_16598_ _16598_/A VGND VGND VPWR VPWR _16598_/X sky130_fd_sc_hd__buf_2
XFILLER_15_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__22475__A _21087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18337_ _20220_/B VGND VGND VPWR VPWR _18932_/B sky130_fd_sc_hd__buf_2
XFILLER_194_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15549_ _24923_/Q VGND VGND VPWR VPWR _15549_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24977__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18268_ _18268_/A VGND VGND VPWR VPWR _18268_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__24906__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_17219_ _23012_/A VGND VGND VPWR VPWR _17219_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22436__B1 _11755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18199_ _18103_/A _19362_/A VGND VGND VPWR VPWR _18199_/X sky130_fd_sc_hd__or2_4
Xclkbuf_6_34_0_HCLK clkbuf_6_35_0_HCLK/A VGND VGND VPWR VPWR clkbuf_7_69_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20230_ _20229_/Y _20227_/X _15762_/X _20227_/X VGND VGND VPWR VPWR _23455_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20161_ _20161_/A VGND VGND VPWR VPWR _20161_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22739__A1 _22520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20092_ _24412_/Q VGND VGND VPWR VPWR _20092_/X sky130_fd_sc_hd__buf_2
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23920_ _23912_/CLK _23920_/D VGND VGND VPWR VPWR _18917_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_130_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14429__B1 _14403_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_245_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23851_ _23853_/CLK _23851_/D VGND VGND VPWR VPWR _19113_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16648__A _16655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__19368__B1 _19301_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22802_ _23178_/A VGND VGND VPWR VPWR _22802_/X sky130_fd_sc_hd__buf_2
XFILLER_38_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20994_ _20994_/A _20994_/B VGND VGND VPWR VPWR _23364_/A sky130_fd_sc_hd__and2_4
X_23782_ _24252_/CLK _19311_/X VGND VGND VPWR VPWR _19310_/A sky130_fd_sc_hd__dfxtp_4
X_25521_ _25521_/CLK _25521_/D HRESETn VGND VGND VPWR VPWR _25521_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22733_ _22539_/A _22733_/B _22732_/X VGND VGND VPWR VPWR _22733_/X sky130_fd_sc_hd__and3_4
XFILLER_26_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22664_ _22572_/X _22660_/Y _21056_/X _22663_/X VGND VGND VPWR VPWR _22665_/D sky130_fd_sc_hd__a2bb2o_4
X_25452_ _24766_/CLK _12430_/X HRESETn VGND VGND VPWR VPWR _12201_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21615_ _14753_/X _21615_/B VGND VGND VPWR VPWR _21615_/X sky130_fd_sc_hd__or2_4
X_24403_ _23427_/CLK _24403_/D HRESETn VGND VGND VPWR VPWR _24403_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_7_116_0_HCLK clkbuf_6_58_0_HCLK/X VGND VGND VPWR VPWR clkbuf_7_116_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_22595_ _21109_/A _22594_/X _22135_/C _24866_/Q _21098_/A VGND VGND VPWR VPWR _22595_/X
+ sky130_fd_sc_hd__a32o_4
X_25383_ _25382_/CLK _25383_/D HRESETn VGND VGND VPWR VPWR _12800_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_138_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_21546_ _17242_/B _22543_/A _25370_/Q _21423_/A VGND VGND VPWR VPWR _21546_/X sky130_fd_sc_hd__a2bb2o_4
X_24334_ _25243_/CLK _24334_/D HRESETn VGND VGND VPWR VPWR _24334_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24647__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16354__B1 _16353_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24265_ _24686_/CLK _17872_/X HRESETn VGND VGND VPWR VPWR _24265_/Q sky130_fd_sc_hd__dfrtp_4
X_21477_ _21453_/X _21469_/X _21477_/C VGND VGND VPWR VPWR _21477_/X sky130_fd_sc_hd__or3_4
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23216_ _23216_/A _22658_/B VGND VGND VPWR VPWR _23216_/X sky130_fd_sc_hd__or2_4
X_20428_ _15482_/B VGND VGND VPWR VPWR _20429_/B sky130_fd_sc_hd__inv_2
X_24196_ _25471_/CLK _24196_/D HRESETn VGND VGND VPWR VPWR _24196_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12391__A1 _12264_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22551__C _22550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23147_ _23103_/A _23146_/X VGND VGND VPWR VPWR _23147_/X sky130_fd_sc_hd__and2_4
X_20359_ _20359_/A VGND VGND VPWR VPWR _21806_/B sky130_fd_sc_hd__inv_2
X_23078_ _23078_/A _22423_/A VGND VGND VPWR VPWR _23081_/B sky130_fd_sc_hd__or2_4
XFILLER_49_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14920_ _25027_/Q VGND VGND VPWR VPWR _14921_/A sky130_fd_sc_hd__inv_2
X_22029_ _21670_/X _22029_/B VGND VGND VPWR VPWR _22029_/X sky130_fd_sc_hd__or2_4
XFILLER_248_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_8_54_0_HCLK clkbuf_8_55_0_HCLK/A VGND VGND VPWR VPWR _24236_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_49_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__25435__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14851_ _14823_/X _14850_/X _24957_/Q _14830_/X VGND VGND VPWR VPWR _14851_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_248_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13802_ _14395_/A _14442_/A VGND VGND VPWR VPWR _17410_/A sky130_fd_sc_hd__or2_4
XFILLER_29_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17570_ _17523_/Y _17646_/A _17569_/X VGND VGND VPWR VPWR _17570_/X sky130_fd_sc_hd__or3_4
XFILLER_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24954__SET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14782_ _18052_/A VGND VGND VPWR VPWR _18020_/A sky130_fd_sc_hd__buf_2
XFILLER_217_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11994_ _11979_/X VGND VGND VPWR VPWR _11994_/Y sky130_fd_sc_hd__inv_2
X_16521_ _16521_/A VGND VGND VPWR VPWR _16521_/X sky130_fd_sc_hd__buf_2
X_13733_ _13732_/X VGND VGND VPWR VPWR _13733_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__20913__B1 _20855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_19240_ _23807_/Q VGND VGND VPWR VPWR _19240_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16452_ _16724_/A _16540_/B VGND VGND VPWR VPWR _16453_/A sky130_fd_sc_hd__nor2_4
XFILLER_231_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13664_ _13682_/A VGND VGND VPWR VPWR _13664_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16593__B1 _16240_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15403_ _15386_/X _15401_/Y _15402_/X VGND VGND VPWR VPWR _15403_/X sky130_fd_sc_hd__and3_4
X_12615_ _12648_/A _12615_/B _12615_/C VGND VGND VPWR VPWR _25432_/D sky130_fd_sc_hd__and3_4
X_19171_ _19169_/Y _19165_/X _19125_/X _19170_/X VGND VGND VPWR VPWR _23832_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16383_ _16380_/Y _16381_/X _16382_/X _16381_/X VGND VGND VPWR VPWR _24606_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13595_ _13594_/X VGND VGND VPWR VPWR _13596_/B sky130_fd_sc_hd__inv_2
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18122_ _18014_/A _18122_/B VGND VGND VPWR VPWR _18123_/C sky130_fd_sc_hd__or2_4
X_15334_ _15282_/B VGND VGND VPWR VPWR _15334_/X sky130_fd_sc_hd__buf_2
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__24388__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12546_ _12507_/X _12519_/X _12532_/X _12546_/D VGND VGND VPWR VPWR _12588_/A sky130_fd_sc_hd__or4_4
XANTENNA__16345__B1 _16059_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18053_ _18053_/A _18053_/B VGND VGND VPWR VPWR _18056_/B sky130_fd_sc_hd__or2_4
XFILLER_185_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22418__B1 _22290_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24317__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15265_ _15265_/A _15269_/B VGND VGND VPWR VPWR _15265_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__16896__B2 _24284_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12477_ _12197_/Y _12480_/B _12382_/X VGND VGND VPWR VPWR _12477_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_126_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17004_ _24393_/Q VGND VGND VPWR VPWR _17004_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14216_ _14215_/Y _14213_/X _13826_/X _14213_/X VGND VGND VPWR VPWR _14216_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15196_ _15195_/X VGND VGND VPWR VPWR _25032_/D sky130_fd_sc_hd__inv_2
XANTENNA__22433__A3 _22432_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14147_ _14133_/X _14146_/Y _14103_/C _14133_/X VGND VGND VPWR VPWR _25216_/D sky130_fd_sc_hd__a2bb2o_4
XANTENNA__15637__A _22111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14078_ _14054_/A VGND VGND VPWR VPWR _20541_/B sky130_fd_sc_hd__buf_2
X_18955_ _17959_/B VGND VGND VPWR VPWR _18955_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__18948__A _19063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13029_ _13028_/X VGND VGND VPWR VPWR _25357_/D sky130_fd_sc_hd__inv_2
X_17906_ _17906_/A _17906_/B VGND VGND VPWR VPWR _17908_/A sky130_fd_sc_hd__or2_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18886_ _23950_/Q _18884_/A VGND VGND VPWR VPWR _18886_/X sky130_fd_sc_hd__or2_4
XFILLER_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__23952__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__25176__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17837_ _17818_/A _17837_/B _17836_/X VGND VGND VPWR VPWR _17837_/X sky130_fd_sc_hd__and3_4
XANTENNA__12295__A2_N _12293_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__25105__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17768_ _16913_/Y _16945_/X _17768_/C _17768_/D VGND VGND VPWR VPWR _17769_/A sky130_fd_sc_hd__or4_4
XFILLER_66_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21157__B1 _14876_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16719_ _16719_/A VGND VGND VPWR VPWR _22844_/A sky130_fd_sc_hd__buf_2
X_19507_ _23712_/Q VGND VGND VPWR VPWR _22027_/B sky130_fd_sc_hd__inv_2
X_17699_ _17529_/A _17698_/Y VGND VGND VPWR VPWR _17700_/B sky130_fd_sc_hd__or2_4
X_19438_ _19437_/Y _19435_/X _19392_/X _19435_/X VGND VGND VPWR VPWR _19438_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19369_ _23761_/Q VGND VGND VPWR VPWR _19369_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__14716__A _13731_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21400_ _22213_/A _21391_/X _21399_/X VGND VGND VPWR VPWR _21400_/X sky130_fd_sc_hd__or3_4
XFILLER_210_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13620__A _13579_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22380_ _22380_/A _22378_/X _22379_/X VGND VGND VPWR VPWR _22380_/X sky130_fd_sc_hd__and3_4
XANTENNA__12070__B1 _11781_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21712__A1_N _17241_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24740__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21331_ _16786_/A _21309_/X _22891_/A VGND VGND VPWR VPWR _21331_/X sky130_fd_sc_hd__o21a_4
XFILLER_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22409__B1 _22407_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24058__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__21880__B2 _21431_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24050_ _24051_/CLK _24050_/D HRESETn VGND VGND VPWR VPWR _13650_/C sky130_fd_sc_hd__dfrtp_4
X_21262_ _21262_/A _19851_/Y VGND VGND VPWR VPWR _21262_/X sky130_fd_sc_hd__or2_4
XANTENNA__23082__B1 _16906_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17746__B _16906_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23001_ _23001_/A VGND VGND VPWR VPWR _23001_/X sky130_fd_sc_hd__buf_2
XFILLER_144_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20213_ _20200_/Y VGND VGND VPWR VPWR _20213_/X sky130_fd_sc_hd__buf_2
XANTENNA__15547__A _16637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21193_ _21209_/A _21193_/B VGND VGND VPWR VPWR _21193_/X sky130_fd_sc_hd__or2_4
XFILLER_131_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20144_ _20142_/Y _20138_/X _20095_/X _20143_/X VGND VGND VPWR VPWR _23488_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__22188__A2 _22174_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17762__A _17755_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20075_ _20074_/Y _20072_/X _19817_/X _20072_/X VGND VGND VPWR VPWR _20075_/X sky130_fd_sc_hd__a2bb2o_4
X_24952_ _24953_/CLK _15474_/X HRESETn VGND VGND VPWR VPWR _24952_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_98_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12402__C _12370_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23903_ _25171_/CLK _18963_/X VGND VGND VPWR VPWR _18078_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_245_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24883_ _24872_/CLK _15716_/X HRESETn VGND VGND VPWR VPWR _24883_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23834_ _24089_/CLK _19166_/X VGND VGND VPWR VPWR _19162_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_45_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__21699__A1 _16637_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _20467_/A _23924_/Q _14530_/A VGND VGND VPWR VPWR _20977_/X sky130_fd_sc_hd__a21o_4
X_23765_ _23767_/CLK _19358_/X VGND VGND VPWR VPWR _18135_/B sky130_fd_sc_hd__dfxtp_4
XANTENNA__22896__B1 _22880_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21699__B2 _22522_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24899__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25504_ _23691_/CLK _11925_/X HRESETn VGND VGND VPWR VPWR _19984_/A sky130_fd_sc_hd__dfrtp_4
XPHY_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22716_ _22716_/A _22713_/X _22715_/X VGND VGND VPWR VPWR _22716_/X sky130_fd_sc_hd__and3_4
XANTENNA__24828__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16575__B1 _16400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23696_ _23406_/CLK _23696_/D VGND VGND VPWR VPWR _23696_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__20628__A _20628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25435_ _25444_/CLK _25435_/D HRESETn VGND VGND VPWR VPWR _25435_/Q sky130_fd_sc_hd__dfrtp_4
X_22647_ _12920_/A _22572_/X _22646_/X VGND VGND VPWR VPWR _22647_/X sky130_fd_sc_hd__o21a_4
XANTENNA__14626__A _18060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__22112__A2 _21019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12400_ _12398_/X _12400_/B _12399_/X VGND VGND VPWR VPWR _12401_/A sky130_fd_sc_hd__or3_4
X_13380_ _13254_/A _13378_/X _13380_/C VGND VGND VPWR VPWR _13380_/X sky130_fd_sc_hd__and3_4
XFILLER_167_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12061__B1 _11761_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__24481__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22578_ _24591_/Q _22532_/B VGND VGND VPWR VPWR _22581_/B sky130_fd_sc_hd__or2_4
X_25366_ _25387_/CLK _25366_/D HRESETn VGND VGND VPWR VPWR _12282_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_222_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22663__A3 _22138_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12331_ _12344_/A _12329_/Y _12330_/Y _24825_/Q VGND VGND VPWR VPWR _12339_/A sky130_fd_sc_hd__a2bb2o_4
X_24317_ _24317_/CLK _17613_/Y HRESETn VGND VGND VPWR VPWR _24317_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__24410__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21529_ _21520_/X _21528_/X _21522_/X _24857_/Q _22522_/B VGND VGND VPWR VPWR _21530_/B
+ sky130_fd_sc_hd__a32o_4
X_25297_ _23916_/CLK _25297_/D HRESETn VGND VGND VPWR VPWR _25297_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12146__A _18372_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12262_ _12261_/X VGND VGND VPWR VPWR _12263_/A sky130_fd_sc_hd__buf_2
X_15050_ _15028_/X _15035_/X _15042_/X _15049_/X VGND VGND VPWR VPWR _15050_/X sky130_fd_sc_hd__or4_4
X_24248_ _23774_/CLK _18025_/X HRESETn VGND VGND VPWR VPWR _24248_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16674__A1_N _16672_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14353__A2 _14340_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__23073__B1 _23060_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14001_ _14001_/A _14028_/B _14000_/Y _13980_/X VGND VGND VPWR VPWR _14002_/B sky130_fd_sc_hd__or4_4
XANTENNA__15457__A _15457_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12364__B2 _24824_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12193_ _25441_/Q _24756_/Q _12191_/X _12192_/Y VGND VGND VPWR VPWR _12193_/X sky130_fd_sc_hd__o22a_4
X_24179_ _24188_/CLK _24179_/D HRESETn VGND VGND VPWR VPWR _18528_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_162_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18740_ _18734_/A _18730_/B _18739_/X VGND VGND VPWR VPWR _24149_/D sky130_fd_sc_hd__and3_4
XFILLER_110_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15952_ _12188_/Y _15949_/X _15951_/X _15949_/X VGND VGND VPWR VPWR _15952_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14903_ _15056_/D VGND VGND VPWR VPWR _14903_/X sky130_fd_sc_hd__buf_2
X_18671_ _18705_/B VGND VGND VPWR VPWR _18744_/A sky130_fd_sc_hd__buf_2
X_15883_ _15879_/X _15880_/X _16226_/A _24800_/Q _15881_/X VGND VGND VPWR VPWR _15883_/X
+ sky130_fd_sc_hd__a32o_4
X_17622_ _17563_/A _17621_/Y VGND VGND VPWR VPWR _17622_/X sky130_fd_sc_hd__or2_4
X_14834_ _14833_/X VGND VGND VPWR VPWR _14834_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16612__A1_N _16610_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17553_ _17553_/A _17550_/X _17551_/X _17553_/D VGND VGND VPWR VPWR _17553_/X sky130_fd_sc_hd__or4_4
X_14765_ _14765_/A _14756_/A _13577_/B VGND VGND VPWR VPWR _14776_/B sky130_fd_sc_hd__and3_4
XANTENNA__19599__A _19598_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11977_ _11977_/A _11977_/B VGND VGND VPWR VPWR _11977_/X sky130_fd_sc_hd__and2_4
XFILLER_205_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16504_ _16503_/Y _16501_/X _16233_/X _16501_/X VGND VGND VPWR VPWR _16504_/X sky130_fd_sc_hd__a2bb2o_4
XANTENNA__19752__B1 _19728_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13716_ _13669_/A _13668_/X VGND VGND VPWR VPWR _13716_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__15920__A _19646_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17484_ _17460_/A _17481_/B _17482_/Y VGND VGND VPWR VPWR _17485_/A sky130_fd_sc_hd__o21a_4
XFILLER_232_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24569__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14696_ _21901_/A _14695_/X _21901_/A _14695_/X VGND VGND VPWR VPWR _14696_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19223_ _23813_/Q VGND VGND VPWR VPWR _19223_/Y sky130_fd_sc_hd__inv_2
X_16435_ _19063_/A VGND VGND VPWR VPWR _16435_/X sky130_fd_sc_hd__buf_2
XFILLER_177_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__22639__B1 _25532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13647_ _24045_/Q _13647_/B VGND VGND VPWR VPWR _13648_/B sky130_fd_sc_hd__or2_4
XFILLER_32_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__22103__A2 _21365_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19154_ _19153_/Y _19149_/X _19106_/X _19149_/X VGND VGND VPWR VPWR _19154_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16366_ _16366_/A _16366_/B VGND VGND VPWR VPWR _16366_/X sky130_fd_sc_hd__or2_4
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _15694_/A VGND VGND VPWR VPWR _13579_/B sky130_fd_sc_hd__inv_2
X_18105_ _18030_/A _18105_/B _18104_/X VGND VGND VPWR VPWR _18109_/B sky130_fd_sc_hd__and3_4
XFILLER_118_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15317_ _25005_/Q _15316_/Y VGND VGND VPWR VPWR _15317_/X sky130_fd_sc_hd__or2_4
XFILLER_158_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__24151__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12529_ _25408_/Q VGND VGND VPWR VPWR _12706_/A sky130_fd_sc_hd__inv_2
X_19085_ _19085_/A VGND VGND VPWR VPWR _21615_/B sky130_fd_sc_hd__inv_2
XFILLER_9_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_16297_ _24636_/Q VGND VGND VPWR VPWR _16297_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__22472__B _22472_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18036_ _17985_/X _18036_/B VGND VGND VPWR VPWR _18036_/X sky130_fd_sc_hd__or2_4
X_15248_ _25019_/Q _15248_/B VGND VGND VPWR VPWR _15250_/B sky130_fd_sc_hd__or2_4
XFILLER_173_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12355__B2 _12354_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11895__A _19600_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15179_ _15067_/B _15311_/B VGND VGND VPWR VPWR _15180_/A sky130_fd_sc_hd__or2_4
XANTENNA__21088__B _22420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__25357__RESET_B HRESETn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19987_ _21185_/B _19980_/X _19874_/X _19962_/Y VGND VGND VPWR VPWR _19987_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18938_ _18938_/A VGND VGND VPWR VPWR _18938_/Y sky130_fd_sc_hd__inv_2
.ends

